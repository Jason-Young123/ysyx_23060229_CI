//Generate the verilog at 2025-09-29T17:15:11 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_B ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ;
wire \myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

AND3_X4 _08999_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [1] ), .A3(\myclint.mtime [0] ), .ZN(_01489_ ) );
AND3_X4 _09000_ ( .A1(_01489_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01490_ ) );
AND3_X4 _09001_ ( .A1(_01490_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01491_ ) );
AND3_X4 _09002_ ( .A1(_01491_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01492_ ) );
AND3_X4 _09003_ ( .A1(_01492_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01493_ ) );
AND3_X4 _09004_ ( .A1(_01493_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01494_ ) );
AND3_X4 _09005_ ( .A1(_01494_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01495_ ) );
AND3_X4 _09006_ ( .A1(_01495_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01496_ ) );
AND3_X4 _09007_ ( .A1(_01496_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01497_ ) );
AND3_X4 _09008_ ( .A1(_01497_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01498_ ) );
AND3_X4 _09009_ ( .A1(_01498_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01499_ ) );
AND3_X4 _09010_ ( .A1(_01499_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01500_ ) );
AND3_X4 _09011_ ( .A1(_01500_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01501_ ) );
AND2_X4 _09012_ ( .A1(_01501_ ), .A2(\myclint.mtime [27] ), .ZN(_01502_ ) );
AND2_X1 _09013_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01503_ ) );
AND2_X2 _09014_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01504_ ) );
AND4_X4 _09015_ ( .A1(\myclint.mtime [33] ), .A2(_01502_ ), .A3(_01503_ ), .A4(_01504_ ), .ZN(_01505_ ) );
AND3_X2 _09016_ ( .A1(_01505_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01506_ ) );
AND3_X2 _09017_ ( .A1(_01506_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [35] ), .ZN(_01507_ ) );
AND2_X2 _09018_ ( .A1(_01507_ ), .A2(\myclint.mtime [37] ), .ZN(_01508_ ) );
AND2_X1 _09019_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [39] ), .ZN(_01509_ ) );
AND2_X2 _09020_ ( .A1(_01508_ ), .A2(_01509_ ), .ZN(_01510_ ) );
AND2_X1 _09021_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01511_ ) );
AND2_X4 _09022_ ( .A1(_01510_ ), .A2(_01511_ ), .ZN(_01512_ ) );
AND2_X1 _09023_ ( .A1(\myclint.mtime [42] ), .A2(\myclint.mtime [43] ), .ZN(_01513_ ) );
AND2_X4 _09024_ ( .A1(_01512_ ), .A2(_01513_ ), .ZN(_01514_ ) );
AND2_X1 _09025_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01515_ ) );
AND3_X1 _09026_ ( .A1(_01515_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01516_ ) );
AND2_X2 _09027_ ( .A1(_01514_ ), .A2(_01516_ ), .ZN(_01517_ ) );
AND2_X1 _09028_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01518_ ) );
AND2_X1 _09029_ ( .A1(_01517_ ), .A2(_01518_ ), .ZN(_01519_ ) );
AND2_X1 _09030_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01520_ ) );
AND2_X2 _09031_ ( .A1(_01519_ ), .A2(_01520_ ), .ZN(_01521_ ) );
AND2_X1 _09032_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01522_ ) );
AND2_X2 _09033_ ( .A1(_01521_ ), .A2(_01522_ ), .ZN(_01523_ ) );
AND2_X1 _09034_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01524_ ) );
AND2_X2 _09035_ ( .A1(_01523_ ), .A2(_01524_ ), .ZN(_01525_ ) );
AND2_X1 _09036_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01526_ ) );
AND2_X2 _09037_ ( .A1(_01525_ ), .A2(_01526_ ), .ZN(_01527_ ) );
AND2_X1 _09038_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01528_ ) );
AND2_X2 _09039_ ( .A1(_01527_ ), .A2(_01528_ ), .ZN(_01529_ ) );
INV_X1 _09040_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01530_ ) );
AND2_X1 _09041_ ( .A1(\myclint.mtime [60] ), .A2(\myclint.mtime [61] ), .ZN(_01531_ ) );
AND3_X4 _09042_ ( .A1(_01529_ ), .A2(_01530_ ), .A3(_01531_ ), .ZN(_01532_ ) );
AND2_X1 _09043_ ( .A1(_01532_ ), .A2(\myclint.mtime [63] ), .ZN(_01533_ ) );
INV_X1 _09044_ ( .A(fanout_net_1 ), .ZN(_01534_ ) );
BUF_X4 _09045_ ( .A(_01534_ ), .Z(_01535_ ) );
BUF_X4 _09046_ ( .A(_01535_ ), .Z(_01536_ ) );
OAI21_X1 _09047_ ( .A(_01536_ ), .B1(_01532_ ), .B2(\myclint.mtime [63] ), .ZN(_01537_ ) );
NOR2_X1 _09048_ ( .A1(_01533_ ), .A2(_01537_ ), .ZN(_00000_ ) );
AND2_X1 _09049_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_01538_ ) );
AND3_X1 _09050_ ( .A1(_01538_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01539_ ) );
AND4_X1 _09051_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01540_ ) );
AND2_X1 _09052_ ( .A1(_01539_ ), .A2(_01540_ ), .ZN(_01541_ ) );
AND2_X1 _09053_ ( .A1(\myclint.mtime [24] ), .A2(\myclint.mtime [25] ), .ZN(_01542_ ) );
AND3_X1 _09054_ ( .A1(_01542_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [27] ), .ZN(_01543_ ) );
NAND4_X1 _09055_ ( .A1(_01541_ ), .A2(_01503_ ), .A3(_01504_ ), .A4(_01543_ ), .ZN(_01544_ ) );
AND2_X1 _09056_ ( .A1(_01489_ ), .A2(\myclint.mtime [3] ), .ZN(_01545_ ) );
AND4_X1 _09057_ ( .A1(\myclint.mtime [6] ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [5] ), .A4(\myclint.mtime [7] ), .ZN(_01546_ ) );
AND2_X1 _09058_ ( .A1(_01545_ ), .A2(_01546_ ), .ZN(_01547_ ) );
AND4_X1 _09059_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01548_ ) );
AND2_X1 _09060_ ( .A1(\myclint.mtime [8] ), .A2(\myclint.mtime [9] ), .ZN(_01549_ ) );
AND4_X1 _09061_ ( .A1(\myclint.mtime [10] ), .A2(_01548_ ), .A3(\myclint.mtime [11] ), .A4(_01549_ ), .ZN(_01550_ ) );
NAND2_X1 _09062_ ( .A1(_01547_ ), .A2(_01550_ ), .ZN(_01551_ ) );
NOR2_X1 _09063_ ( .A1(_01544_ ), .A2(_01551_ ), .ZN(_01552_ ) );
AND2_X1 _09064_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01553_ ) );
AND3_X1 _09065_ ( .A1(_01553_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01554_ ) );
AND2_X1 _09066_ ( .A1(_01513_ ), .A2(_01511_ ), .ZN(_01555_ ) );
AND4_X1 _09067_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01556_ ) );
AND4_X1 _09068_ ( .A1(_01516_ ), .A2(_01554_ ), .A3(_01555_ ), .A4(_01556_ ), .ZN(_01557_ ) );
AND2_X1 _09069_ ( .A1(_01552_ ), .A2(_01557_ ), .ZN(_01558_ ) );
AND4_X1 _09070_ ( .A1(_01524_ ), .A2(_01522_ ), .A3(_01520_ ), .A4(_01518_ ), .ZN(_01559_ ) );
AND2_X1 _09071_ ( .A1(_01558_ ), .A2(_01559_ ), .ZN(_01560_ ) );
AND4_X1 _09072_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01561_ ) );
NAND3_X1 _09073_ ( .A1(_01560_ ), .A2(_01531_ ), .A3(_01561_ ), .ZN(_01562_ ) );
OR2_X1 _09074_ ( .A1(_01562_ ), .A2(\myclint.mtime [62] ), .ZN(_01563_ ) );
NAND2_X1 _09075_ ( .A1(_01562_ ), .A2(\myclint.mtime [62] ), .ZN(_01564_ ) );
AOI21_X1 _09076_ ( .A(fanout_net_1 ), .B1(_01563_ ), .B2(_01564_ ), .ZN(_00001_ ) );
AND2_X1 _09077_ ( .A1(_01520_ ), .A2(_01518_ ), .ZN(_01565_ ) );
NAND2_X1 _09078_ ( .A1(_01558_ ), .A2(_01565_ ), .ZN(_01566_ ) );
OR3_X1 _09079_ ( .A1(_01566_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [53] ), .ZN(_01567_ ) );
OAI21_X1 _09080_ ( .A(\myclint.mtime [53] ), .B1(_01566_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01568_ ) );
AOI21_X1 _09081_ ( .A(fanout_net_1 ), .B1(_01567_ ), .B2(_01568_ ), .ZN(_00002_ ) );
XNOR2_X1 _09082_ ( .A(_01566_ ), .B(\myclint.mtime [52] ), .ZN(_01569_ ) );
CLKBUF_X3 _09083_ ( .A(_01535_ ), .Z(_01570_ ) );
AND2_X1 _09084_ ( .A1(_01569_ ), .A2(_01570_ ), .ZN(_00003_ ) );
NAND3_X1 _09085_ ( .A1(_01552_ ), .A2(_01518_ ), .A3(_01557_ ), .ZN(_01571_ ) );
OR3_X1 _09086_ ( .A1(_01571_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [51] ), .ZN(_01572_ ) );
OAI21_X1 _09087_ ( .A(\myclint.mtime [51] ), .B1(_01571_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01573_ ) );
AOI21_X1 _09088_ ( .A(fanout_net_1 ), .B1(_01572_ ), .B2(_01573_ ), .ZN(_00004_ ) );
OR2_X1 _09089_ ( .A1(_01571_ ), .A2(\myclint.mtime [50] ), .ZN(_01574_ ) );
NAND2_X1 _09090_ ( .A1(_01571_ ), .A2(\myclint.mtime [50] ), .ZN(_01575_ ) );
AOI21_X1 _09091_ ( .A(fanout_net_1 ), .B1(_01574_ ), .B2(_01575_ ), .ZN(_00005_ ) );
INV_X1 _09092_ ( .A(_01514_ ), .ZN(_01576_ ) );
INV_X1 _09093_ ( .A(_01516_ ), .ZN(_01577_ ) );
NOR3_X1 _09094_ ( .A1(_01576_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01577_ ), .ZN(_01578_ ) );
AND2_X1 _09095_ ( .A1(_01578_ ), .A2(\myclint.mtime [49] ), .ZN(_01579_ ) );
OAI21_X1 _09096_ ( .A(_01536_ ), .B1(_01578_ ), .B2(\myclint.mtime [49] ), .ZN(_01580_ ) );
NOR2_X1 _09097_ ( .A1(_01579_ ), .A2(_01580_ ), .ZN(_00006_ ) );
INV_X1 _09098_ ( .A(_01552_ ), .ZN(_01581_ ) );
INV_X1 _09099_ ( .A(_01557_ ), .ZN(_01582_ ) );
OAI21_X1 _09100_ ( .A(\myclint.mtime [48] ), .B1(_01581_ ), .B2(_01582_ ), .ZN(_01583_ ) );
OR4_X1 _09101_ ( .A1(\myclint.mtime [48] ), .A2(_01544_ ), .A3(_01582_ ), .A4(_01551_ ), .ZN(_01584_ ) );
AOI21_X1 _09102_ ( .A(fanout_net_1 ), .B1(_01583_ ), .B2(_01584_ ), .ZN(_00007_ ) );
NAND3_X1 _09103_ ( .A1(_01512_ ), .A2(\myclint.mtime [44] ), .A3(_01513_ ), .ZN(_01585_ ) );
INV_X1 _09104_ ( .A(\myclint.mtime [45] ), .ZN(_01586_ ) );
NOR3_X1 _09105_ ( .A1(_01585_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01586_ ), .ZN(_01587_ ) );
AND2_X1 _09106_ ( .A1(_01587_ ), .A2(\myclint.mtime [47] ), .ZN(_01588_ ) );
NAND3_X1 _09107_ ( .A1(_01512_ ), .A2(_01515_ ), .A3(_01513_ ), .ZN(_01589_ ) );
NOR2_X1 _09108_ ( .A1(_01589_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01590_ ) );
OAI21_X1 _09109_ ( .A(_01536_ ), .B1(_01590_ ), .B2(\myclint.mtime [47] ), .ZN(_01591_ ) );
NOR2_X1 _09110_ ( .A1(_01588_ ), .A2(_01591_ ), .ZN(_00008_ ) );
AND2_X1 _09111_ ( .A1(_01554_ ), .A2(_01556_ ), .ZN(_01592_ ) );
AND2_X1 _09112_ ( .A1(_01552_ ), .A2(_01592_ ), .ZN(_01593_ ) );
AND3_X1 _09113_ ( .A1(_01593_ ), .A2(_01515_ ), .A3(_01555_ ), .ZN(_01594_ ) );
XNOR2_X1 _09114_ ( .A(_01594_ ), .B(\myclint.mtime [46] ), .ZN(_01595_ ) );
NOR2_X1 _09115_ ( .A1(_01595_ ), .A2(fanout_net_1 ), .ZN(_00009_ ) );
INV_X1 _09116_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01596_ ) );
AND3_X1 _09117_ ( .A1(_01512_ ), .A2(_01596_ ), .A3(_01513_ ), .ZN(_01597_ ) );
AND2_X1 _09118_ ( .A1(_01597_ ), .A2(\myclint.mtime [45] ), .ZN(_01598_ ) );
BUF_X4 _09119_ ( .A(_01535_ ), .Z(_01599_ ) );
OAI21_X1 _09120_ ( .A(_01599_ ), .B1(_01597_ ), .B2(\myclint.mtime [45] ), .ZN(_01600_ ) );
NOR2_X1 _09121_ ( .A1(_01598_ ), .A2(_01600_ ), .ZN(_00010_ ) );
AND2_X1 _09122_ ( .A1(_01593_ ), .A2(_01555_ ), .ZN(_01601_ ) );
XNOR2_X1 _09123_ ( .A(_01601_ ), .B(\myclint.mtime [44] ), .ZN(_01602_ ) );
NOR2_X1 _09124_ ( .A1(_01602_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
AND2_X1 _09125_ ( .A1(_01560_ ), .A2(_01561_ ), .ZN(_01603_ ) );
INV_X1 _09126_ ( .A(_01603_ ), .ZN(_01604_ ) );
OR3_X1 _09127_ ( .A1(_01604_ ), .A2(\myclint.mtime [61] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01605_ ) );
OAI21_X1 _09128_ ( .A(\myclint.mtime [61] ), .B1(_01604_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01606_ ) );
AOI21_X1 _09129_ ( .A(fanout_net_1 ), .B1(_01605_ ), .B2(_01606_ ), .ZN(_00012_ ) );
NAND3_X1 _09130_ ( .A1(_01552_ ), .A2(_01511_ ), .A3(_01592_ ), .ZN(_01607_ ) );
OR3_X1 _09131_ ( .A1(_01607_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [43] ), .ZN(_01608_ ) );
OAI21_X1 _09132_ ( .A(\myclint.mtime [43] ), .B1(_01607_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01609_ ) );
AOI21_X1 _09133_ ( .A(fanout_net_1 ), .B1(_01608_ ), .B2(_01609_ ), .ZN(_00013_ ) );
OR2_X1 _09134_ ( .A1(_01607_ ), .A2(\myclint.mtime [42] ), .ZN(_01610_ ) );
NAND2_X1 _09135_ ( .A1(_01607_ ), .A2(\myclint.mtime [42] ), .ZN(_01611_ ) );
AOI21_X1 _09136_ ( .A(fanout_net_1 ), .B1(_01610_ ), .B2(_01611_ ), .ZN(_00014_ ) );
INV_X1 _09137_ ( .A(_01593_ ), .ZN(_01612_ ) );
OR3_X1 _09138_ ( .A1(_01612_ ), .A2(\myclint.mtime [41] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01613_ ) );
OAI21_X1 _09139_ ( .A(\myclint.mtime [41] ), .B1(_01612_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01614_ ) );
AOI21_X1 _09140_ ( .A(fanout_net_1 ), .B1(_01613_ ), .B2(_01614_ ), .ZN(_00015_ ) );
XNOR2_X1 _09141_ ( .A(_01593_ ), .B(\myclint.mtime [40] ), .ZN(_01615_ ) );
NOR2_X1 _09142_ ( .A1(_01615_ ), .A2(fanout_net_1 ), .ZN(_00016_ ) );
INV_X1 _09143_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01616_ ) );
AND3_X1 _09144_ ( .A1(_01507_ ), .A2(_01616_ ), .A3(\myclint.mtime [37] ), .ZN(_01617_ ) );
AND2_X1 _09145_ ( .A1(_01617_ ), .A2(\myclint.mtime [39] ), .ZN(_01618_ ) );
OAI21_X1 _09146_ ( .A(_01599_ ), .B1(_01617_ ), .B2(\myclint.mtime [39] ), .ZN(_01619_ ) );
NOR2_X1 _09147_ ( .A1(_01618_ ), .A2(_01619_ ), .ZN(_00017_ ) );
AND2_X1 _09148_ ( .A1(_01552_ ), .A2(_01554_ ), .ZN(_01620_ ) );
NAND3_X1 _09149_ ( .A1(_01620_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .ZN(_01621_ ) );
OR2_X1 _09150_ ( .A1(_01621_ ), .A2(\myclint.mtime [38] ), .ZN(_01622_ ) );
NAND2_X1 _09151_ ( .A1(_01621_ ), .A2(\myclint.mtime [38] ), .ZN(_01623_ ) );
AOI21_X1 _09152_ ( .A(fanout_net_1 ), .B1(_01622_ ), .B2(_01623_ ), .ZN(_00018_ ) );
BUF_X4 _09153_ ( .A(_01535_ ), .Z(_01624_ ) );
INV_X1 _09154_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01625_ ) );
AND3_X1 _09155_ ( .A1(_01506_ ), .A2(_01625_ ), .A3(\myclint.mtime [35] ), .ZN(_01626_ ) );
OAI21_X1 _09156_ ( .A(_01624_ ), .B1(_01626_ ), .B2(\myclint.mtime [37] ), .ZN(_01627_ ) );
NAND4_X1 _09157_ ( .A1(_01502_ ), .A2(\myclint.mtime [33] ), .A3(_01503_ ), .A4(_01504_ ), .ZN(_01628_ ) );
INV_X1 _09158_ ( .A(\myclint.mtime [32] ), .ZN(_01629_ ) );
NOR2_X1 _09159_ ( .A1(_01628_ ), .A2(_01629_ ), .ZN(_01630_ ) );
AND3_X1 _09160_ ( .A1(_01630_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01631_ ) );
AND3_X1 _09161_ ( .A1(_01631_ ), .A2(\myclint.mtime [37] ), .A3(_01625_ ), .ZN(_01632_ ) );
NOR2_X1 _09162_ ( .A1(_01627_ ), .A2(_01632_ ), .ZN(_00019_ ) );
OAI21_X1 _09163_ ( .A(_01624_ ), .B1(_01631_ ), .B2(\myclint.mtime [36] ), .ZN(_01633_ ) );
NOR2_X1 _09164_ ( .A1(_01633_ ), .A2(_01507_ ), .ZN(_00020_ ) );
NOR3_X1 _09165_ ( .A1(_01628_ ), .A2(_01629_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01634_ ) );
OAI21_X1 _09166_ ( .A(_01624_ ), .B1(_01634_ ), .B2(\myclint.mtime [35] ), .ZN(_01635_ ) );
INV_X1 _09167_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01636_ ) );
AND3_X1 _09168_ ( .A1(_01630_ ), .A2(_01636_ ), .A3(\myclint.mtime [35] ), .ZN(_01637_ ) );
NOR2_X1 _09169_ ( .A1(_01635_ ), .A2(_01637_ ), .ZN(_00021_ ) );
OAI21_X1 _09170_ ( .A(_01624_ ), .B1(_01630_ ), .B2(\myclint.mtime [34] ), .ZN(_01638_ ) );
NOR2_X1 _09171_ ( .A1(_01638_ ), .A2(_01506_ ), .ZN(_00022_ ) );
XNOR2_X1 _09172_ ( .A(_01603_ ), .B(\myclint.mtime [60] ), .ZN(_01639_ ) );
NOR2_X1 _09173_ ( .A1(_01639_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
AND2_X1 _09174_ ( .A1(_01502_ ), .A2(_01504_ ), .ZN(_01640_ ) );
INV_X1 _09175_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01641_ ) );
AND3_X1 _09176_ ( .A1(_01640_ ), .A2(_01641_ ), .A3(_01503_ ), .ZN(_01642_ ) );
AND2_X1 _09177_ ( .A1(_01642_ ), .A2(\myclint.mtime [33] ), .ZN(_01643_ ) );
OAI21_X1 _09178_ ( .A(_01599_ ), .B1(_01642_ ), .B2(\myclint.mtime [33] ), .ZN(_01644_ ) );
NOR2_X1 _09179_ ( .A1(_01643_ ), .A2(_01644_ ), .ZN(_00024_ ) );
AND4_X1 _09180_ ( .A1(_01503_ ), .A2(_01541_ ), .A3(_01504_ ), .A4(_01543_ ), .ZN(_01645_ ) );
AND2_X1 _09181_ ( .A1(_01547_ ), .A2(_01550_ ), .ZN(_01646_ ) );
NAND3_X1 _09182_ ( .A1(_01645_ ), .A2(_01629_ ), .A3(_01646_ ), .ZN(_01647_ ) );
OAI21_X1 _09183_ ( .A(\myclint.mtime [32] ), .B1(_01544_ ), .B2(_01551_ ), .ZN(_01648_ ) );
AOI21_X1 _09184_ ( .A(fanout_net_1 ), .B1(_01647_ ), .B2(_01648_ ), .ZN(_00025_ ) );
INV_X1 _09185_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01649_ ) );
AND3_X1 _09186_ ( .A1(_01502_ ), .A2(_01649_ ), .A3(_01504_ ), .ZN(_01650_ ) );
AND2_X1 _09187_ ( .A1(_01650_ ), .A2(\myclint.mtime [31] ), .ZN(_01651_ ) );
OAI21_X1 _09188_ ( .A(_01599_ ), .B1(_01650_ ), .B2(\myclint.mtime [31] ), .ZN(_01652_ ) );
NOR2_X1 _09189_ ( .A1(_01651_ ), .A2(_01652_ ), .ZN(_00026_ ) );
AND2_X1 _09190_ ( .A1(_01646_ ), .A2(_01541_ ), .ZN(_01653_ ) );
NAND3_X1 _09191_ ( .A1(_01653_ ), .A2(_01504_ ), .A3(_01543_ ), .ZN(_01654_ ) );
OR2_X1 _09192_ ( .A1(_01654_ ), .A2(\myclint.mtime [30] ), .ZN(_01655_ ) );
NAND2_X1 _09193_ ( .A1(_01654_ ), .A2(\myclint.mtime [30] ), .ZN(_01656_ ) );
AOI21_X1 _09194_ ( .A(fanout_net_1 ), .B1(_01655_ ), .B2(_01656_ ), .ZN(_00027_ ) );
INV_X1 _09195_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01657_ ) );
AND3_X1 _09196_ ( .A1(_01501_ ), .A2(_01657_ ), .A3(\myclint.mtime [27] ), .ZN(_01658_ ) );
AND2_X1 _09197_ ( .A1(_01658_ ), .A2(\myclint.mtime [29] ), .ZN(_01659_ ) );
OAI21_X1 _09198_ ( .A(_01599_ ), .B1(_01658_ ), .B2(\myclint.mtime [29] ), .ZN(_01660_ ) );
NOR2_X1 _09199_ ( .A1(_01659_ ), .A2(_01660_ ), .ZN(_00028_ ) );
NAND2_X1 _09200_ ( .A1(_01653_ ), .A2(_01543_ ), .ZN(_01661_ ) );
OR2_X1 _09201_ ( .A1(_01661_ ), .A2(\myclint.mtime [28] ), .ZN(_01662_ ) );
NAND2_X1 _09202_ ( .A1(_01661_ ), .A2(\myclint.mtime [28] ), .ZN(_01663_ ) );
AOI21_X1 _09203_ ( .A(fanout_net_1 ), .B1(_01662_ ), .B2(_01663_ ), .ZN(_00029_ ) );
NAND3_X1 _09204_ ( .A1(_01646_ ), .A2(_01542_ ), .A3(_01541_ ), .ZN(_01664_ ) );
OR3_X1 _09205_ ( .A1(_01664_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01665_ ) );
OAI21_X1 _09206_ ( .A(\myclint.mtime [27] ), .B1(_01664_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01666_ ) );
AOI21_X1 _09207_ ( .A(fanout_net_1 ), .B1(_01665_ ), .B2(_01666_ ), .ZN(_00030_ ) );
AND2_X1 _09208_ ( .A1(_01500_ ), .A2(\myclint.mtime [25] ), .ZN(_01667_ ) );
OAI21_X1 _09209_ ( .A(_01624_ ), .B1(_01667_ ), .B2(\myclint.mtime [26] ), .ZN(_01668_ ) );
NOR2_X1 _09210_ ( .A1(_01668_ ), .A2(_01501_ ), .ZN(_00031_ ) );
INV_X1 _09211_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01669_ ) );
AND3_X1 _09212_ ( .A1(_01499_ ), .A2(_01669_ ), .A3(\myclint.mtime [23] ), .ZN(_01670_ ) );
AND2_X1 _09213_ ( .A1(_01670_ ), .A2(\myclint.mtime [25] ), .ZN(_01671_ ) );
OAI21_X1 _09214_ ( .A(_01599_ ), .B1(_01670_ ), .B2(\myclint.mtime [25] ), .ZN(_01672_ ) );
NOR2_X1 _09215_ ( .A1(_01671_ ), .A2(_01672_ ), .ZN(_00032_ ) );
AND2_X1 _09216_ ( .A1(_01499_ ), .A2(\myclint.mtime [23] ), .ZN(_01673_ ) );
OAI21_X1 _09217_ ( .A(_01624_ ), .B1(_01673_ ), .B2(\myclint.mtime [24] ), .ZN(_01674_ ) );
NOR2_X1 _09218_ ( .A1(_01674_ ), .A2(_01500_ ), .ZN(_00033_ ) );
NAND3_X1 _09219_ ( .A1(_01558_ ), .A2(_01526_ ), .A3(_01559_ ), .ZN(_01675_ ) );
OR3_X1 _09220_ ( .A1(_01675_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [59] ), .ZN(_01676_ ) );
OAI21_X1 _09221_ ( .A(\myclint.mtime [59] ), .B1(_01675_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01677_ ) );
AOI21_X1 _09222_ ( .A(fanout_net_1 ), .B1(_01676_ ), .B2(_01677_ ), .ZN(_00034_ ) );
AND2_X1 _09223_ ( .A1(_01646_ ), .A2(_01539_ ), .ZN(_01678_ ) );
NAND3_X1 _09224_ ( .A1(_01678_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01679_ ) );
OR3_X1 _09225_ ( .A1(_01679_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01680_ ) );
OAI21_X1 _09226_ ( .A(\myclint.mtime [23] ), .B1(_01679_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01681_ ) );
AOI21_X1 _09227_ ( .A(fanout_net_1 ), .B1(_01680_ ), .B2(_01681_ ), .ZN(_00035_ ) );
AND2_X1 _09228_ ( .A1(_01498_ ), .A2(\myclint.mtime [21] ), .ZN(_01682_ ) );
OAI21_X1 _09229_ ( .A(_01624_ ), .B1(_01682_ ), .B2(\myclint.mtime [22] ), .ZN(_01683_ ) );
NOR2_X1 _09230_ ( .A1(_01683_ ), .A2(_01499_ ), .ZN(_00036_ ) );
INV_X1 _09231_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01684_ ) );
AND3_X1 _09232_ ( .A1(_01497_ ), .A2(_01684_ ), .A3(\myclint.mtime [19] ), .ZN(_01685_ ) );
AND2_X1 _09233_ ( .A1(_01685_ ), .A2(\myclint.mtime [21] ), .ZN(_01686_ ) );
OAI21_X1 _09234_ ( .A(_01599_ ), .B1(_01685_ ), .B2(\myclint.mtime [21] ), .ZN(_01687_ ) );
NOR2_X1 _09235_ ( .A1(_01686_ ), .A2(_01687_ ), .ZN(_00037_ ) );
AND2_X1 _09236_ ( .A1(_01497_ ), .A2(\myclint.mtime [19] ), .ZN(_01688_ ) );
OAI21_X1 _09237_ ( .A(_01624_ ), .B1(_01688_ ), .B2(\myclint.mtime [20] ), .ZN(_01689_ ) );
NOR2_X1 _09238_ ( .A1(_01689_ ), .A2(_01498_ ), .ZN(_00038_ ) );
NAND3_X1 _09239_ ( .A1(_01646_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01690_ ) );
OR3_X1 _09240_ ( .A1(_01690_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01691_ ) );
OAI21_X1 _09241_ ( .A(\myclint.mtime [19] ), .B1(_01690_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01692_ ) );
AOI21_X1 _09242_ ( .A(fanout_net_1 ), .B1(_01691_ ), .B2(_01692_ ), .ZN(_00039_ ) );
AND2_X1 _09243_ ( .A1(_01496_ ), .A2(\myclint.mtime [17] ), .ZN(_01693_ ) );
OAI21_X1 _09244_ ( .A(_01624_ ), .B1(_01693_ ), .B2(\myclint.mtime [18] ), .ZN(_01694_ ) );
NOR2_X1 _09245_ ( .A1(_01694_ ), .A2(_01497_ ), .ZN(_00040_ ) );
INV_X1 _09246_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01695_ ) );
AND3_X1 _09247_ ( .A1(_01495_ ), .A2(_01695_ ), .A3(\myclint.mtime [15] ), .ZN(_01696_ ) );
AND2_X1 _09248_ ( .A1(_01696_ ), .A2(\myclint.mtime [17] ), .ZN(_01697_ ) );
OAI21_X1 _09249_ ( .A(_01599_ ), .B1(_01696_ ), .B2(\myclint.mtime [17] ), .ZN(_01698_ ) );
NOR2_X1 _09250_ ( .A1(_01697_ ), .A2(_01698_ ), .ZN(_00041_ ) );
AND2_X1 _09251_ ( .A1(_01495_ ), .A2(\myclint.mtime [15] ), .ZN(_01699_ ) );
OAI21_X1 _09252_ ( .A(_01536_ ), .B1(_01699_ ), .B2(\myclint.mtime [16] ), .ZN(_01700_ ) );
NOR2_X1 _09253_ ( .A1(_01700_ ), .A2(_01496_ ), .ZN(_00042_ ) );
AND3_X1 _09254_ ( .A1(_01549_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [11] ), .ZN(_01701_ ) );
AND2_X1 _09255_ ( .A1(_01547_ ), .A2(_01701_ ), .ZN(_01702_ ) );
NAND3_X1 _09256_ ( .A1(_01702_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01703_ ) );
OR3_X1 _09257_ ( .A1(_01703_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01704_ ) );
OAI21_X1 _09258_ ( .A(\myclint.mtime [15] ), .B1(_01703_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01705_ ) );
AOI21_X1 _09259_ ( .A(fanout_net_1 ), .B1(_01704_ ), .B2(_01705_ ), .ZN(_00043_ ) );
AND2_X1 _09260_ ( .A1(_01494_ ), .A2(\myclint.mtime [13] ), .ZN(_01706_ ) );
OAI21_X1 _09261_ ( .A(_01536_ ), .B1(_01706_ ), .B2(\myclint.mtime [14] ), .ZN(_01707_ ) );
NOR2_X1 _09262_ ( .A1(_01707_ ), .A2(_01495_ ), .ZN(_00044_ ) );
OR2_X1 _09263_ ( .A1(_01675_ ), .A2(\myclint.mtime [58] ), .ZN(_01708_ ) );
NAND2_X1 _09264_ ( .A1(_01675_ ), .A2(\myclint.mtime [58] ), .ZN(_01709_ ) );
AOI21_X1 _09265_ ( .A(fanout_net_1 ), .B1(_01708_ ), .B2(_01709_ ), .ZN(_00045_ ) );
INV_X1 _09266_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01710_ ) );
AND3_X1 _09267_ ( .A1(_01493_ ), .A2(_01710_ ), .A3(\myclint.mtime [11] ), .ZN(_01711_ ) );
AND2_X1 _09268_ ( .A1(_01711_ ), .A2(\myclint.mtime [13] ), .ZN(_01712_ ) );
OAI21_X1 _09269_ ( .A(_01599_ ), .B1(_01711_ ), .B2(\myclint.mtime [13] ), .ZN(_01713_ ) );
NOR2_X1 _09270_ ( .A1(_01712_ ), .A2(_01713_ ), .ZN(_00046_ ) );
AND2_X1 _09271_ ( .A1(_01493_ ), .A2(\myclint.mtime [11] ), .ZN(_01714_ ) );
OAI21_X1 _09272_ ( .A(_01536_ ), .B1(_01714_ ), .B2(\myclint.mtime [12] ), .ZN(_01715_ ) );
NOR2_X1 _09273_ ( .A1(_01715_ ), .A2(_01494_ ), .ZN(_00047_ ) );
NAND3_X1 _09274_ ( .A1(_01545_ ), .A2(_01546_ ), .A3(_01549_ ), .ZN(_01716_ ) );
OR3_X1 _09275_ ( .A1(_01716_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_01717_ ) );
OAI21_X1 _09276_ ( .A(\myclint.mtime [11] ), .B1(_01716_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01718_ ) );
AOI21_X1 _09277_ ( .A(fanout_net_1 ), .B1(_01717_ ), .B2(_01718_ ), .ZN(_00048_ ) );
OR2_X1 _09278_ ( .A1(_01716_ ), .A2(\myclint.mtime [10] ), .ZN(_01719_ ) );
NAND2_X1 _09279_ ( .A1(_01716_ ), .A2(\myclint.mtime [10] ), .ZN(_01720_ ) );
AOI21_X1 _09280_ ( .A(fanout_net_1 ), .B1(_01719_ ), .B2(_01720_ ), .ZN(_00049_ ) );
AND2_X1 _09281_ ( .A1(_01491_ ), .A2(\myclint.mtime [7] ), .ZN(_01721_ ) );
INV_X1 _09282_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01722_ ) );
AND3_X1 _09283_ ( .A1(_01721_ ), .A2(\myclint.mtime [9] ), .A3(_01722_ ), .ZN(_01723_ ) );
AOI21_X1 _09284_ ( .A(\myclint.mtime [9] ), .B1(_01721_ ), .B2(_01722_ ), .ZN(_01724_ ) );
NOR3_X1 _09285_ ( .A1(_01723_ ), .A2(_01724_ ), .A3(fanout_net_1 ), .ZN(_00050_ ) );
OAI21_X1 _09286_ ( .A(_01536_ ), .B1(_01721_ ), .B2(\myclint.mtime [8] ), .ZN(_01725_ ) );
NOR2_X1 _09287_ ( .A1(_01725_ ), .A2(_01492_ ), .ZN(_00051_ ) );
AND2_X1 _09288_ ( .A1(_01490_ ), .A2(\myclint.mtime [5] ), .ZN(_01726_ ) );
INV_X1 _09289_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01727_ ) );
AND3_X1 _09290_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(\myclint.mtime [7] ), .ZN(_01728_ ) );
AOI21_X1 _09291_ ( .A(\myclint.mtime [7] ), .B1(_01726_ ), .B2(_01727_ ), .ZN(_01729_ ) );
NOR3_X1 _09292_ ( .A1(_01728_ ), .A2(_01729_ ), .A3(fanout_net_1 ), .ZN(_00052_ ) );
OAI21_X1 _09293_ ( .A(_01536_ ), .B1(_01726_ ), .B2(\myclint.mtime [6] ), .ZN(_01730_ ) );
NOR2_X1 _09294_ ( .A1(_01730_ ), .A2(_01491_ ), .ZN(_00053_ ) );
INV_X1 _09295_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01731_ ) );
AND3_X1 _09296_ ( .A1(_01545_ ), .A2(\myclint.mtime [5] ), .A3(_01731_ ), .ZN(_01732_ ) );
AOI21_X1 _09297_ ( .A(\myclint.mtime [5] ), .B1(_01545_ ), .B2(_01731_ ), .ZN(_01733_ ) );
NOR3_X1 _09298_ ( .A1(_01732_ ), .A2(_01733_ ), .A3(fanout_net_1 ), .ZN(_00054_ ) );
OAI21_X1 _09299_ ( .A(_01536_ ), .B1(_01545_ ), .B2(\myclint.mtime [4] ), .ZN(_01734_ ) );
NOR2_X1 _09300_ ( .A1(_01734_ ), .A2(_01490_ ), .ZN(_00055_ ) );
INV_X1 _09301_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01735_ ) );
AND3_X1 _09302_ ( .A1(_01523_ ), .A2(_01735_ ), .A3(_01524_ ), .ZN(_01736_ ) );
AND2_X1 _09303_ ( .A1(_01736_ ), .A2(\myclint.mtime [57] ), .ZN(_01737_ ) );
OAI21_X1 _09304_ ( .A(_01599_ ), .B1(_01736_ ), .B2(\myclint.mtime [57] ), .ZN(_01738_ ) );
NOR2_X1 _09305_ ( .A1(_01737_ ), .A2(_01738_ ), .ZN(_00056_ ) );
AND2_X1 _09306_ ( .A1(\myclint.mtime [1] ), .A2(\myclint.mtime [0] ), .ZN(_01739_ ) );
INV_X1 _09307_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01740_ ) );
AND3_X1 _09308_ ( .A1(_01739_ ), .A2(_01740_ ), .A3(\myclint.mtime [3] ), .ZN(_01741_ ) );
AOI21_X1 _09309_ ( .A(\myclint.mtime [3] ), .B1(_01739_ ), .B2(_01740_ ), .ZN(_01742_ ) );
NOR3_X1 _09310_ ( .A1(_01741_ ), .A2(_01742_ ), .A3(fanout_net_1 ), .ZN(_00057_ ) );
AOI21_X1 _09311_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [1] ), .B2(\myclint.mtime [0] ), .ZN(_01743_ ) );
NOR3_X1 _09312_ ( .A1(_01489_ ), .A2(_01743_ ), .A3(fanout_net_2 ), .ZN(_00058_ ) );
NOR2_X1 _09313_ ( .A1(\myclint.mtime [1] ), .A2(\myclint.mtime [0] ), .ZN(_01744_ ) );
NOR3_X1 _09314_ ( .A1(_01739_ ), .A2(_01744_ ), .A3(fanout_net_2 ), .ZN(_00059_ ) );
INV_X1 _09315_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_01745_ ) );
NOR2_X1 _09316_ ( .A1(_01745_ ), .A2(fanout_net_2 ), .ZN(_00060_ ) );
INV_X1 _09317_ ( .A(_01560_ ), .ZN(_01746_ ) );
OR2_X1 _09318_ ( .A1(_01746_ ), .A2(\myclint.mtime [56] ), .ZN(_01747_ ) );
NAND2_X1 _09319_ ( .A1(_01746_ ), .A2(\myclint.mtime [56] ), .ZN(_01748_ ) );
AOI21_X1 _09320_ ( .A(fanout_net_2 ), .B1(_01747_ ), .B2(_01748_ ), .ZN(_00061_ ) );
NAND3_X1 _09321_ ( .A1(_01558_ ), .A2(_01522_ ), .A3(_01565_ ), .ZN(_01749_ ) );
OR3_X1 _09322_ ( .A1(_01749_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01750_ ) );
OAI21_X1 _09323_ ( .A(\myclint.mtime [55] ), .B1(_01749_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01751_ ) );
AOI21_X1 _09324_ ( .A(fanout_net_2 ), .B1(_01750_ ), .B2(_01751_ ), .ZN(_00062_ ) );
OR2_X1 _09325_ ( .A1(_01749_ ), .A2(\myclint.mtime [54] ), .ZN(_01752_ ) );
NAND2_X1 _09326_ ( .A1(_01749_ ), .A2(\myclint.mtime [54] ), .ZN(_01753_ ) );
AOI21_X1 _09327_ ( .A(fanout_net_2 ), .B1(_01752_ ), .B2(_01753_ ), .ZN(_00063_ ) );
MUX2_X1 _09328_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(fanout_net_40 ), .Z(_01754_ ) );
MUX2_X1 _09329_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_40 ), .Z(_01755_ ) );
MUX2_X1 _09330_ ( .A(_01754_ ), .B(_01755_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01756_ ) );
INV_X1 _09331_ ( .A(\IF_ID_pc [25] ), .ZN(_01757_ ) );
NAND2_X1 _09332_ ( .A1(_01756_ ), .A2(_01757_ ), .ZN(_01758_ ) );
INV_X1 _09333_ ( .A(\IF_ID_pc [24] ), .ZN(_01759_ ) );
INV_X32 _09334_ ( .A(fanout_net_40 ), .ZN(_01760_ ) );
CLKBUF_X2 _09335_ ( .A(_01760_ ), .Z(_01761_ ) );
OR2_X1 _09336_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[1][19] ), .ZN(_01762_ ) );
INV_X32 _09337_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01763_ ) );
BUF_X4 _09338_ ( .A(_01763_ ), .Z(_01764_ ) );
BUF_X4 _09339_ ( .A(_01764_ ), .Z(_01765_ ) );
OAI211_X1 _09340_ ( .A(_01762_ ), .B(_01765_ ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[0][19] ), .ZN(_01766_ ) );
OR2_X1 _09341_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][19] ), .ZN(_01767_ ) );
OAI211_X1 _09342_ ( .A(_01767_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01761_ ), .C2(\myifu.myicache.tag[3][19] ), .ZN(_01768_ ) );
NAND2_X1 _09343_ ( .A1(_01766_ ), .A2(_01768_ ), .ZN(_01769_ ) );
OR2_X1 _09344_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[1][14] ), .ZN(_01770_ ) );
OAI211_X1 _09345_ ( .A(_01770_ ), .B(_01765_ ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[0][14] ), .ZN(_01771_ ) );
INV_X1 _09346_ ( .A(\IF_ID_pc [19] ), .ZN(_01772_ ) );
OR2_X1 _09347_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][14] ), .ZN(_01773_ ) );
OAI211_X1 _09348_ ( .A(_01773_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01761_ ), .C2(\myifu.myicache.tag[3][14] ), .ZN(_01774_ ) );
AND3_X1 _09349_ ( .A1(_01771_ ), .A2(_01772_ ), .A3(_01774_ ), .ZN(_01775_ ) );
AOI21_X1 _09350_ ( .A(_01772_ ), .B1(_01771_ ), .B2(_01774_ ), .ZN(_01776_ ) );
OAI221_X1 _09351_ ( .A(_01758_ ), .B1(_01759_ ), .B2(_01769_ ), .C1(_01775_ ), .C2(_01776_ ), .ZN(_01777_ ) );
OR2_X1 _09352_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_01778_ ) );
OAI211_X1 _09353_ ( .A(_01778_ ), .B(_01765_ ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_01779_ ) );
OR2_X1 _09354_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[3][6] ), .ZN(_01780_ ) );
OAI211_X1 _09355_ ( .A(_01780_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[2][6] ), .ZN(_01781_ ) );
INV_X1 _09356_ ( .A(\IF_ID_pc [11] ), .ZN(_01782_ ) );
AND3_X1 _09357_ ( .A1(_01779_ ), .A2(_01781_ ), .A3(_01782_ ), .ZN(_01783_ ) );
AOI21_X1 _09358_ ( .A(_01782_ ), .B1(_01779_ ), .B2(_01781_ ), .ZN(_01784_ ) );
OR2_X2 _09359_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[1][23] ), .ZN(_01785_ ) );
OAI211_X1 _09360_ ( .A(_01785_ ), .B(_01765_ ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[0][23] ), .ZN(_01786_ ) );
INV_X1 _09361_ ( .A(\IF_ID_pc [28] ), .ZN(_01787_ ) );
OR2_X1 _09362_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][23] ), .ZN(_01788_ ) );
OAI211_X1 _09363_ ( .A(_01788_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01761_ ), .C2(\myifu.myicache.tag[3][23] ), .ZN(_01789_ ) );
AND3_X1 _09364_ ( .A1(_01786_ ), .A2(_01787_ ), .A3(_01789_ ), .ZN(_01790_ ) );
AOI21_X1 _09365_ ( .A(_01787_ ), .B1(_01786_ ), .B2(_01789_ ), .ZN(_01791_ ) );
OAI22_X1 _09366_ ( .A1(_01783_ ), .A2(_01784_ ), .B1(_01790_ ), .B2(_01791_ ), .ZN(_01792_ ) );
NOR2_X1 _09367_ ( .A1(_01777_ ), .A2(_01792_ ), .ZN(_01793_ ) );
MUX2_X1 _09368_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(fanout_net_40 ), .Z(_01794_ ) );
MUX2_X1 _09369_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(fanout_net_40 ), .Z(_01795_ ) );
MUX2_X2 _09370_ ( .A(_01794_ ), .B(_01795_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01796_ ) );
INV_X1 _09371_ ( .A(\IF_ID_pc [20] ), .ZN(_01797_ ) );
XNOR2_X1 _09372_ ( .A(_01796_ ), .B(_01797_ ), .ZN(_01798_ ) );
MUX2_X1 _09373_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(fanout_net_40 ), .Z(_01799_ ) );
OR2_X2 _09374_ ( .A1(_01799_ ), .A2(_01763_ ), .ZN(_01800_ ) );
MUX2_X2 _09375_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(fanout_net_40 ), .Z(_01801_ ) );
OAI21_X4 _09376_ ( .A(_01800_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01801_ ), .ZN(_01802_ ) );
INV_X1 _09377_ ( .A(\IF_ID_pc [8] ), .ZN(_01803_ ) );
MUX2_X1 _09378_ ( .A(\myifu.myicache.tag[0][3] ), .B(\myifu.myicache.tag[1][3] ), .S(fanout_net_40 ), .Z(_01804_ ) );
MUX2_X1 _09379_ ( .A(\myifu.myicache.tag[2][3] ), .B(\myifu.myicache.tag[3][3] ), .S(fanout_net_40 ), .Z(_01805_ ) );
MUX2_X2 _09380_ ( .A(_01804_ ), .B(_01805_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01806_ ) );
AOI221_X1 _09381_ ( .A(_01798_ ), .B1(\IF_ID_pc [12] ), .B2(_01802_ ), .C1(_01803_ ), .C2(_01806_ ), .ZN(_01807_ ) );
MUX2_X1 _09382_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(fanout_net_40 ), .Z(_01808_ ) );
AND2_X2 _09383_ ( .A1(_01808_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01809_ ) );
MUX2_X1 _09384_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(fanout_net_40 ), .Z(_01810_ ) );
AOI21_X4 _09385_ ( .A(_01809_ ), .B1(_01764_ ), .B2(_01810_ ), .ZN(_01811_ ) );
OAI22_X2 _09386_ ( .A1(_01811_ ), .A2(\IF_ID_pc [21] ), .B1(_01802_ ), .B2(\IF_ID_pc [12] ), .ZN(_01812_ ) );
MUX2_X1 _09387_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(fanout_net_40 ), .Z(_01813_ ) );
OR2_X2 _09388_ ( .A1(_01813_ ), .A2(_01764_ ), .ZN(_01814_ ) );
MUX2_X1 _09389_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(fanout_net_40 ), .Z(_01815_ ) );
OAI21_X1 _09390_ ( .A(_01814_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01815_ ), .ZN(_01816_ ) );
MUX2_X1 _09391_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(fanout_net_40 ), .Z(_01817_ ) );
OR2_X1 _09392_ ( .A1(_01817_ ), .A2(_01764_ ), .ZN(_01818_ ) );
MUX2_X1 _09393_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(fanout_net_40 ), .Z(_01819_ ) );
OAI21_X1 _09394_ ( .A(_01818_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01819_ ), .ZN(_01820_ ) );
AOI221_X2 _09395_ ( .A(_01812_ ), .B1(\IF_ID_pc [27] ), .B2(_01816_ ), .C1(\IF_ID_pc [23] ), .C2(_01820_ ), .ZN(_01821_ ) );
AND2_X2 _09396_ ( .A1(_01807_ ), .A2(_01821_ ), .ZN(_01822_ ) );
MUX2_X1 _09397_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(fanout_net_40 ), .Z(_01823_ ) );
OR2_X2 _09398_ ( .A1(_01823_ ), .A2(_01764_ ), .ZN(_01824_ ) );
MUX2_X1 _09399_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(fanout_net_40 ), .Z(_01825_ ) );
OAI21_X2 _09400_ ( .A(_01824_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01825_ ), .ZN(_01826_ ) );
NOR2_X1 _09401_ ( .A1(_01826_ ), .A2(\IF_ID_pc [18] ), .ZN(_01827_ ) );
OAI22_X1 _09402_ ( .A1(_01757_ ), .A2(_01756_ ), .B1(_01806_ ), .B2(_01803_ ), .ZN(_01828_ ) );
MUX2_X1 _09403_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_40 ), .Z(_01829_ ) );
OR2_X1 _09404_ ( .A1(_01829_ ), .A2(_01764_ ), .ZN(_01830_ ) );
MUX2_X1 _09405_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_40 ), .Z(_01831_ ) );
OAI21_X1 _09406_ ( .A(_01830_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01831_ ), .ZN(_01832_ ) );
AOI211_X2 _09407_ ( .A(_01827_ ), .B(_01828_ ), .C1(\IF_ID_pc [16] ), .C2(_01832_ ), .ZN(_01833_ ) );
MUX2_X1 _09408_ ( .A(\myifu.myicache.tag[0][26] ), .B(\myifu.myicache.tag[1][26] ), .S(fanout_net_40 ), .Z(_01834_ ) );
MUX2_X1 _09409_ ( .A(\myifu.myicache.tag[2][26] ), .B(\myifu.myicache.tag[3][26] ), .S(fanout_net_40 ), .Z(_01835_ ) );
MUX2_X1 _09410_ ( .A(_01834_ ), .B(_01835_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01836_ ) );
INV_X1 _09411_ ( .A(\IF_ID_pc [31] ), .ZN(_01837_ ) );
NOR2_X1 _09412_ ( .A1(_01836_ ), .A2(_01837_ ), .ZN(_01838_ ) );
AOI21_X1 _09413_ ( .A(_01838_ ), .B1(\IF_ID_pc [21] ), .B2(_01811_ ), .ZN(_01839_ ) );
MUX2_X1 _09414_ ( .A(\myifu.myicache.tag[2][0] ), .B(\myifu.myicache.tag[3][0] ), .S(fanout_net_40 ), .Z(_01840_ ) );
OR2_X1 _09415_ ( .A1(_01840_ ), .A2(_01764_ ), .ZN(_01841_ ) );
MUX2_X1 _09416_ ( .A(\myifu.myicache.tag[0][0] ), .B(\myifu.myicache.tag[1][0] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01842_ ) );
OR2_X1 _09417_ ( .A1(_01842_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01843_ ) );
AOI21_X1 _09418_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_01841_ ), .B2(_01843_ ), .ZN(_01844_ ) );
AOI21_X1 _09419_ ( .A(_01844_ ), .B1(_01837_ ), .B2(_01836_ ), .ZN(_01845_ ) );
AND4_X4 _09420_ ( .A1(_01822_ ), .A2(_01833_ ), .A3(_01839_ ), .A4(_01845_ ), .ZN(_01846_ ) );
AND2_X1 _09421_ ( .A1(_01826_ ), .A2(\IF_ID_pc [18] ), .ZN(_01847_ ) );
MUX2_X1 _09422_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01848_ ) );
MUX2_X1 _09423_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01849_ ) );
MUX2_X1 _09424_ ( .A(_01848_ ), .B(_01849_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01850_ ) );
INV_X1 _09425_ ( .A(_01850_ ), .ZN(_01851_ ) );
INV_X1 _09426_ ( .A(\IF_ID_pc [7] ), .ZN(_01852_ ) );
CLKBUF_X2 _09427_ ( .A(_01760_ ), .Z(_01853_ ) );
OR2_X1 _09428_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[1][2] ), .ZN(_01854_ ) );
OAI211_X1 _09429_ ( .A(_01854_ ), .B(_01765_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][2] ), .ZN(_01855_ ) );
OR2_X1 _09430_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[3][2] ), .ZN(_01856_ ) );
OAI211_X1 _09431_ ( .A(_01856_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][2] ), .ZN(_01857_ ) );
NAND2_X1 _09432_ ( .A1(_01855_ ), .A2(_01857_ ), .ZN(_01858_ ) );
AOI221_X4 _09433_ ( .A(_01847_ ), .B1(\IF_ID_pc [10] ), .B2(_01851_ ), .C1(_01852_ ), .C2(_01858_ ), .ZN(_01859_ ) );
AND3_X1 _09434_ ( .A1(_01855_ ), .A2(_01857_ ), .A3(\IF_ID_pc [7] ), .ZN(_01860_ ) );
OR2_X2 _09435_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_01861_ ) );
OAI211_X1 _09436_ ( .A(_01861_ ), .B(_01765_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_01862_ ) );
OR2_X1 _09437_ ( .A1(_01760_ ), .A2(\myifu.myicache.tag[3][25] ), .ZN(_01863_ ) );
OAI211_X1 _09438_ ( .A(_01863_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][25] ), .ZN(_01864_ ) );
NAND2_X1 _09439_ ( .A1(_01862_ ), .A2(_01864_ ), .ZN(_01865_ ) );
INV_X1 _09440_ ( .A(\IF_ID_pc [30] ), .ZN(_01866_ ) );
XNOR2_X1 _09441_ ( .A(_01865_ ), .B(_01866_ ), .ZN(_01867_ ) );
AOI211_X1 _09442_ ( .A(_01860_ ), .B(_01867_ ), .C1(_01759_ ), .C2(_01769_ ), .ZN(_01868_ ) );
AND4_X4 _09443_ ( .A1(_01793_ ), .A2(_01846_ ), .A3(_01859_ ), .A4(_01868_ ), .ZN(_01869_ ) );
OR2_X1 _09444_ ( .A1(_01760_ ), .A2(\myifu.myicache.tag[1][9] ), .ZN(_01870_ ) );
OAI211_X1 _09445_ ( .A(_01870_ ), .B(_01764_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][9] ), .ZN(_01871_ ) );
OR2_X1 _09446_ ( .A1(_01760_ ), .A2(\myifu.myicache.tag[3][9] ), .ZN(_01872_ ) );
OAI211_X1 _09447_ ( .A(_01872_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][9] ), .ZN(_01873_ ) );
AND3_X1 _09448_ ( .A1(_01871_ ), .A2(_01873_ ), .A3(\IF_ID_pc [14] ), .ZN(_01874_ ) );
INV_X1 _09449_ ( .A(\IF_ID_pc [29] ), .ZN(_01875_ ) );
MUX2_X1 _09450_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01876_ ) );
MUX2_X1 _09451_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01877_ ) );
MUX2_X1 _09452_ ( .A(_01876_ ), .B(_01877_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01878_ ) );
AOI21_X1 _09453_ ( .A(_01874_ ), .B1(_01875_ ), .B2(_01878_ ), .ZN(_01879_ ) );
OAI221_X1 _09454_ ( .A(_01879_ ), .B1(\IF_ID_pc [16] ), .B2(_01832_ ), .C1(\IF_ID_pc [10] ), .C2(_01851_ ), .ZN(_01880_ ) );
NAND3_X1 _09455_ ( .A1(_01841_ ), .A2(_01843_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01881_ ) );
OAI21_X1 _09456_ ( .A(_01881_ ), .B1(_01875_ ), .B2(_01878_ ), .ZN(_01882_ ) );
NOR2_X1 _09457_ ( .A1(_01820_ ), .A2(\IF_ID_pc [23] ), .ZN(_01883_ ) );
AOI21_X1 _09458_ ( .A(\IF_ID_pc [14] ), .B1(_01871_ ), .B2(_01873_ ), .ZN(_01884_ ) );
NOR4_X1 _09459_ ( .A1(_01880_ ), .A2(_01882_ ), .A3(_01883_ ), .A4(_01884_ ), .ZN(_01885_ ) );
MUX2_X1 _09460_ ( .A(\myifu.myicache.tag[0][8] ), .B(\myifu.myicache.tag[1][8] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01886_ ) );
MUX2_X1 _09461_ ( .A(\myifu.myicache.tag[2][8] ), .B(\myifu.myicache.tag[3][8] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01887_ ) );
MUX2_X1 _09462_ ( .A(_01886_ ), .B(_01887_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01888_ ) );
XNOR2_X1 _09463_ ( .A(_01888_ ), .B(\IF_ID_pc [13] ), .ZN(_01889_ ) );
MUX2_X1 _09464_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01890_ ) );
MUX2_X1 _09465_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01891_ ) );
MUX2_X1 _09466_ ( .A(_01890_ ), .B(_01891_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01892_ ) );
OAI211_X1 _09467_ ( .A(_01889_ ), .B(_01892_ ), .C1(\IF_ID_pc [27] ), .C2(_01816_ ), .ZN(_01893_ ) );
OR2_X1 _09468_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[1][21] ), .ZN(_01894_ ) );
OAI211_X1 _09469_ ( .A(_01894_ ), .B(_01765_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][21] ), .ZN(_01895_ ) );
OR2_X1 _09470_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[3][21] ), .ZN(_01896_ ) );
OAI211_X1 _09471_ ( .A(_01896_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][21] ), .ZN(_01897_ ) );
NAND2_X1 _09472_ ( .A1(_01895_ ), .A2(_01897_ ), .ZN(_01898_ ) );
INV_X1 _09473_ ( .A(\IF_ID_pc [26] ), .ZN(_01899_ ) );
XNOR2_X1 _09474_ ( .A(_01898_ ), .B(_01899_ ), .ZN(_01900_ ) );
OR2_X1 _09475_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01901_ ) );
OAI211_X1 _09476_ ( .A(_01901_ ), .B(_01765_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01902_ ) );
OR2_X1 _09477_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[3][12] ), .ZN(_01903_ ) );
OAI211_X1 _09478_ ( .A(_01903_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][12] ), .ZN(_01904_ ) );
AND3_X1 _09479_ ( .A1(_01902_ ), .A2(_01904_ ), .A3(\IF_ID_pc [17] ), .ZN(_01905_ ) );
AOI21_X1 _09480_ ( .A(\IF_ID_pc [17] ), .B1(_01902_ ), .B2(_01904_ ), .ZN(_01906_ ) );
NOR4_X1 _09481_ ( .A1(_01893_ ), .A2(_01900_ ), .A3(_01905_ ), .A4(_01906_ ), .ZN(_01907_ ) );
OR2_X1 _09482_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[1][1] ), .ZN(_01908_ ) );
OAI211_X1 _09483_ ( .A(_01908_ ), .B(_01765_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][1] ), .ZN(_01909_ ) );
OR2_X1 _09484_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[3][1] ), .ZN(_01910_ ) );
OAI211_X1 _09485_ ( .A(_01910_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][1] ), .ZN(_01911_ ) );
NAND2_X1 _09486_ ( .A1(_01909_ ), .A2(_01911_ ), .ZN(_01912_ ) );
XNOR2_X1 _09487_ ( .A(_01912_ ), .B(\IF_ID_pc [6] ), .ZN(_01913_ ) );
OR2_X1 _09488_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[1][10] ), .ZN(_01914_ ) );
OAI211_X1 _09489_ ( .A(_01914_ ), .B(_01765_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][10] ), .ZN(_01915_ ) );
OR2_X1 _09490_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[3][10] ), .ZN(_01916_ ) );
OAI211_X1 _09491_ ( .A(_01916_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][10] ), .ZN(_01917_ ) );
NAND2_X1 _09492_ ( .A1(_01915_ ), .A2(_01917_ ), .ZN(_01918_ ) );
XNOR2_X1 _09493_ ( .A(_01918_ ), .B(\IF_ID_pc [15] ), .ZN(_01919_ ) );
OR2_X2 _09494_ ( .A1(_01853_ ), .A2(\myifu.myicache.tag[1][17] ), .ZN(_01920_ ) );
OAI211_X1 _09495_ ( .A(_01920_ ), .B(_01764_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][17] ), .ZN(_01921_ ) );
OR2_X1 _09496_ ( .A1(_01760_ ), .A2(\myifu.myicache.tag[3][17] ), .ZN(_01922_ ) );
OAI211_X1 _09497_ ( .A(_01922_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][17] ), .ZN(_01923_ ) );
NAND2_X1 _09498_ ( .A1(_01921_ ), .A2(_01923_ ), .ZN(_01924_ ) );
XNOR2_X1 _09499_ ( .A(_01924_ ), .B(\IF_ID_pc [22] ), .ZN(_01925_ ) );
OR2_X1 _09500_ ( .A1(_01760_ ), .A2(\myifu.myicache.tag[1][4] ), .ZN(_01926_ ) );
OAI211_X1 _09501_ ( .A(_01926_ ), .B(_01764_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][4] ), .ZN(_01927_ ) );
OR2_X1 _09502_ ( .A1(_01760_ ), .A2(\myifu.myicache.tag[3][4] ), .ZN(_01928_ ) );
OAI211_X1 _09503_ ( .A(_01928_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][4] ), .ZN(_01929_ ) );
NAND2_X1 _09504_ ( .A1(_01927_ ), .A2(_01929_ ), .ZN(_01930_ ) );
XNOR2_X1 _09505_ ( .A(_01930_ ), .B(\IF_ID_pc [9] ), .ZN(_01931_ ) );
AND4_X1 _09506_ ( .A1(_01913_ ), .A2(_01919_ ), .A3(_01925_ ), .A4(_01931_ ), .ZN(_01932_ ) );
AND3_X1 _09507_ ( .A1(_01885_ ), .A2(_01907_ ), .A3(_01932_ ), .ZN(_01933_ ) );
AND2_X4 _09508_ ( .A1(_01869_ ), .A2(_01933_ ), .ZN(_01934_ ) );
INV_X1 _09509_ ( .A(\myifu.state [0] ), .ZN(_01935_ ) );
NOR2_X4 _09510_ ( .A1(_01934_ ), .A2(_01935_ ), .ZN(_01936_ ) );
INV_X2 _09511_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01937_ ) );
NOR2_X4 _09512_ ( .A1(_01936_ ), .A2(_01937_ ), .ZN(_01938_ ) );
NOR2_X1 _09513_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01939_ ) );
NOR2_X4 _09514_ ( .A1(_01938_ ), .A2(_01939_ ), .ZN(_01940_ ) );
INV_X32 _09515_ ( .A(\EX_LS_flag [2] ), .ZN(_01941_ ) );
NAND4_X1 _09516_ ( .A1(_01941_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(EXU_valid_LSU ), .ZN(_01942_ ) );
NOR2_X1 _09517_ ( .A1(_01942_ ), .A2(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01943_ ) );
INV_X1 _09518_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01944_ ) );
NOR2_X1 _09519_ ( .A1(_01943_ ), .A2(_01944_ ), .ZN(_01945_ ) );
NOR2_X4 _09520_ ( .A1(_01940_ ), .A2(_01945_ ), .ZN(_01946_ ) );
BUF_X8 _09521_ ( .A(_01946_ ), .Z(_01947_ ) );
CLKBUF_X2 _09522_ ( .A(_01942_ ), .Z(_01948_ ) );
OR3_X1 _09523_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01949_ ) );
BUF_X4 _09524_ ( .A(_01943_ ), .Z(_01950_ ) );
OAI211_X1 _09525_ ( .A(_01947_ ), .B(_01949_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01950_ ), .ZN(_01951_ ) );
INV_X1 _09526_ ( .A(\IF_ID_pc [23] ), .ZN(_01952_ ) );
BUF_X16 _09527_ ( .A(_01940_ ), .Z(_01953_ ) );
INV_X16 _09528_ ( .A(_01953_ ), .ZN(_01954_ ) );
OAI21_X2 _09529_ ( .A(_01951_ ), .B1(_01952_ ), .B2(_01954_ ), .ZN(\io_master_araddr [23] ) );
OR3_X1 _09530_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01955_ ) );
OAI211_X2 _09531_ ( .A(_01947_ ), .B(_01955_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01950_ ), .ZN(_01956_ ) );
INV_X1 _09532_ ( .A(\IF_ID_pc [17] ), .ZN(_01957_ ) );
OAI21_X2 _09533_ ( .A(_01956_ ), .B1(_01957_ ), .B2(_01954_ ), .ZN(\io_master_araddr [17] ) );
OR2_X1 _09534_ ( .A1(\io_master_araddr [23] ), .A2(\io_master_araddr [17] ), .ZN(_01958_ ) );
INV_X1 _09535_ ( .A(_01945_ ), .ZN(_01959_ ) );
MUX2_X1 _09536_ ( .A(\mylsu.araddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_01943_ ), .Z(_01960_ ) );
AND3_X4 _09537_ ( .A1(_01954_ ), .A2(_01959_ ), .A3(_01960_ ), .ZN(_01961_ ) );
AOI21_X2 _09538_ ( .A(_01961_ ), .B1(\IF_ID_pc [25] ), .B2(_01953_ ), .ZN(_01962_ ) );
INV_X4 _09539_ ( .A(_01962_ ), .ZN(\io_master_araddr [25] ) );
CLKBUF_X2 _09540_ ( .A(_01948_ ), .Z(_01963_ ) );
OR3_X1 _09541_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01964_ ) );
BUF_X4 _09542_ ( .A(_01943_ ), .Z(_01965_ ) );
OAI211_X1 _09543_ ( .A(_01947_ ), .B(_01964_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01965_ ), .ZN(_01966_ ) );
BUF_X4 _09544_ ( .A(_01936_ ), .Z(_01967_ ) );
BUF_X4 _09545_ ( .A(_01937_ ), .Z(_01968_ ) );
OAI221_X1 _09546_ ( .A(\IF_ID_pc [30] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_01969_ ) );
AND2_X1 _09547_ ( .A1(_01966_ ), .A2(_01969_ ), .ZN(_01970_ ) );
OR3_X1 _09548_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01971_ ) );
OAI211_X1 _09549_ ( .A(_01947_ ), .B(_01971_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01950_ ), .ZN(_01972_ ) );
OAI221_X1 _09550_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01937_ ), .ZN(_01973_ ) );
AND2_X2 _09551_ ( .A1(_01972_ ), .A2(_01973_ ), .ZN(_01974_ ) );
BUF_X4 _09552_ ( .A(_01946_ ), .Z(_01975_ ) );
OR3_X1 _09553_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01976_ ) );
OAI211_X1 _09554_ ( .A(_01975_ ), .B(_01976_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01965_ ), .ZN(_01977_ ) );
OAI221_X1 _09555_ ( .A(\IF_ID_pc [24] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_01978_ ) );
AND2_X2 _09556_ ( .A1(_01977_ ), .A2(_01978_ ), .ZN(_01979_ ) );
NAND4_X1 _09557_ ( .A1(\io_master_araddr [25] ), .A2(_01970_ ), .A3(_01974_ ), .A4(_01979_ ), .ZN(_01980_ ) );
OR3_X1 _09558_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01981_ ) );
OAI211_X2 _09559_ ( .A(_01947_ ), .B(_01981_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01950_ ), .ZN(_01982_ ) );
OAI21_X4 _09560_ ( .A(_01982_ ), .B1(_01797_ ), .B2(_01954_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09561_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01983_ ) );
OAI211_X2 _09562_ ( .A(_01947_ ), .B(_01983_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01950_ ), .ZN(_01984_ ) );
INV_X1 _09563_ ( .A(\IF_ID_pc [18] ), .ZN(_01985_ ) );
OAI21_X4 _09564_ ( .A(_01984_ ), .B1(_01985_ ), .B2(_01954_ ), .ZN(\io_master_araddr [18] ) );
OR4_X2 _09565_ ( .A1(_01958_ ), .A2(_01980_ ), .A3(\io_master_araddr [20] ), .A4(\io_master_araddr [18] ), .ZN(_01986_ ) );
INV_X1 _09566_ ( .A(\myclint.rvalid ), .ZN(_01987_ ) );
OR3_X1 _09567_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01988_ ) );
OAI211_X1 _09568_ ( .A(_01947_ ), .B(_01988_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01950_ ), .ZN(_01989_ ) );
OAI221_X1 _09569_ ( .A(\IF_ID_pc [28] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01936_ ), .C2(_01937_ ), .ZN(_01990_ ) );
AND2_X2 _09570_ ( .A1(_01989_ ), .A2(_01990_ ), .ZN(_01991_ ) );
OR3_X1 _09571_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01992_ ) );
OAI211_X1 _09572_ ( .A(_01947_ ), .B(_01992_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01965_ ), .ZN(_01993_ ) );
OAI221_X1 _09573_ ( .A(\IF_ID_pc [26] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_01994_ ) );
AND2_X2 _09574_ ( .A1(_01993_ ), .A2(_01994_ ), .ZN(_01995_ ) );
OR3_X1 _09575_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01996_ ) );
OAI211_X1 _09576_ ( .A(_01946_ ), .B(_01996_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01950_ ), .ZN(_01997_ ) );
OAI221_X1 _09577_ ( .A(\IF_ID_pc [21] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01936_ ), .C2(_01937_ ), .ZN(_01998_ ) );
AND2_X1 _09578_ ( .A1(_01997_ ), .A2(_01998_ ), .ZN(_01999_ ) );
OR3_X1 _09579_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02000_ ) );
OAI211_X1 _09580_ ( .A(_01946_ ), .B(_02000_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01950_ ), .ZN(_02001_ ) );
OAI221_X1 _09581_ ( .A(\IF_ID_pc [19] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01936_ ), .C2(_01937_ ), .ZN(_02002_ ) );
AND2_X1 _09582_ ( .A1(_02001_ ), .A2(_02002_ ), .ZN(_02003_ ) );
AND4_X1 _09583_ ( .A1(_01991_ ), .A2(_01995_ ), .A3(_01999_ ), .A4(_02003_ ), .ZN(_02004_ ) );
OR3_X1 _09584_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02005_ ) );
OAI211_X1 _09585_ ( .A(_01947_ ), .B(_02005_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01950_ ), .ZN(_02006_ ) );
OAI221_X1 _09586_ ( .A(\IF_ID_pc [29] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01936_ ), .C2(_01937_ ), .ZN(_02007_ ) );
AND2_X2 _09587_ ( .A1(_02006_ ), .A2(_02007_ ), .ZN(_02008_ ) );
OR3_X1 _09588_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02009_ ) );
OAI211_X1 _09589_ ( .A(_01947_ ), .B(_02009_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01965_ ), .ZN(_02010_ ) );
OAI221_X1 _09590_ ( .A(\IF_ID_pc [27] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_02011_ ) );
AND2_X2 _09591_ ( .A1(_02010_ ), .A2(_02011_ ), .ZN(_02012_ ) );
OR3_X1 _09592_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02013_ ) );
OAI211_X1 _09593_ ( .A(_01946_ ), .B(_02013_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01950_ ), .ZN(_02014_ ) );
OAI221_X1 _09594_ ( .A(\IF_ID_pc [22] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01936_ ), .C2(_01937_ ), .ZN(_02015_ ) );
AND2_X1 _09595_ ( .A1(_02014_ ), .A2(_02015_ ), .ZN(_02016_ ) );
OR3_X1 _09596_ ( .A1(_01948_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02017_ ) );
OAI211_X1 _09597_ ( .A(_01946_ ), .B(_02017_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01943_ ), .ZN(_02018_ ) );
OAI221_X1 _09598_ ( .A(\IF_ID_pc [16] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01936_ ), .C2(_01937_ ), .ZN(_02019_ ) );
AND2_X1 _09599_ ( .A1(_02018_ ), .A2(_02019_ ), .ZN(_02020_ ) );
AND4_X1 _09600_ ( .A1(_02008_ ), .A2(_02012_ ), .A3(_02016_ ), .A4(_02020_ ), .ZN(_02021_ ) );
NAND2_X1 _09601_ ( .A1(_02004_ ), .A2(_02021_ ), .ZN(_02022_ ) );
NOR3_X1 _09602_ ( .A1(_01986_ ), .A2(_01987_ ), .A3(_02022_ ), .ZN(_02023_ ) );
CLKBUF_X2 _09603_ ( .A(_01953_ ), .Z(_02024_ ) );
CLKBUF_X2 _09604_ ( .A(_02024_ ), .Z(_02025_ ) );
CLKBUF_X2 _09605_ ( .A(_02025_ ), .Z(_02026_ ) );
CLKBUF_X2 _09606_ ( .A(_02026_ ), .Z(_02027_ ) );
INV_X1 _09607_ ( .A(\EX_LS_typ [0] ), .ZN(_02028_ ) );
NOR2_X1 _09608_ ( .A1(fanout_net_3 ), .A2(\EX_LS_dest_csreg_mem [1] ), .ZN(_02029_ ) );
INV_X1 _09609_ ( .A(\EX_LS_typ [2] ), .ZN(_02030_ ) );
NOR4_X1 _09610_ ( .A1(_02029_ ), .A2(_02030_ ), .A3(\EX_LS_typ [1] ), .A4(\EX_LS_typ [3] ), .ZN(_02031_ ) );
AND2_X1 _09611_ ( .A1(fanout_net_3 ), .A2(\EX_LS_typ [1] ), .ZN(_02032_ ) );
NOR2_X1 _09612_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02033_ ) );
AND2_X1 _09613_ ( .A1(_02032_ ), .A2(_02033_ ), .ZN(_02034_ ) );
OAI21_X1 _09614_ ( .A(_02028_ ), .B1(_02031_ ), .B2(_02034_ ), .ZN(_02035_ ) );
NAND3_X1 _09615_ ( .A1(_02032_ ), .A2(_02033_ ), .A3(\EX_LS_typ [0] ), .ZN(_02036_ ) );
NAND2_X1 _09616_ ( .A1(_02035_ ), .A2(_02036_ ), .ZN(_02037_ ) );
AND2_X4 _09617_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02038_ ) );
AND2_X2 _09618_ ( .A1(_02038_ ), .A2(_01941_ ), .ZN(_02039_ ) );
INV_X1 _09619_ ( .A(_02039_ ), .ZN(_02040_ ) );
NOR2_X1 _09620_ ( .A1(_02040_ ), .A2(\EX_LS_typ [4] ), .ZN(_02041_ ) );
AND2_X1 _09621_ ( .A1(_02037_ ), .A2(_02041_ ), .ZN(_02042_ ) );
OR2_X1 _09622_ ( .A1(\EX_LS_dest_csreg_mem [27] ), .A2(\EX_LS_dest_csreg_mem [25] ), .ZN(_02043_ ) );
NOR3_X1 _09623_ ( .A1(_02043_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(\EX_LS_dest_csreg_mem [24] ), .ZN(_02044_ ) );
NOR4_X1 _09624_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\EX_LS_dest_csreg_mem [29] ), .A4(\EX_LS_dest_csreg_mem [28] ), .ZN(_02045_ ) );
AND2_X1 _09625_ ( .A1(_02044_ ), .A2(_02045_ ), .ZN(_02046_ ) );
AND2_X1 _09626_ ( .A1(_02046_ ), .A2(_02039_ ), .ZN(_02047_ ) );
NOR2_X1 _09627_ ( .A1(_02042_ ), .A2(_02047_ ), .ZN(_02048_ ) );
INV_X32 _09628_ ( .A(\EX_LS_flag [1] ), .ZN(_02049_ ) );
NOR2_X4 _09629_ ( .A1(_02049_ ), .A2(\EX_LS_flag [0] ), .ZN(_02050_ ) );
AND2_X1 _09630_ ( .A1(_02050_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02051_ ) );
AND2_X1 _09631_ ( .A1(_02046_ ), .A2(_02051_ ), .ZN(_02052_ ) );
INV_X1 _09632_ ( .A(_02029_ ), .ZN(_02053_ ) );
AND3_X1 _09633_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02054_ ) );
AOI22_X1 _09634_ ( .A1(_02053_ ), .A2(_02054_ ), .B1(_02032_ ), .B2(_02033_ ), .ZN(_02055_ ) );
NOR3_X1 _09635_ ( .A1(_02028_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_typ [4] ), .ZN(_02056_ ) );
NAND2_X1 _09636_ ( .A1(_02056_ ), .A2(_02050_ ), .ZN(_02057_ ) );
NOR2_X1 _09637_ ( .A1(_02055_ ), .A2(_02057_ ), .ZN(_02058_ ) );
NOR2_X1 _09638_ ( .A1(_02052_ ), .A2(_02058_ ), .ZN(_02059_ ) );
AND2_X1 _09639_ ( .A1(_02048_ ), .A2(_02059_ ), .ZN(_02060_ ) );
AOI211_X1 _09640_ ( .A(_01944_ ), .B(_02027_ ), .C1(_01965_ ), .C2(_02060_ ), .ZN(_02061_ ) );
NOR2_X1 _09641_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02062_ ) );
INV_X2 _09642_ ( .A(_02062_ ), .ZN(_02063_ ) );
NOR3_X1 _09643_ ( .A1(_01934_ ), .A2(_01935_ ), .A3(_02063_ ), .ZN(_02064_ ) );
NOR4_X1 _09644_ ( .A1(_01938_ ), .A2(_02064_ ), .A3(_01968_ ), .A4(_01939_ ), .ZN(_02065_ ) );
NOR2_X1 _09645_ ( .A1(_02061_ ), .A2(_02065_ ), .ZN(_02066_ ) );
NAND4_X1 _09646_ ( .A1(\io_master_araddr [25] ), .A2(_01970_ ), .A3(_02008_ ), .A4(_02012_ ), .ZN(_02067_ ) );
NOR4_X2 _09647_ ( .A1(_02067_ ), .A2(_01958_ ), .A3(\io_master_araddr [20] ), .A4(\io_master_araddr [18] ), .ZN(_02068_ ) );
NAND4_X1 _09648_ ( .A1(_01974_ ), .A2(_01979_ ), .A3(_01991_ ), .A4(_01995_ ), .ZN(_02069_ ) );
NAND4_X1 _09649_ ( .A1(_01999_ ), .A2(_02003_ ), .A3(_02016_ ), .A4(_02020_ ), .ZN(_02070_ ) );
NOR2_X1 _09650_ ( .A1(_02069_ ), .A2(_02070_ ), .ZN(_02071_ ) );
AND2_X2 _09651_ ( .A1(_02068_ ), .A2(_02071_ ), .ZN(_02072_ ) );
INV_X1 _09652_ ( .A(_02072_ ), .ZN(_02073_ ) );
AOI21_X1 _09653_ ( .A(_02027_ ), .B1(_01965_ ), .B2(_02060_ ), .ZN(_02074_ ) );
AOI211_X1 _09654_ ( .A(_01939_ ), .B(_01938_ ), .C1(\myifu.state [0] ), .C2(_02062_ ), .ZN(_02075_ ) );
OR3_X1 _09655_ ( .A1(_02073_ ), .A2(_02074_ ), .A3(_02075_ ), .ZN(_02076_ ) );
AOI221_X4 _09656_ ( .A(fanout_net_2 ), .B1(_02023_ ), .B2(_02066_ ), .C1(_02076_ ), .C2(_01987_ ), .ZN(_00064_ ) );
INV_X1 _09657_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02077_ ) );
CLKBUF_X2 _09658_ ( .A(_02077_ ), .Z(_02078_ ) );
AND2_X1 _09659_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00065_ ) );
AND2_X1 _09660_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00066_ ) );
AND2_X1 _09661_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00067_ ) );
INV_X1 _09662_ ( .A(\LS_WB_wdata_csreg [20] ), .ZN(_02079_ ) );
NOR2_X1 _09663_ ( .A1(_02079_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00068_ ) );
AND2_X1 _09664_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [19] ), .ZN(_00069_ ) );
AND2_X1 _09665_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [18] ), .ZN(_00070_ ) );
AND2_X1 _09666_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [17] ), .ZN(_00071_ ) );
AND2_X1 _09667_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00072_ ) );
AND2_X1 _09668_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00073_ ) );
AND2_X1 _09669_ ( .A1(_02078_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00074_ ) );
CLKBUF_X2 _09670_ ( .A(_02077_ ), .Z(_02080_ ) );
AND2_X1 _09671_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00075_ ) );
AND2_X1 _09672_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00076_ ) );
AND2_X1 _09673_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00077_ ) );
AND2_X1 _09674_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00078_ ) );
AND2_X1 _09675_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00079_ ) );
AND2_X1 _09676_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00080_ ) );
AND2_X1 _09677_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00081_ ) );
AND2_X1 _09678_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00082_ ) );
INV_X1 _09679_ ( .A(\LS_WB_wdata_csreg [6] ), .ZN(_02081_ ) );
NOR2_X1 _09680_ ( .A1(_02081_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00083_ ) );
AND2_X1 _09681_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00084_ ) );
AND2_X1 _09682_ ( .A1(_02080_ ), .A2(\LS_WB_wdata_csreg [4] ), .ZN(_00085_ ) );
AND2_X1 _09683_ ( .A1(_02077_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00086_ ) );
AND2_X1 _09684_ ( .A1(_02077_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00087_ ) );
AND2_X1 _09685_ ( .A1(_02077_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00088_ ) );
AND2_X1 _09686_ ( .A1(_02077_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00089_ ) );
AND2_X1 _09687_ ( .A1(_02077_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00090_ ) );
AND2_X1 _09688_ ( .A1(_02077_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00091_ ) );
AND2_X1 _09689_ ( .A1(_02077_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00092_ ) );
AOI21_X1 _09690_ ( .A(excp_written ), .B1(\LS_WB_wen_csreg [6] ), .B2(\LS_WB_wen_csreg [7] ), .ZN(_02082_ ) );
NOR2_X1 _09691_ ( .A1(_02082_ ), .A2(fanout_net_2 ), .ZN(_00093_ ) );
INV_X1 _09692_ ( .A(_02048_ ), .ZN(_02083_ ) );
INV_X1 _09693_ ( .A(_02059_ ), .ZN(_02084_ ) );
OR2_X1 _09694_ ( .A1(\myexu.pc_jump [26] ), .A2(\myexu.pc_jump [25] ), .ZN(_02085_ ) );
OR3_X1 _09695_ ( .A1(_02085_ ), .A2(\myexu.pc_jump [27] ), .A3(\myexu.pc_jump [24] ), .ZN(_02086_ ) );
OR4_X1 _09696_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02087_ ) );
NOR2_X1 _09697_ ( .A1(_02086_ ), .A2(_02087_ ), .ZN(_02088_ ) );
NOR2_X1 _09698_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02089_ ) );
INV_X1 _09699_ ( .A(_02089_ ), .ZN(_02090_ ) );
NOR3_X1 _09700_ ( .A1(_02088_ ), .A2(exception_quest_IDU ), .A3(_02090_ ), .ZN(_02091_ ) );
NOR2_X1 _09701_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02092_ ) );
AND2_X1 _09702_ ( .A1(_02092_ ), .A2(_01534_ ), .ZN(_02093_ ) );
INV_X1 _09703_ ( .A(_02093_ ), .ZN(_02094_ ) );
NOR4_X1 _09704_ ( .A1(_02083_ ), .A2(_02084_ ), .A3(_02091_ ), .A4(_02094_ ), .ZN(_00094_ ) );
AOI21_X1 _09705_ ( .A(_02094_ ), .B1(_02060_ ), .B2(exception_quest_IDU ), .ZN(_00095_ ) );
INV_X1 _09706_ ( .A(fanout_net_26 ), .ZN(_02095_ ) );
BUF_X4 _09707_ ( .A(_02095_ ), .Z(_02096_ ) );
BUF_X4 _09708_ ( .A(_02096_ ), .Z(_02097_ ) );
BUF_X4 _09709_ ( .A(_02097_ ), .Z(_02098_ ) );
INV_X2 _09710_ ( .A(fanout_net_25 ), .ZN(_02099_ ) );
BUF_X4 _09711_ ( .A(_02099_ ), .Z(_02100_ ) );
BUF_X4 _09712_ ( .A(_02100_ ), .Z(_02101_ ) );
BUF_X4 _09713_ ( .A(_02101_ ), .Z(_02102_ ) );
MUX2_X1 _09714_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02103_ ) );
AND2_X1 _09715_ ( .A1(_02103_ ), .A2(fanout_net_23 ), .ZN(_02104_ ) );
INV_X2 _09716_ ( .A(fanout_net_23 ), .ZN(_02105_ ) );
BUF_X4 _09717_ ( .A(_02105_ ), .Z(_02106_ ) );
BUF_X4 _09718_ ( .A(_02106_ ), .Z(_02107_ ) );
BUF_X4 _09719_ ( .A(_02107_ ), .Z(_02108_ ) );
BUF_X4 _09720_ ( .A(_02108_ ), .Z(_02109_ ) );
BUF_X4 _09721_ ( .A(_02109_ ), .Z(_02110_ ) );
MUX2_X1 _09722_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02111_ ) );
AOI211_X1 _09723_ ( .A(_02102_ ), .B(_02104_ ), .C1(_02110_ ), .C2(_02111_ ), .ZN(_02112_ ) );
BUF_X4 _09724_ ( .A(_02102_ ), .Z(_02113_ ) );
AND2_X1 _09725_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02114_ ) );
INV_X1 _09726_ ( .A(fanout_net_14 ), .ZN(_02115_ ) );
BUF_X2 _09727_ ( .A(_02115_ ), .Z(_02116_ ) );
BUF_X2 _09728_ ( .A(_02116_ ), .Z(_02117_ ) );
BUF_X2 _09729_ ( .A(_02117_ ), .Z(_02118_ ) );
BUF_X2 _09730_ ( .A(_02118_ ), .Z(_02119_ ) );
CLKBUF_X2 _09731_ ( .A(_02119_ ), .Z(_02120_ ) );
BUF_X4 _09732_ ( .A(_02120_ ), .Z(_02121_ ) );
AOI21_X1 _09733_ ( .A(_02114_ ), .B1(_02121_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02122_ ) );
AND2_X1 _09734_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02123_ ) );
AOI21_X1 _09735_ ( .A(_02123_ ), .B1(_02121_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02124_ ) );
BUF_X4 _09736_ ( .A(_02108_ ), .Z(_02125_ ) );
MUX2_X1 _09737_ ( .A(_02122_ ), .B(_02124_ ), .S(_02125_ ), .Z(_02126_ ) );
AOI211_X1 _09738_ ( .A(_02098_ ), .B(_02112_ ), .C1(_02113_ ), .C2(_02126_ ), .ZN(_02127_ ) );
AND2_X4 _09739_ ( .A1(_02050_ ), .A2(\EX_LS_flag [2] ), .ZN(_02128_ ) );
NOR2_X2 _09740_ ( .A1(_02128_ ), .A2(_02039_ ), .ZN(_02129_ ) );
OAI211_X1 _09741_ ( .A(_02049_ ), .B(\EX_LS_flag [0] ), .C1(\EX_LS_flag [2] ), .C2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02130_ ) );
AND2_X4 _09742_ ( .A1(_02129_ ), .A2(_02130_ ), .ZN(_02131_ ) );
XNOR2_X1 _09743_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02132_ ) );
INV_X4 _09744_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02133_ ) );
NAND2_X1 _09745_ ( .A1(_02133_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02134_ ) );
OR3_X1 _09746_ ( .A1(\EX_LS_dest_reg [2] ), .A2(\EX_LS_dest_reg [1] ), .A3(\EX_LS_dest_reg [0] ), .ZN(_02135_ ) );
OR2_X1 _09747_ ( .A1(\EX_LS_dest_reg [4] ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02136_ ) );
OAI211_X1 _09748_ ( .A(_02132_ ), .B(_02134_ ), .C1(_02135_ ), .C2(_02136_ ), .ZN(_02137_ ) );
OR2_X2 _09749_ ( .A1(_02131_ ), .A2(_02137_ ), .ZN(_02138_ ) );
BUF_X4 _09750_ ( .A(_02138_ ), .Z(_02139_ ) );
XNOR2_X1 _09751_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .ZN(_02140_ ) );
INV_X1 _09752_ ( .A(\ID_EX_rs1 [3] ), .ZN(_02141_ ) );
NAND2_X1 _09753_ ( .A1(_02141_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02142_ ) );
NAND3_X1 _09754_ ( .A1(_02140_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y ), .A3(_02142_ ), .ZN(_02143_ ) );
XOR2_X2 _09755_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .Z(_02144_ ) );
OAI22_X1 _09756_ ( .A1(_02141_ ), .A2(\EX_LS_dest_reg [3] ), .B1(_02133_ ), .B2(\ID_EX_rs1 [1] ), .ZN(_02145_ ) );
OR3_X4 _09757_ ( .A1(_02143_ ), .A2(_02144_ ), .A3(_02145_ ), .ZN(_02146_ ) );
CLKBUF_X2 _09758_ ( .A(_02146_ ), .Z(_02147_ ) );
NOR2_X1 _09759_ ( .A1(_02139_ ), .A2(_02147_ ), .ZN(_02148_ ) );
BUF_X4 _09760_ ( .A(_02102_ ), .Z(_02149_ ) );
MUX2_X1 _09761_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02150_ ) );
AND2_X1 _09762_ ( .A1(_02150_ ), .A2(fanout_net_23 ), .ZN(_02151_ ) );
MUX2_X1 _09763_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02152_ ) );
AOI211_X1 _09764_ ( .A(_02149_ ), .B(_02151_ ), .C1(_02110_ ), .C2(_02152_ ), .ZN(_02153_ ) );
INV_X1 _09765_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02154_ ) );
AOI21_X1 _09766_ ( .A(fanout_net_23 ), .B1(_02154_ ), .B2(fanout_net_14 ), .ZN(_02155_ ) );
OR2_X1 _09767_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02156_ ) );
MUX2_X1 _09768_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02157_ ) );
AOI221_X4 _09769_ ( .A(fanout_net_25 ), .B1(_02155_ ), .B2(_02156_ ), .C1(_02157_ ), .C2(fanout_net_23 ), .ZN(_02158_ ) );
NOR3_X1 _09770_ ( .A1(_02153_ ), .A2(fanout_net_26 ), .A3(_02158_ ), .ZN(_02159_ ) );
OR3_X1 _09771_ ( .A1(_02127_ ), .A2(_02148_ ), .A3(_02159_ ), .ZN(_02160_ ) );
BUF_X4 _09772_ ( .A(_02131_ ), .Z(_02161_ ) );
CLKBUF_X2 _09773_ ( .A(_02161_ ), .Z(_02162_ ) );
BUF_X2 _09774_ ( .A(_02162_ ), .Z(_02163_ ) );
BUF_X2 _09775_ ( .A(_02163_ ), .Z(_02164_ ) );
CLKBUF_X2 _09776_ ( .A(_02146_ ), .Z(_02165_ ) );
BUF_X2 _09777_ ( .A(_02165_ ), .Z(_02166_ ) );
BUF_X2 _09778_ ( .A(_02166_ ), .Z(_02167_ ) );
BUF_X2 _09779_ ( .A(_02167_ ), .Z(_02168_ ) );
CLKBUF_X2 _09780_ ( .A(_02137_ ), .Z(_02169_ ) );
CLKBUF_X2 _09781_ ( .A(_02169_ ), .Z(_02170_ ) );
OR4_X1 _09782_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A2(_02164_ ), .A3(_02168_ ), .A4(_02170_ ), .ZN(_02171_ ) );
AND2_X2 _09783_ ( .A1(_02160_ ), .A2(_02171_ ), .ZN(_02172_ ) );
INV_X1 _09784_ ( .A(\ID_EX_imm [30] ), .ZN(_02173_ ) );
XNOR2_X1 _09785_ ( .A(_02172_ ), .B(_02173_ ), .ZN(_02174_ ) );
OR2_X1 _09786_ ( .A1(_02120_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02175_ ) );
OAI211_X1 _09787_ ( .A(_02175_ ), .B(fanout_net_23 ), .C1(fanout_net_14 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02176_ ) );
INV_X1 _09788_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02177_ ) );
NAND2_X1 _09789_ ( .A1(_02177_ ), .A2(fanout_net_14 ), .ZN(_02178_ ) );
OAI211_X1 _09790_ ( .A(_02178_ ), .B(_02109_ ), .C1(fanout_net_14 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02179_ ) );
NAND3_X1 _09791_ ( .A1(_02176_ ), .A2(_02149_ ), .A3(_02179_ ), .ZN(_02180_ ) );
MUX2_X1 _09792_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02181_ ) );
MUX2_X1 _09793_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02182_ ) );
MUX2_X1 _09794_ ( .A(_02181_ ), .B(_02182_ ), .S(_02109_ ), .Z(_02183_ ) );
OAI211_X1 _09795_ ( .A(fanout_net_26 ), .B(_02180_ ), .C1(_02183_ ), .C2(_02113_ ), .ZN(_02184_ ) );
OR2_X1 _09796_ ( .A1(fanout_net_14 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02185_ ) );
OAI211_X1 _09797_ ( .A(_02185_ ), .B(_02109_ ), .C1(_02121_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02186_ ) );
INV_X1 _09798_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02187_ ) );
NAND2_X1 _09799_ ( .A1(_02187_ ), .A2(fanout_net_14 ), .ZN(_02188_ ) );
OAI211_X1 _09800_ ( .A(_02188_ ), .B(fanout_net_23 ), .C1(fanout_net_14 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02189_ ) );
NAND3_X1 _09801_ ( .A1(_02186_ ), .A2(_02189_ ), .A3(_02149_ ), .ZN(_02190_ ) );
MUX2_X1 _09802_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02191_ ) );
MUX2_X1 _09803_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02192_ ) );
MUX2_X1 _09804_ ( .A(_02191_ ), .B(_02192_ ), .S(_02109_ ), .Z(_02193_ ) );
OAI211_X1 _09805_ ( .A(_02098_ ), .B(_02190_ ), .C1(_02193_ ), .C2(_02149_ ), .ZN(_02194_ ) );
BUF_X4 _09806_ ( .A(_02139_ ), .Z(_02195_ ) );
OAI211_X1 _09807_ ( .A(_02184_ ), .B(_02194_ ), .C1(_02195_ ), .C2(_02168_ ), .ZN(_02196_ ) );
CLKBUF_X2 _09808_ ( .A(_02163_ ), .Z(_02197_ ) );
OR4_X1 _09809_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02197_ ), .A3(_02167_ ), .A4(_02170_ ), .ZN(_02198_ ) );
NAND2_X1 _09810_ ( .A1(_02196_ ), .A2(_02198_ ), .ZN(_02199_ ) );
INV_X1 _09811_ ( .A(\ID_EX_imm [29] ), .ZN(_02200_ ) );
XNOR2_X1 _09812_ ( .A(_02199_ ), .B(_02200_ ), .ZN(_02201_ ) );
NAND2_X1 _09813_ ( .A1(_02148_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_02202_ ) );
OR2_X1 _09814_ ( .A1(_02120_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02203_ ) );
OAI211_X1 _09815_ ( .A(_02203_ ), .B(fanout_net_23 ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02204_ ) );
INV_X1 _09816_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02205_ ) );
NAND2_X1 _09817_ ( .A1(_02205_ ), .A2(fanout_net_14 ), .ZN(_02206_ ) );
OAI211_X1 _09818_ ( .A(_02206_ ), .B(_02125_ ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02207_ ) );
NAND3_X1 _09819_ ( .A1(_02204_ ), .A2(_02149_ ), .A3(_02207_ ), .ZN(_02208_ ) );
MUX2_X1 _09820_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02209_ ) );
MUX2_X1 _09821_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02210_ ) );
MUX2_X1 _09822_ ( .A(_02209_ ), .B(_02210_ ), .S(_02125_ ), .Z(_02211_ ) );
OAI211_X1 _09823_ ( .A(_02098_ ), .B(_02208_ ), .C1(_02211_ ), .C2(_02113_ ), .ZN(_02212_ ) );
OR2_X1 _09824_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02213_ ) );
OAI211_X1 _09825_ ( .A(_02213_ ), .B(_02125_ ), .C1(_02121_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02214_ ) );
INV_X1 _09826_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02215_ ) );
NAND2_X1 _09827_ ( .A1(_02215_ ), .A2(fanout_net_14 ), .ZN(_02216_ ) );
OAI211_X1 _09828_ ( .A(_02216_ ), .B(fanout_net_23 ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02217_ ) );
NAND3_X1 _09829_ ( .A1(_02214_ ), .A2(_02217_ ), .A3(fanout_net_25 ), .ZN(_02218_ ) );
MUX2_X1 _09830_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02219_ ) );
MUX2_X1 _09831_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_02220_ ) );
MUX2_X1 _09832_ ( .A(_02219_ ), .B(_02220_ ), .S(fanout_net_23 ), .Z(_02221_ ) );
OAI211_X1 _09833_ ( .A(fanout_net_26 ), .B(_02218_ ), .C1(_02221_ ), .C2(fanout_net_25 ), .ZN(_02222_ ) );
NAND2_X1 _09834_ ( .A1(_02212_ ), .A2(_02222_ ), .ZN(_02223_ ) );
OAI21_X1 _09835_ ( .A(_02223_ ), .B1(_02168_ ), .B2(_02195_ ), .ZN(_02224_ ) );
AND2_X1 _09836_ ( .A1(_02202_ ), .A2(_02224_ ), .ZN(_02225_ ) );
BUF_X2 _09837_ ( .A(_02225_ ), .Z(_02226_ ) );
XNOR2_X1 _09838_ ( .A(_02226_ ), .B(\ID_EX_imm [28] ), .ZN(_02227_ ) );
INV_X1 _09839_ ( .A(_02227_ ), .ZN(_02228_ ) );
OR2_X1 _09840_ ( .A1(_02120_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02229_ ) );
OAI211_X1 _09841_ ( .A(_02229_ ), .B(_02110_ ), .C1(fanout_net_15 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02230_ ) );
OR2_X1 _09842_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02231_ ) );
OAI211_X1 _09843_ ( .A(_02231_ ), .B(fanout_net_23 ), .C1(_02121_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02232_ ) );
NAND3_X1 _09844_ ( .A1(_02230_ ), .A2(fanout_net_25 ), .A3(_02232_ ), .ZN(_02233_ ) );
MUX2_X1 _09845_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02234_ ) );
MUX2_X1 _09846_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02235_ ) );
MUX2_X1 _09847_ ( .A(_02234_ ), .B(_02235_ ), .S(_02125_ ), .Z(_02236_ ) );
OAI211_X1 _09848_ ( .A(_02098_ ), .B(_02233_ ), .C1(_02236_ ), .C2(fanout_net_25 ), .ZN(_02237_ ) );
MUX2_X1 _09849_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02238_ ) );
AND2_X1 _09850_ ( .A1(_02238_ ), .A2(fanout_net_23 ), .ZN(_02239_ ) );
MUX2_X1 _09851_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02240_ ) );
AOI211_X1 _09852_ ( .A(fanout_net_25 ), .B(_02239_ ), .C1(_02110_ ), .C2(_02240_ ), .ZN(_02241_ ) );
MUX2_X1 _09853_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02242_ ) );
MUX2_X1 _09854_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02243_ ) );
MUX2_X1 _09855_ ( .A(_02242_ ), .B(_02243_ ), .S(fanout_net_23 ), .Z(_02244_ ) );
OAI21_X1 _09856_ ( .A(fanout_net_26 ), .B1(_02244_ ), .B2(_02113_ ), .ZN(_02245_ ) );
OAI221_X1 _09857_ ( .A(_02237_ ), .B1(_02241_ ), .B2(_02245_ ), .C1(_02195_ ), .C2(_02168_ ), .ZN(_02246_ ) );
OR4_X1 _09858_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A2(_02197_ ), .A3(_02168_ ), .A4(_02170_ ), .ZN(_02247_ ) );
NAND2_X1 _09859_ ( .A1(_02246_ ), .A2(_02247_ ), .ZN(_02248_ ) );
INV_X1 _09860_ ( .A(\ID_EX_imm [27] ), .ZN(_02249_ ) );
XNOR2_X1 _09861_ ( .A(_02248_ ), .B(_02249_ ), .ZN(_02250_ ) );
OR2_X1 _09862_ ( .A1(_02120_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02251_ ) );
OAI211_X1 _09863_ ( .A(_02251_ ), .B(fanout_net_23 ), .C1(fanout_net_15 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02252_ ) );
OR2_X1 _09864_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02253_ ) );
OAI211_X1 _09865_ ( .A(_02253_ ), .B(_02125_ ), .C1(_02121_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02254_ ) );
NAND3_X1 _09866_ ( .A1(_02252_ ), .A2(_02149_ ), .A3(_02254_ ), .ZN(_02255_ ) );
MUX2_X1 _09867_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02256_ ) );
MUX2_X1 _09868_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02257_ ) );
MUX2_X1 _09869_ ( .A(_02256_ ), .B(_02257_ ), .S(_02125_ ), .Z(_02258_ ) );
OAI211_X1 _09870_ ( .A(_02098_ ), .B(_02255_ ), .C1(_02258_ ), .C2(_02113_ ), .ZN(_02259_ ) );
OR2_X1 _09871_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02260_ ) );
OAI211_X1 _09872_ ( .A(_02260_ ), .B(_02125_ ), .C1(_02121_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02261_ ) );
NOR2_X1 _09873_ ( .A1(_02121_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02262_ ) );
OAI21_X1 _09874_ ( .A(fanout_net_23 ), .B1(fanout_net_15 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02263_ ) );
OAI211_X1 _09875_ ( .A(_02261_ ), .B(fanout_net_25 ), .C1(_02262_ ), .C2(_02263_ ), .ZN(_02264_ ) );
MUX2_X1 _09876_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02265_ ) );
MUX2_X1 _09877_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02266_ ) );
MUX2_X1 _09878_ ( .A(_02265_ ), .B(_02266_ ), .S(fanout_net_23 ), .Z(_02267_ ) );
OAI211_X1 _09879_ ( .A(fanout_net_26 ), .B(_02264_ ), .C1(_02267_ ), .C2(fanout_net_25 ), .ZN(_02268_ ) );
OAI211_X1 _09880_ ( .A(_02259_ ), .B(_02268_ ), .C1(_02195_ ), .C2(_02168_ ), .ZN(_02269_ ) );
OR4_X1 _09881_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A2(_02197_ ), .A3(_02167_ ), .A4(_02170_ ), .ZN(_02270_ ) );
NAND2_X1 _09882_ ( .A1(_02269_ ), .A2(_02270_ ), .ZN(_02271_ ) );
INV_X1 _09883_ ( .A(\ID_EX_imm [24] ), .ZN(_02272_ ) );
XNOR2_X1 _09884_ ( .A(_02271_ ), .B(_02272_ ), .ZN(_02273_ ) );
INV_X1 _09885_ ( .A(_02273_ ), .ZN(_02274_ ) );
OR2_X1 _09886_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02275_ ) );
BUF_X4 _09887_ ( .A(_02106_ ), .Z(_02276_ ) );
BUF_X4 _09888_ ( .A(_02276_ ), .Z(_02277_ ) );
CLKBUF_X2 _09889_ ( .A(_02117_ ), .Z(_02278_ ) );
BUF_X2 _09890_ ( .A(_02278_ ), .Z(_02279_ ) );
OAI211_X1 _09891_ ( .A(_02275_ ), .B(_02277_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02280_ ) );
OR2_X1 _09892_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02281_ ) );
OAI211_X1 _09893_ ( .A(_02281_ ), .B(fanout_net_23 ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02282_ ) );
BUF_X4 _09894_ ( .A(_02100_ ), .Z(_02283_ ) );
NAND3_X1 _09895_ ( .A1(_02280_ ), .A2(_02282_ ), .A3(_02283_ ), .ZN(_02284_ ) );
MUX2_X1 _09896_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02285_ ) );
MUX2_X1 _09897_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02286_ ) );
BUF_X4 _09898_ ( .A(_02276_ ), .Z(_02287_ ) );
MUX2_X1 _09899_ ( .A(_02285_ ), .B(_02286_ ), .S(_02287_ ), .Z(_02288_ ) );
BUF_X4 _09900_ ( .A(_02099_ ), .Z(_02289_ ) );
BUF_X4 _09901_ ( .A(_02289_ ), .Z(_02290_ ) );
OAI211_X1 _09902_ ( .A(_02097_ ), .B(_02284_ ), .C1(_02288_ ), .C2(_02290_ ), .ZN(_02291_ ) );
OR2_X1 _09903_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02292_ ) );
OAI211_X1 _09904_ ( .A(_02292_ ), .B(fanout_net_23 ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02293_ ) );
OR2_X1 _09905_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02294_ ) );
OAI211_X1 _09906_ ( .A(_02294_ ), .B(_02277_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02295_ ) );
NAND3_X1 _09907_ ( .A1(_02293_ ), .A2(_02295_ ), .A3(fanout_net_25 ), .ZN(_02296_ ) );
MUX2_X1 _09908_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02297_ ) );
MUX2_X1 _09909_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02298_ ) );
MUX2_X1 _09910_ ( .A(_02297_ ), .B(_02298_ ), .S(fanout_net_23 ), .Z(_02299_ ) );
OAI211_X1 _09911_ ( .A(fanout_net_26 ), .B(_02296_ ), .C1(_02299_ ), .C2(fanout_net_25 ), .ZN(_02300_ ) );
BUF_X4 _09912_ ( .A(_02138_ ), .Z(_02301_ ) );
OAI211_X1 _09913_ ( .A(_02291_ ), .B(_02300_ ), .C1(_02301_ ), .C2(_02167_ ), .ZN(_02302_ ) );
BUF_X8 _09914_ ( .A(_02131_ ), .Z(_02303_ ) );
CLKBUF_X2 _09915_ ( .A(_02303_ ), .Z(_02304_ ) );
CLKBUF_X2 _09916_ ( .A(_02169_ ), .Z(_02305_ ) );
OR4_X1 _09917_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02304_ ), .A3(_02147_ ), .A4(_02305_ ), .ZN(_02306_ ) );
NAND2_X2 _09918_ ( .A1(_02302_ ), .A2(_02306_ ), .ZN(_02307_ ) );
INV_X1 _09919_ ( .A(\ID_EX_imm [23] ), .ZN(_02308_ ) );
XNOR2_X1 _09920_ ( .A(_02307_ ), .B(_02308_ ), .ZN(_02309_ ) );
OR2_X1 _09921_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02310_ ) );
OAI211_X1 _09922_ ( .A(_02310_ ), .B(_02108_ ), .C1(_02119_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02311_ ) );
OR2_X1 _09923_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02312_ ) );
OAI211_X1 _09924_ ( .A(_02312_ ), .B(fanout_net_23 ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02313_ ) );
NAND3_X1 _09925_ ( .A1(_02311_ ), .A2(_02313_ ), .A3(fanout_net_25 ), .ZN(_02314_ ) );
MUX2_X1 _09926_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02315_ ) );
MUX2_X1 _09927_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02316_ ) );
MUX2_X1 _09928_ ( .A(_02315_ ), .B(_02316_ ), .S(_02277_ ), .Z(_02317_ ) );
OAI211_X1 _09929_ ( .A(_02097_ ), .B(_02314_ ), .C1(_02317_ ), .C2(fanout_net_25 ), .ZN(_02318_ ) );
BUF_X2 _09930_ ( .A(_02117_ ), .Z(_02319_ ) );
BUF_X4 _09931_ ( .A(_02319_ ), .Z(_02320_ ) );
NOR2_X1 _09932_ ( .A1(_02320_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02321_ ) );
OAI21_X1 _09933_ ( .A(fanout_net_23 ), .B1(fanout_net_15 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02322_ ) );
NOR2_X1 _09934_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02323_ ) );
OAI21_X1 _09935_ ( .A(_02277_ ), .B1(_02320_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02324_ ) );
OAI221_X1 _09936_ ( .A(_02283_ ), .B1(_02321_ ), .B2(_02322_ ), .C1(_02323_ ), .C2(_02324_ ), .ZN(_02325_ ) );
MUX2_X1 _09937_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02326_ ) );
MUX2_X1 _09938_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02327_ ) );
MUX2_X1 _09939_ ( .A(_02326_ ), .B(_02327_ ), .S(fanout_net_23 ), .Z(_02328_ ) );
OAI211_X1 _09940_ ( .A(fanout_net_26 ), .B(_02325_ ), .C1(_02328_ ), .C2(_02102_ ), .ZN(_02329_ ) );
OAI211_X1 _09941_ ( .A(_02318_ ), .B(_02329_ ), .C1(_02195_ ), .C2(_02167_ ), .ZN(_02330_ ) );
BUF_X2 _09942_ ( .A(_02303_ ), .Z(_02331_ ) );
OR4_X1 _09943_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02331_ ), .A3(_02166_ ), .A4(_02170_ ), .ZN(_02332_ ) );
NAND2_X2 _09944_ ( .A1(_02330_ ), .A2(_02332_ ), .ZN(_02333_ ) );
INV_X1 _09945_ ( .A(\ID_EX_imm [22] ), .ZN(_02334_ ) );
XNOR2_X1 _09946_ ( .A(_02333_ ), .B(_02334_ ), .ZN(_02335_ ) );
AND2_X1 _09947_ ( .A1(_02309_ ), .A2(_02335_ ), .ZN(_02336_ ) );
OR2_X1 _09948_ ( .A1(_02278_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02337_ ) );
OAI211_X1 _09949_ ( .A(_02337_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02338_ ) );
OR2_X1 _09950_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02339_ ) );
OAI211_X1 _09951_ ( .A(_02339_ ), .B(_02277_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02340_ ) );
NAND3_X1 _09952_ ( .A1(_02338_ ), .A2(_02283_ ), .A3(_02340_ ), .ZN(_02341_ ) );
MUX2_X1 _09953_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02342_ ) );
MUX2_X1 _09954_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02343_ ) );
MUX2_X1 _09955_ ( .A(_02342_ ), .B(_02343_ ), .S(_02287_ ), .Z(_02344_ ) );
OAI211_X1 _09956_ ( .A(_02097_ ), .B(_02341_ ), .C1(_02344_ ), .C2(_02290_ ), .ZN(_02345_ ) );
OR2_X1 _09957_ ( .A1(_02278_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02346_ ) );
OAI211_X1 _09958_ ( .A(_02346_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02347_ ) );
OR2_X1 _09959_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02348_ ) );
OAI211_X1 _09960_ ( .A(_02348_ ), .B(_02277_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02349_ ) );
NAND3_X1 _09961_ ( .A1(_02347_ ), .A2(fanout_net_25 ), .A3(_02349_ ), .ZN(_02350_ ) );
MUX2_X1 _09962_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02351_ ) );
MUX2_X1 _09963_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02352_ ) );
MUX2_X1 _09964_ ( .A(_02351_ ), .B(_02352_ ), .S(fanout_net_23 ), .Z(_02353_ ) );
OAI211_X1 _09965_ ( .A(fanout_net_26 ), .B(_02350_ ), .C1(_02353_ ), .C2(fanout_net_25 ), .ZN(_02354_ ) );
BUF_X2 _09966_ ( .A(_02165_ ), .Z(_02355_ ) );
OAI211_X1 _09967_ ( .A(_02345_ ), .B(_02354_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02356_ ) );
INV_X1 _09968_ ( .A(\ID_EX_imm [21] ), .ZN(_02357_ ) );
OR4_X1 _09969_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02304_ ), .A3(_02166_ ), .A4(_02305_ ), .ZN(_02358_ ) );
AND3_X1 _09970_ ( .A1(_02356_ ), .A2(_02357_ ), .A3(_02358_ ), .ZN(_02359_ ) );
AOI21_X1 _09971_ ( .A(_02357_ ), .B1(_02356_ ), .B2(_02358_ ), .ZN(_02360_ ) );
NOR2_X1 _09972_ ( .A1(_02359_ ), .A2(_02360_ ), .ZN(_02361_ ) );
OR2_X1 _09973_ ( .A1(_02279_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02362_ ) );
OAI211_X1 _09974_ ( .A(_02362_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02363_ ) );
OR2_X1 _09975_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02364_ ) );
OAI211_X1 _09976_ ( .A(_02364_ ), .B(_02108_ ), .C1(_02119_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02365_ ) );
NAND3_X1 _09977_ ( .A1(_02363_ ), .A2(_02102_ ), .A3(_02365_ ), .ZN(_02366_ ) );
MUX2_X1 _09978_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02367_ ) );
MUX2_X1 _09979_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02368_ ) );
MUX2_X1 _09980_ ( .A(_02367_ ), .B(_02368_ ), .S(_02108_ ), .Z(_02369_ ) );
OAI211_X1 _09981_ ( .A(_02098_ ), .B(_02366_ ), .C1(_02369_ ), .C2(_02102_ ), .ZN(_02370_ ) );
OR2_X1 _09982_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02371_ ) );
OAI211_X1 _09983_ ( .A(_02371_ ), .B(fanout_net_23 ), .C1(_02119_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02372_ ) );
OR2_X1 _09984_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02373_ ) );
OAI211_X1 _09985_ ( .A(_02373_ ), .B(_02108_ ), .C1(_02119_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02374_ ) );
NAND3_X1 _09986_ ( .A1(_02372_ ), .A2(_02374_ ), .A3(fanout_net_25 ), .ZN(_02375_ ) );
MUX2_X1 _09987_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02376_ ) );
MUX2_X1 _09988_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02377_ ) );
MUX2_X1 _09989_ ( .A(_02376_ ), .B(_02377_ ), .S(fanout_net_23 ), .Z(_02378_ ) );
OAI211_X1 _09990_ ( .A(fanout_net_26 ), .B(_02375_ ), .C1(_02378_ ), .C2(fanout_net_25 ), .ZN(_02379_ ) );
OAI211_X1 _09991_ ( .A(_02370_ ), .B(_02379_ ), .C1(_02195_ ), .C2(_02167_ ), .ZN(_02380_ ) );
OR4_X1 _09992_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02163_ ), .A3(_02355_ ), .A4(_02170_ ), .ZN(_02381_ ) );
NAND2_X2 _09993_ ( .A1(_02380_ ), .A2(_02381_ ), .ZN(_02382_ ) );
INV_X1 _09994_ ( .A(\ID_EX_imm [20] ), .ZN(_02383_ ) );
XNOR2_X1 _09995_ ( .A(_02382_ ), .B(_02383_ ), .ZN(_02384_ ) );
AND3_X1 _09996_ ( .A1(_02336_ ), .A2(_02361_ ), .A3(_02384_ ), .ZN(_02385_ ) );
OR2_X1 _09997_ ( .A1(_02118_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02386_ ) );
OAI211_X1 _09998_ ( .A(_02386_ ), .B(_02108_ ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02387_ ) );
OR2_X1 _09999_ ( .A1(_02118_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02388_ ) );
OAI211_X1 _10000_ ( .A(_02388_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02389_ ) );
NAND3_X1 _10001_ ( .A1(_02387_ ), .A2(_02389_ ), .A3(_02283_ ), .ZN(_02390_ ) );
MUX2_X1 _10002_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02391_ ) );
MUX2_X1 _10003_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02392_ ) );
MUX2_X1 _10004_ ( .A(_02391_ ), .B(_02392_ ), .S(_02277_ ), .Z(_02393_ ) );
OAI211_X1 _10005_ ( .A(fanout_net_26 ), .B(_02390_ ), .C1(_02393_ ), .C2(_02102_ ), .ZN(_02394_ ) );
OR2_X1 _10006_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02395_ ) );
OAI211_X1 _10007_ ( .A(_02395_ ), .B(_02277_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02396_ ) );
NOR2_X1 _10008_ ( .A1(_02119_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02397_ ) );
OAI21_X1 _10009_ ( .A(fanout_net_23 ), .B1(fanout_net_16 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02398_ ) );
OAI211_X1 _10010_ ( .A(_02396_ ), .B(_02283_ ), .C1(_02397_ ), .C2(_02398_ ), .ZN(_02399_ ) );
MUX2_X1 _10011_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02400_ ) );
MUX2_X1 _10012_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02401_ ) );
MUX2_X1 _10013_ ( .A(_02400_ ), .B(_02401_ ), .S(_02287_ ), .Z(_02402_ ) );
OAI211_X1 _10014_ ( .A(_02097_ ), .B(_02399_ ), .C1(_02402_ ), .C2(_02290_ ), .ZN(_02403_ ) );
OAI211_X1 _10015_ ( .A(_02394_ ), .B(_02403_ ), .C1(_02301_ ), .C2(_02167_ ), .ZN(_02404_ ) );
OR4_X1 _10016_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02331_ ), .A3(_02166_ ), .A4(_02305_ ), .ZN(_02405_ ) );
NAND2_X2 _10017_ ( .A1(_02404_ ), .A2(_02405_ ), .ZN(_02406_ ) );
XOR2_X1 _10018_ ( .A(_02406_ ), .B(\ID_EX_imm [18] ), .Z(_02407_ ) );
OR2_X1 _10019_ ( .A1(_02319_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02408_ ) );
OAI211_X1 _10020_ ( .A(_02408_ ), .B(_02287_ ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02409_ ) );
OR2_X1 _10021_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02410_ ) );
OAI211_X1 _10022_ ( .A(_02410_ ), .B(fanout_net_24 ), .C1(_02320_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02411_ ) );
NAND3_X1 _10023_ ( .A1(_02409_ ), .A2(_02101_ ), .A3(_02411_ ), .ZN(_02412_ ) );
MUX2_X1 _10024_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02413_ ) );
MUX2_X1 _10025_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02414_ ) );
BUF_X4 _10026_ ( .A(_02105_ ), .Z(_02415_ ) );
BUF_X4 _10027_ ( .A(_02415_ ), .Z(_02416_ ) );
MUX2_X1 _10028_ ( .A(_02413_ ), .B(_02414_ ), .S(_02416_ ), .Z(_02417_ ) );
OAI211_X1 _10029_ ( .A(fanout_net_26 ), .B(_02412_ ), .C1(_02417_ ), .C2(_02290_ ), .ZN(_02418_ ) );
OR2_X1 _10030_ ( .A1(_02319_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02419_ ) );
OAI211_X1 _10031_ ( .A(_02419_ ), .B(_02416_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02420_ ) );
OR2_X1 _10032_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02421_ ) );
BUF_X4 _10033_ ( .A(_02117_ ), .Z(_02422_ ) );
OAI211_X1 _10034_ ( .A(_02421_ ), .B(fanout_net_24 ), .C1(_02422_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02423_ ) );
NAND3_X1 _10035_ ( .A1(_02420_ ), .A2(_02101_ ), .A3(_02423_ ), .ZN(_02424_ ) );
MUX2_X1 _10036_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02425_ ) );
MUX2_X1 _10037_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02426_ ) );
MUX2_X1 _10038_ ( .A(_02425_ ), .B(_02426_ ), .S(_02416_ ), .Z(_02427_ ) );
OAI211_X1 _10039_ ( .A(_02097_ ), .B(_02424_ ), .C1(_02427_ ), .C2(_02290_ ), .ZN(_02428_ ) );
OAI211_X1 _10040_ ( .A(_02418_ ), .B(_02428_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02429_ ) );
INV_X1 _10041_ ( .A(\ID_EX_imm [19] ), .ZN(_02430_ ) );
OR4_X1 _10042_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02162_ ), .A3(_02147_ ), .A4(_02305_ ), .ZN(_02431_ ) );
AND3_X1 _10043_ ( .A1(_02429_ ), .A2(_02430_ ), .A3(_02431_ ), .ZN(_02432_ ) );
AOI21_X1 _10044_ ( .A(_02430_ ), .B1(_02429_ ), .B2(_02431_ ), .ZN(_02433_ ) );
NOR2_X1 _10045_ ( .A1(_02432_ ), .A2(_02433_ ), .ZN(_02434_ ) );
AND2_X1 _10046_ ( .A1(_02407_ ), .A2(_02434_ ), .ZN(_02435_ ) );
BUF_X2 _10047_ ( .A(_02116_ ), .Z(_02436_ ) );
OR2_X1 _10048_ ( .A1(_02436_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02437_ ) );
OAI211_X1 _10049_ ( .A(_02437_ ), .B(fanout_net_24 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02438_ ) );
OR2_X1 _10050_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02439_ ) );
OAI211_X1 _10051_ ( .A(_02439_ ), .B(_02107_ ), .C1(_02422_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02440_ ) );
NAND3_X1 _10052_ ( .A1(_02438_ ), .A2(fanout_net_25 ), .A3(_02440_ ), .ZN(_02441_ ) );
MUX2_X1 _10053_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02442_ ) );
MUX2_X1 _10054_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02443_ ) );
MUX2_X1 _10055_ ( .A(_02442_ ), .B(_02443_ ), .S(_02107_ ), .Z(_02444_ ) );
OAI211_X1 _10056_ ( .A(_02096_ ), .B(_02441_ ), .C1(_02444_ ), .C2(fanout_net_25 ), .ZN(_02445_ ) );
NOR2_X1 _10057_ ( .A1(_02118_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02446_ ) );
OAI21_X1 _10058_ ( .A(fanout_net_24 ), .B1(fanout_net_17 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02447_ ) );
NOR2_X1 _10059_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02448_ ) );
OAI21_X1 _10060_ ( .A(_02107_ ), .B1(_02118_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02449_ ) );
OAI221_X1 _10061_ ( .A(_02289_ ), .B1(_02446_ ), .B2(_02447_ ), .C1(_02448_ ), .C2(_02449_ ), .ZN(_02450_ ) );
MUX2_X1 _10062_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02451_ ) );
MUX2_X1 _10063_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02452_ ) );
MUX2_X1 _10064_ ( .A(_02451_ ), .B(_02452_ ), .S(fanout_net_24 ), .Z(_02453_ ) );
OAI211_X1 _10065_ ( .A(fanout_net_26 ), .B(_02450_ ), .C1(_02453_ ), .C2(_02283_ ), .ZN(_02454_ ) );
OAI211_X1 _10066_ ( .A(_02445_ ), .B(_02454_ ), .C1(_02139_ ), .C2(_02166_ ), .ZN(_02455_ ) );
CLKBUF_X2 _10067_ ( .A(_02161_ ), .Z(_02456_ ) );
OR4_X1 _10068_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02456_ ), .A3(_02165_ ), .A4(_02169_ ), .ZN(_02457_ ) );
NAND2_X2 _10069_ ( .A1(_02455_ ), .A2(_02457_ ), .ZN(_02458_ ) );
XOR2_X1 _10070_ ( .A(_02458_ ), .B(\ID_EX_imm [17] ), .Z(_02459_ ) );
OR2_X1 _10071_ ( .A1(_02279_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02460_ ) );
OAI211_X1 _10072_ ( .A(_02460_ ), .B(fanout_net_24 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02461_ ) );
OR2_X1 _10073_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02462_ ) );
OAI211_X1 _10074_ ( .A(_02462_ ), .B(_02108_ ), .C1(_02119_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02463_ ) );
NAND3_X1 _10075_ ( .A1(_02461_ ), .A2(_02102_ ), .A3(_02463_ ), .ZN(_02464_ ) );
MUX2_X1 _10076_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02465_ ) );
MUX2_X1 _10077_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02466_ ) );
MUX2_X1 _10078_ ( .A(_02465_ ), .B(_02466_ ), .S(_02108_ ), .Z(_02467_ ) );
OAI211_X1 _10079_ ( .A(_02098_ ), .B(_02464_ ), .C1(_02467_ ), .C2(_02102_ ), .ZN(_02468_ ) );
OR2_X1 _10080_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02469_ ) );
OAI211_X1 _10081_ ( .A(_02469_ ), .B(fanout_net_24 ), .C1(_02119_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02470_ ) );
OR2_X1 _10082_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02471_ ) );
OAI211_X1 _10083_ ( .A(_02471_ ), .B(_02108_ ), .C1(_02119_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02472_ ) );
NAND3_X1 _10084_ ( .A1(_02470_ ), .A2(_02472_ ), .A3(fanout_net_25 ), .ZN(_02473_ ) );
MUX2_X1 _10085_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02474_ ) );
MUX2_X1 _10086_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02475_ ) );
MUX2_X1 _10087_ ( .A(_02474_ ), .B(_02475_ ), .S(fanout_net_24 ), .Z(_02476_ ) );
OAI211_X1 _10088_ ( .A(fanout_net_26 ), .B(_02473_ ), .C1(_02476_ ), .C2(fanout_net_25 ), .ZN(_02477_ ) );
OAI211_X1 _10089_ ( .A(_02468_ ), .B(_02477_ ), .C1(_02195_ ), .C2(_02167_ ), .ZN(_02478_ ) );
OR4_X1 _10090_ ( .A1(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02163_ ), .A3(_02355_ ), .A4(_02170_ ), .ZN(_02479_ ) );
NAND2_X2 _10091_ ( .A1(_02478_ ), .A2(_02479_ ), .ZN(_02480_ ) );
INV_X1 _10092_ ( .A(\ID_EX_imm [16] ), .ZN(_02481_ ) );
XNOR2_X1 _10093_ ( .A(_02480_ ), .B(_02481_ ), .ZN(_02482_ ) );
AND3_X1 _10094_ ( .A1(_02435_ ), .A2(_02459_ ), .A3(_02482_ ), .ZN(_02483_ ) );
OR2_X1 _10095_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02484_ ) );
OAI211_X1 _10096_ ( .A(_02484_ ), .B(_02106_ ), .C1(_02436_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02485_ ) );
OR2_X1 _10097_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02486_ ) );
OAI211_X1 _10098_ ( .A(_02486_ ), .B(fanout_net_24 ), .C1(_02117_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02487_ ) );
NAND3_X1 _10099_ ( .A1(_02485_ ), .A2(_02487_ ), .A3(_02099_ ), .ZN(_02488_ ) );
MUX2_X1 _10100_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02489_ ) );
MUX2_X1 _10101_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02490_ ) );
MUX2_X1 _10102_ ( .A(_02489_ ), .B(_02490_ ), .S(_02106_ ), .Z(_02491_ ) );
OAI211_X1 _10103_ ( .A(fanout_net_26 ), .B(_02488_ ), .C1(_02491_ ), .C2(_02100_ ), .ZN(_02492_ ) );
MUX2_X1 _10104_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02493_ ) );
AND2_X1 _10105_ ( .A1(_02493_ ), .A2(fanout_net_24 ), .ZN(_02494_ ) );
MUX2_X1 _10106_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02495_ ) );
AOI211_X1 _10107_ ( .A(fanout_net_25 ), .B(_02494_ ), .C1(_02107_ ), .C2(_02495_ ), .ZN(_02496_ ) );
MUX2_X1 _10108_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02497_ ) );
MUX2_X1 _10109_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02498_ ) );
MUX2_X1 _10110_ ( .A(_02497_ ), .B(_02498_ ), .S(_02106_ ), .Z(_02499_ ) );
OAI21_X1 _10111_ ( .A(_02095_ ), .B1(_02499_ ), .B2(_02099_ ), .ZN(_02500_ ) );
OAI221_X1 _10112_ ( .A(_02492_ ), .B1(_02496_ ), .B2(_02500_ ), .C1(_02138_ ), .C2(_02165_ ), .ZN(_02501_ ) );
OR4_X4 _10113_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02161_ ), .A3(_02146_ ), .A4(_02169_ ), .ZN(_02502_ ) );
NAND2_X2 _10114_ ( .A1(_02501_ ), .A2(_02502_ ), .ZN(_02503_ ) );
XNOR2_X1 _10115_ ( .A(_02503_ ), .B(\ID_EX_imm [15] ), .ZN(_02504_ ) );
OR2_X1 _10116_ ( .A1(_02116_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02505_ ) );
OAI211_X1 _10117_ ( .A(_02505_ ), .B(_02415_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02506_ ) );
OR2_X1 _10118_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02507_ ) );
OAI211_X1 _10119_ ( .A(_02507_ ), .B(fanout_net_24 ), .C1(_02436_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02508_ ) );
NAND3_X1 _10120_ ( .A1(_02506_ ), .A2(_02100_ ), .A3(_02508_ ), .ZN(_02509_ ) );
MUX2_X1 _10121_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02510_ ) );
MUX2_X1 _10122_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02511_ ) );
MUX2_X1 _10123_ ( .A(_02510_ ), .B(_02511_ ), .S(_02106_ ), .Z(_02512_ ) );
OAI211_X1 _10124_ ( .A(_02096_ ), .B(_02509_ ), .C1(_02512_ ), .C2(_02289_ ), .ZN(_02513_ ) );
OR2_X1 _10125_ ( .A1(_02116_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02514_ ) );
OAI211_X1 _10126_ ( .A(_02514_ ), .B(fanout_net_24 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02515_ ) );
OR2_X1 _10127_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02516_ ) );
OAI211_X1 _10128_ ( .A(_02516_ ), .B(_02106_ ), .C1(_02436_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02517_ ) );
NAND3_X1 _10129_ ( .A1(_02515_ ), .A2(fanout_net_25 ), .A3(_02517_ ), .ZN(_02518_ ) );
MUX2_X1 _10130_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02519_ ) );
MUX2_X1 _10131_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02520_ ) );
MUX2_X1 _10132_ ( .A(_02519_ ), .B(_02520_ ), .S(fanout_net_24 ), .Z(_02521_ ) );
OAI211_X1 _10133_ ( .A(fanout_net_26 ), .B(_02518_ ), .C1(_02521_ ), .C2(fanout_net_25 ), .ZN(_02522_ ) );
OAI211_X1 _10134_ ( .A(_02513_ ), .B(_02522_ ), .C1(_02139_ ), .C2(_02147_ ), .ZN(_02523_ ) );
OR4_X4 _10135_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02303_ ), .A3(_02165_ ), .A4(_02169_ ), .ZN(_02524_ ) );
NAND2_X2 _10136_ ( .A1(_02523_ ), .A2(_02524_ ), .ZN(_02525_ ) );
BUF_X4 _10137_ ( .A(_02525_ ), .Z(_02526_ ) );
INV_X1 _10138_ ( .A(\ID_EX_imm [14] ), .ZN(_02527_ ) );
XNOR2_X1 _10139_ ( .A(_02526_ ), .B(_02527_ ), .ZN(_02528_ ) );
INV_X1 _10140_ ( .A(_02528_ ), .ZN(_02529_ ) );
OR2_X1 _10141_ ( .A1(_02504_ ), .A2(_02529_ ), .ZN(_02530_ ) );
OR2_X1 _10142_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02531_ ) );
OAI211_X1 _10143_ ( .A(_02531_ ), .B(_02276_ ), .C1(_02118_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02532_ ) );
OR2_X1 _10144_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02533_ ) );
OAI211_X1 _10145_ ( .A(_02533_ ), .B(fanout_net_24 ), .C1(_02278_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02534_ ) );
NAND3_X1 _10146_ ( .A1(_02532_ ), .A2(_02534_ ), .A3(_02100_ ), .ZN(_02535_ ) );
MUX2_X1 _10147_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02536_ ) );
MUX2_X1 _10148_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02537_ ) );
MUX2_X1 _10149_ ( .A(_02536_ ), .B(_02537_ ), .S(_02276_ ), .Z(_02538_ ) );
OAI211_X1 _10150_ ( .A(fanout_net_26 ), .B(_02535_ ), .C1(_02538_ ), .C2(_02101_ ), .ZN(_02539_ ) );
OR2_X1 _10151_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02540_ ) );
OAI211_X1 _10152_ ( .A(_02540_ ), .B(_02276_ ), .C1(_02118_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02541_ ) );
OR2_X1 _10153_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02542_ ) );
OAI211_X1 _10154_ ( .A(_02542_ ), .B(fanout_net_24 ), .C1(_02278_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02543_ ) );
NAND3_X1 _10155_ ( .A1(_02541_ ), .A2(_02543_ ), .A3(_02100_ ), .ZN(_02544_ ) );
MUX2_X1 _10156_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02545_ ) );
MUX2_X1 _10157_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02546_ ) );
MUX2_X1 _10158_ ( .A(_02545_ ), .B(_02546_ ), .S(_02415_ ), .Z(_02547_ ) );
OAI211_X1 _10159_ ( .A(_02096_ ), .B(_02544_ ), .C1(_02547_ ), .C2(_02101_ ), .ZN(_02548_ ) );
OAI211_X1 _10160_ ( .A(_02539_ ), .B(_02548_ ), .C1(_02139_ ), .C2(_02166_ ), .ZN(_02549_ ) );
OR4_X1 _10161_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02303_ ), .A3(_02165_ ), .A4(_02169_ ), .ZN(_02550_ ) );
NAND2_X1 _10162_ ( .A1(_02549_ ), .A2(_02550_ ), .ZN(_02551_ ) );
BUF_X4 _10163_ ( .A(_02551_ ), .Z(_02552_ ) );
XNOR2_X1 _10164_ ( .A(_02552_ ), .B(\ID_EX_imm [13] ), .ZN(_02553_ ) );
OR2_X1 _10165_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02554_ ) );
OAI211_X1 _10166_ ( .A(_02554_ ), .B(_02107_ ), .C1(_02422_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02555_ ) );
OR2_X1 _10167_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02556_ ) );
OAI211_X1 _10168_ ( .A(_02556_ ), .B(fanout_net_24 ), .C1(_02118_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02557_ ) );
NAND3_X1 _10169_ ( .A1(_02555_ ), .A2(_02557_ ), .A3(_02289_ ), .ZN(_02558_ ) );
MUX2_X1 _10170_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02559_ ) );
MUX2_X1 _10171_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02560_ ) );
MUX2_X1 _10172_ ( .A(_02559_ ), .B(_02560_ ), .S(_02276_ ), .Z(_02561_ ) );
OAI211_X1 _10173_ ( .A(_02096_ ), .B(_02558_ ), .C1(_02561_ ), .C2(_02101_ ), .ZN(_02562_ ) );
OR2_X1 _10174_ ( .A1(_02117_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02563_ ) );
OAI211_X1 _10175_ ( .A(_02563_ ), .B(fanout_net_24 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02564_ ) );
OR2_X1 _10176_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02565_ ) );
OAI211_X1 _10177_ ( .A(_02565_ ), .B(_02276_ ), .C1(_02118_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02566_ ) );
NAND3_X1 _10178_ ( .A1(_02564_ ), .A2(fanout_net_25 ), .A3(_02566_ ), .ZN(_02567_ ) );
MUX2_X1 _10179_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02568_ ) );
MUX2_X1 _10180_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02569_ ) );
MUX2_X1 _10181_ ( .A(_02568_ ), .B(_02569_ ), .S(fanout_net_24 ), .Z(_02570_ ) );
OAI211_X1 _10182_ ( .A(fanout_net_26 ), .B(_02567_ ), .C1(_02570_ ), .C2(fanout_net_25 ), .ZN(_02571_ ) );
OAI211_X1 _10183_ ( .A(_02562_ ), .B(_02571_ ), .C1(_02139_ ), .C2(_02166_ ), .ZN(_02572_ ) );
OR4_X1 _10184_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02456_ ), .A3(_02165_ ), .A4(_02169_ ), .ZN(_02573_ ) );
NAND2_X4 _10185_ ( .A1(_02572_ ), .A2(_02573_ ), .ZN(_02574_ ) );
INV_X1 _10186_ ( .A(\ID_EX_imm [12] ), .ZN(_02575_ ) );
XNOR2_X1 _10187_ ( .A(_02574_ ), .B(_02575_ ), .ZN(_02576_ ) );
INV_X1 _10188_ ( .A(_02576_ ), .ZN(_02577_ ) );
OR3_X1 _10189_ ( .A1(_02530_ ), .A2(_02553_ ), .A3(_02577_ ), .ZN(_02578_ ) );
OR2_X1 _10190_ ( .A1(_02278_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02579_ ) );
OAI211_X1 _10191_ ( .A(_02579_ ), .B(_02277_ ), .C1(fanout_net_18 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02580_ ) );
OR2_X1 _10192_ ( .A1(fanout_net_18 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02581_ ) );
OAI211_X1 _10193_ ( .A(_02581_ ), .B(fanout_net_24 ), .C1(_02320_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02582_ ) );
NAND3_X1 _10194_ ( .A1(_02580_ ), .A2(_02283_ ), .A3(_02582_ ), .ZN(_02583_ ) );
MUX2_X1 _10195_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02584_ ) );
MUX2_X1 _10196_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02585_ ) );
MUX2_X1 _10197_ ( .A(_02584_ ), .B(_02585_ ), .S(_02287_ ), .Z(_02586_ ) );
OAI211_X1 _10198_ ( .A(_02097_ ), .B(_02583_ ), .C1(_02586_ ), .C2(_02290_ ), .ZN(_02587_ ) );
OR2_X1 _10199_ ( .A1(_02278_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02588_ ) );
OAI211_X1 _10200_ ( .A(_02588_ ), .B(fanout_net_24 ), .C1(fanout_net_18 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02589_ ) );
OR2_X1 _10201_ ( .A1(fanout_net_18 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02590_ ) );
OAI211_X1 _10202_ ( .A(_02590_ ), .B(_02287_ ), .C1(_02320_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02591_ ) );
NAND3_X1 _10203_ ( .A1(_02589_ ), .A2(fanout_net_25 ), .A3(_02591_ ), .ZN(_02592_ ) );
MUX2_X1 _10204_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02593_ ) );
MUX2_X1 _10205_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02594_ ) );
MUX2_X1 _10206_ ( .A(_02593_ ), .B(_02594_ ), .S(fanout_net_24 ), .Z(_02595_ ) );
OAI211_X1 _10207_ ( .A(fanout_net_26 ), .B(_02592_ ), .C1(_02595_ ), .C2(fanout_net_25 ), .ZN(_02596_ ) );
OAI211_X1 _10208_ ( .A(_02587_ ), .B(_02596_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02597_ ) );
OR4_X1 _10209_ ( .A1(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02304_ ), .A3(_02147_ ), .A4(_02305_ ), .ZN(_02598_ ) );
NAND2_X1 _10210_ ( .A1(_02597_ ), .A2(_02598_ ), .ZN(_02599_ ) );
BUF_X4 _10211_ ( .A(_02599_ ), .Z(_02600_ ) );
INV_X1 _10212_ ( .A(\ID_EX_imm [8] ), .ZN(_02601_ ) );
XNOR2_X1 _10213_ ( .A(_02600_ ), .B(_02601_ ), .ZN(_02602_ ) );
INV_X1 _10214_ ( .A(_02602_ ), .ZN(_02603_ ) );
OR2_X1 _10215_ ( .A1(_02117_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02604_ ) );
OAI211_X1 _10216_ ( .A(_02604_ ), .B(_02415_ ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02605_ ) );
OR2_X1 _10217_ ( .A1(_02117_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02606_ ) );
OAI211_X1 _10218_ ( .A(_02606_ ), .B(fanout_net_24 ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02607_ ) );
NAND3_X1 _10219_ ( .A1(_02605_ ), .A2(_02607_ ), .A3(_02100_ ), .ZN(_02608_ ) );
MUX2_X1 _10220_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02609_ ) );
MUX2_X1 _10221_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02610_ ) );
MUX2_X1 _10222_ ( .A(_02609_ ), .B(_02610_ ), .S(_02415_ ), .Z(_02611_ ) );
OAI211_X1 _10223_ ( .A(fanout_net_26 ), .B(_02608_ ), .C1(_02611_ ), .C2(_02289_ ), .ZN(_02612_ ) );
OR2_X1 _10224_ ( .A1(_02117_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02613_ ) );
OAI211_X1 _10225_ ( .A(_02613_ ), .B(fanout_net_24 ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02614_ ) );
OR2_X1 _10226_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02615_ ) );
OAI211_X1 _10227_ ( .A(_02615_ ), .B(_02415_ ), .C1(_02436_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02616_ ) );
NAND3_X1 _10228_ ( .A1(_02614_ ), .A2(_02100_ ), .A3(_02616_ ), .ZN(_02617_ ) );
MUX2_X1 _10229_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02618_ ) );
MUX2_X1 _10230_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02619_ ) );
MUX2_X1 _10231_ ( .A(_02618_ ), .B(_02619_ ), .S(_02106_ ), .Z(_02620_ ) );
OAI211_X1 _10232_ ( .A(_02096_ ), .B(_02617_ ), .C1(_02620_ ), .C2(_02289_ ), .ZN(_02621_ ) );
OAI211_X1 _10233_ ( .A(_02612_ ), .B(_02621_ ), .C1(_02139_ ), .C2(_02147_ ), .ZN(_02622_ ) );
OR4_X1 _10234_ ( .A1(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02303_ ), .A3(_02165_ ), .A4(_02169_ ), .ZN(_02623_ ) );
NAND2_X2 _10235_ ( .A1(_02622_ ), .A2(_02623_ ), .ZN(_02624_ ) );
XNOR2_X1 _10236_ ( .A(_02624_ ), .B(\ID_EX_imm [9] ), .ZN(_02625_ ) );
NOR2_X1 _10237_ ( .A1(_02603_ ), .A2(_02625_ ), .ZN(_02626_ ) );
OR2_X1 _10238_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02627_ ) );
OAI211_X1 _10239_ ( .A(_02627_ ), .B(_02416_ ), .C1(_02320_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02628_ ) );
OR2_X1 _10240_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02629_ ) );
OAI211_X1 _10241_ ( .A(_02629_ ), .B(fanout_net_24 ), .C1(_02422_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02630_ ) );
NAND3_X1 _10242_ ( .A1(_02628_ ), .A2(_02630_ ), .A3(_02101_ ), .ZN(_02631_ ) );
MUX2_X1 _10243_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02632_ ) );
MUX2_X1 _10244_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02633_ ) );
MUX2_X1 _10245_ ( .A(_02632_ ), .B(_02633_ ), .S(_02416_ ), .Z(_02634_ ) );
OAI211_X1 _10246_ ( .A(fanout_net_26 ), .B(_02631_ ), .C1(_02634_ ), .C2(_02290_ ), .ZN(_02635_ ) );
OR2_X1 _10247_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02636_ ) );
OAI211_X1 _10248_ ( .A(_02636_ ), .B(_02416_ ), .C1(_02422_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02637_ ) );
NOR2_X1 _10249_ ( .A1(_02320_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02638_ ) );
OAI21_X1 _10250_ ( .A(fanout_net_24 ), .B1(fanout_net_19 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02639_ ) );
OAI211_X1 _10251_ ( .A(_02637_ ), .B(_02289_ ), .C1(_02638_ ), .C2(_02639_ ), .ZN(_02640_ ) );
MUX2_X1 _10252_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02641_ ) );
MUX2_X1 _10253_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02642_ ) );
MUX2_X1 _10254_ ( .A(_02641_ ), .B(_02642_ ), .S(_02416_ ), .Z(_02643_ ) );
OAI211_X1 _10255_ ( .A(_02097_ ), .B(_02640_ ), .C1(_02643_ ), .C2(_02290_ ), .ZN(_02644_ ) );
OAI211_X1 _10256_ ( .A(_02635_ ), .B(_02644_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02645_ ) );
OR4_X1 _10257_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02162_ ), .A3(_02147_ ), .A4(_02305_ ), .ZN(_02646_ ) );
NAND2_X2 _10258_ ( .A1(_02645_ ), .A2(_02646_ ), .ZN(_02647_ ) );
INV_X1 _10259_ ( .A(\ID_EX_imm [10] ), .ZN(_02648_ ) );
XNOR2_X1 _10260_ ( .A(_02647_ ), .B(_02648_ ), .ZN(_02649_ ) );
OR2_X1 _10261_ ( .A1(_02278_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02650_ ) );
OAI211_X1 _10262_ ( .A(_02650_ ), .B(fanout_net_24 ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02651_ ) );
OR2_X1 _10263_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02652_ ) );
OAI211_X1 _10264_ ( .A(_02652_ ), .B(_02287_ ), .C1(_02320_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02653_ ) );
NAND3_X1 _10265_ ( .A1(_02651_ ), .A2(_02283_ ), .A3(_02653_ ), .ZN(_02654_ ) );
MUX2_X1 _10266_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02655_ ) );
MUX2_X1 _10267_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02656_ ) );
MUX2_X1 _10268_ ( .A(_02655_ ), .B(_02656_ ), .S(_02416_ ), .Z(_02657_ ) );
OAI211_X1 _10269_ ( .A(_02097_ ), .B(_02654_ ), .C1(_02657_ ), .C2(_02290_ ), .ZN(_02658_ ) );
OR2_X1 _10270_ ( .A1(_02319_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02659_ ) );
OAI211_X1 _10271_ ( .A(_02659_ ), .B(fanout_net_24 ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02660_ ) );
OR2_X1 _10272_ ( .A1(_02319_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02661_ ) );
OAI211_X1 _10273_ ( .A(_02661_ ), .B(_02287_ ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02662_ ) );
NAND3_X1 _10274_ ( .A1(_02660_ ), .A2(_02662_ ), .A3(fanout_net_25 ), .ZN(_02663_ ) );
MUX2_X1 _10275_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02664_ ) );
MUX2_X1 _10276_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02665_ ) );
MUX2_X1 _10277_ ( .A(_02664_ ), .B(_02665_ ), .S(fanout_net_24 ), .Z(_02666_ ) );
OAI211_X1 _10278_ ( .A(fanout_net_26 ), .B(_02663_ ), .C1(_02666_ ), .C2(fanout_net_25 ), .ZN(_02667_ ) );
OAI211_X1 _10279_ ( .A(_02658_ ), .B(_02667_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02668_ ) );
OR4_X4 _10280_ ( .A1(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A2(_02304_ ), .A3(_02147_ ), .A4(_02305_ ), .ZN(_02669_ ) );
NAND2_X2 _10281_ ( .A1(_02668_ ), .A2(_02669_ ), .ZN(_02670_ ) );
INV_X1 _10282_ ( .A(\ID_EX_imm [11] ), .ZN(_02671_ ) );
XNOR2_X1 _10283_ ( .A(_02670_ ), .B(_02671_ ), .ZN(_02672_ ) );
AND2_X1 _10284_ ( .A1(_02649_ ), .A2(_02672_ ), .ZN(_02673_ ) );
NAND2_X1 _10285_ ( .A1(_02626_ ), .A2(_02673_ ), .ZN(_02674_ ) );
OR2_X1 _10286_ ( .A1(_02116_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02675_ ) );
OAI211_X1 _10287_ ( .A(_02675_ ), .B(_02415_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02676_ ) );
OR2_X1 _10288_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02677_ ) );
OAI211_X1 _10289_ ( .A(_02677_ ), .B(fanout_net_24 ), .C1(_02436_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02678_ ) );
NAND3_X1 _10290_ ( .A1(_02676_ ), .A2(_02099_ ), .A3(_02678_ ), .ZN(_02679_ ) );
MUX2_X1 _10291_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02680_ ) );
MUX2_X1 _10292_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02681_ ) );
MUX2_X1 _10293_ ( .A(_02680_ ), .B(_02681_ ), .S(_02106_ ), .Z(_02682_ ) );
OAI211_X1 _10294_ ( .A(_02095_ ), .B(_02679_ ), .C1(_02682_ ), .C2(_02289_ ), .ZN(_02683_ ) );
OR2_X1 _10295_ ( .A1(_02116_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02684_ ) );
OAI211_X1 _10296_ ( .A(_02684_ ), .B(_02106_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02685_ ) );
OR2_X1 _10297_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02686_ ) );
OAI211_X1 _10298_ ( .A(_02686_ ), .B(fanout_net_24 ), .C1(_02436_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02687_ ) );
NAND3_X1 _10299_ ( .A1(_02685_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02687_ ), .ZN(_02688_ ) );
MUX2_X1 _10300_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02689_ ) );
MUX2_X1 _10301_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02690_ ) );
MUX2_X1 _10302_ ( .A(_02689_ ), .B(_02690_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02691_ ) );
OAI211_X1 _10303_ ( .A(fanout_net_26 ), .B(_02688_ ), .C1(_02691_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02692_ ) );
OAI211_X1 _10304_ ( .A(_02683_ ), .B(_02692_ ), .C1(_02139_ ), .C2(_02147_ ), .ZN(_02693_ ) );
OR4_X1 _10305_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02161_ ), .A3(_02146_ ), .A4(_02169_ ), .ZN(_02694_ ) );
NAND2_X2 _10306_ ( .A1(_02693_ ), .A2(_02694_ ), .ZN(_02695_ ) );
NAND2_X1 _10307_ ( .A1(_02695_ ), .A2(\ID_EX_imm [2] ), .ZN(_02696_ ) );
OR2_X1 _10308_ ( .A1(_02115_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02697_ ) );
OAI211_X1 _10309_ ( .A(_02697_ ), .B(_02105_ ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02698_ ) );
OR2_X1 _10310_ ( .A1(_02115_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02699_ ) );
OAI211_X1 _10311_ ( .A(_02699_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02700_ ) );
NAND3_X1 _10312_ ( .A1(_02698_ ), .A2(_02700_ ), .A3(_02099_ ), .ZN(_02701_ ) );
MUX2_X1 _10313_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02702_ ) );
MUX2_X1 _10314_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02703_ ) );
MUX2_X1 _10315_ ( .A(_02702_ ), .B(_02703_ ), .S(_02105_ ), .Z(_02704_ ) );
OAI211_X1 _10316_ ( .A(_02095_ ), .B(_02701_ ), .C1(_02704_ ), .C2(_02099_ ), .ZN(_02705_ ) );
OR2_X1 _10317_ ( .A1(_02115_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02706_ ) );
OAI211_X1 _10318_ ( .A(_02706_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02707_ ) );
OR2_X1 _10319_ ( .A1(_02115_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02708_ ) );
OAI211_X1 _10320_ ( .A(_02708_ ), .B(_02105_ ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02709_ ) );
NAND3_X1 _10321_ ( .A1(_02707_ ), .A2(_02709_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02710_ ) );
MUX2_X1 _10322_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02711_ ) );
MUX2_X1 _10323_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02712_ ) );
MUX2_X1 _10324_ ( .A(_02711_ ), .B(_02712_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02713_ ) );
OAI211_X1 _10325_ ( .A(fanout_net_26 ), .B(_02710_ ), .C1(_02713_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02714_ ) );
OAI211_X1 _10326_ ( .A(_02705_ ), .B(_02714_ ), .C1(_02138_ ), .C2(_02146_ ), .ZN(_02715_ ) );
OR4_X1 _10327_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02131_ ), .A3(_02146_ ), .A4(_02137_ ), .ZN(_02716_ ) );
NAND2_X2 _10328_ ( .A1(_02715_ ), .A2(_02716_ ), .ZN(_02717_ ) );
INV_X1 _10329_ ( .A(\ID_EX_imm [1] ), .ZN(_02718_ ) );
XNOR2_X1 _10330_ ( .A(_02717_ ), .B(_02718_ ), .ZN(_02719_ ) );
INV_X1 _10331_ ( .A(\ID_EX_imm [0] ), .ZN(_02720_ ) );
OR2_X1 _10332_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(fanout_net_20 ), .ZN(_02721_ ) );
OAI211_X1 _10333_ ( .A(_02721_ ), .B(_02105_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_02116_ ), .ZN(_02722_ ) );
OR2_X1 _10334_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02723_ ) );
OAI211_X1 _10335_ ( .A(_02723_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02116_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02724_ ) );
NAND3_X1 _10336_ ( .A1(_02722_ ), .A2(_02724_ ), .A3(_02099_ ), .ZN(_02725_ ) );
MUX2_X1 _10337_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02726_ ) );
MUX2_X1 _10338_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02727_ ) );
MUX2_X1 _10339_ ( .A(_02726_ ), .B(_02727_ ), .S(_02105_ ), .Z(_02728_ ) );
OAI211_X1 _10340_ ( .A(_02095_ ), .B(_02725_ ), .C1(_02728_ ), .C2(_02099_ ), .ZN(_02729_ ) );
OR2_X1 _10341_ ( .A1(_02116_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02730_ ) );
OAI211_X1 _10342_ ( .A(_02730_ ), .B(_02105_ ), .C1(fanout_net_20 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02731_ ) );
OR2_X1 _10343_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02732_ ) );
OAI211_X1 _10344_ ( .A(_02732_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02116_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02733_ ) );
NAND3_X1 _10345_ ( .A1(_02731_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02733_ ), .ZN(_02734_ ) );
MUX2_X1 _10346_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02735_ ) );
MUX2_X1 _10347_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02736_ ) );
MUX2_X1 _10348_ ( .A(_02735_ ), .B(_02736_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02737_ ) );
OAI211_X1 _10349_ ( .A(fanout_net_26 ), .B(_02734_ ), .C1(_02737_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02738_ ) );
OAI211_X1 _10350_ ( .A(_02729_ ), .B(_02738_ ), .C1(_02138_ ), .C2(_02146_ ), .ZN(_02739_ ) );
OR4_X1 _10351_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A2(_02131_ ), .A3(_02146_ ), .A4(_02137_ ), .ZN(_02740_ ) );
AOI21_X1 _10352_ ( .A(_02720_ ), .B1(_02739_ ), .B2(_02740_ ), .ZN(_02741_ ) );
AND2_X1 _10353_ ( .A1(_02719_ ), .A2(_02741_ ), .ZN(_02742_ ) );
AOI21_X1 _10354_ ( .A(_02742_ ), .B1(\ID_EX_imm [1] ), .B2(_02717_ ), .ZN(_02743_ ) );
XNOR2_X1 _10355_ ( .A(_02695_ ), .B(\ID_EX_imm [2] ), .ZN(_02744_ ) );
OAI21_X1 _10356_ ( .A(_02696_ ), .B1(_02743_ ), .B2(_02744_ ), .ZN(_02745_ ) );
OR2_X1 _10357_ ( .A1(_02117_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02746_ ) );
OAI211_X1 _10358_ ( .A(_02746_ ), .B(_02276_ ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02747_ ) );
OR2_X1 _10359_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02748_ ) );
OAI211_X1 _10360_ ( .A(_02748_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02118_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02749_ ) );
NAND3_X1 _10361_ ( .A1(_02747_ ), .A2(_02749_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02750_ ) );
MUX2_X1 _10362_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02751_ ) );
MUX2_X1 _10363_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02752_ ) );
MUX2_X1 _10364_ ( .A(_02751_ ), .B(_02752_ ), .S(_02276_ ), .Z(_02753_ ) );
OAI211_X1 _10365_ ( .A(_02096_ ), .B(_02750_ ), .C1(_02753_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02754_ ) );
NOR2_X1 _10366_ ( .A1(_02319_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02755_ ) );
OAI21_X1 _10367_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_20 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02756_ ) );
NOR2_X1 _10368_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02757_ ) );
OAI21_X1 _10369_ ( .A(_02276_ ), .B1(_02319_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02758_ ) );
OAI221_X1 _10370_ ( .A(_02100_ ), .B1(_02755_ ), .B2(_02756_ ), .C1(_02757_ ), .C2(_02758_ ), .ZN(_02759_ ) );
MUX2_X1 _10371_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02760_ ) );
MUX2_X1 _10372_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02761_ ) );
MUX2_X1 _10373_ ( .A(_02760_ ), .B(_02761_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02762_ ) );
OAI211_X1 _10374_ ( .A(fanout_net_26 ), .B(_02759_ ), .C1(_02762_ ), .C2(_02101_ ), .ZN(_02763_ ) );
OAI211_X1 _10375_ ( .A(_02754_ ), .B(_02763_ ), .C1(_02139_ ), .C2(_02166_ ), .ZN(_02764_ ) );
OR4_X1 _10376_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02456_ ), .A3(_02165_ ), .A4(_02169_ ), .ZN(_02765_ ) );
NAND2_X1 _10377_ ( .A1(_02764_ ), .A2(_02765_ ), .ZN(_02766_ ) );
XOR2_X1 _10378_ ( .A(_02766_ ), .B(\ID_EX_imm [3] ), .Z(_02767_ ) );
NAND2_X1 _10379_ ( .A1(_02745_ ), .A2(_02767_ ), .ZN(_02768_ ) );
INV_X1 _10380_ ( .A(_02766_ ), .ZN(_02769_ ) );
OR2_X1 _10381_ ( .A1(_02769_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02770_ ) );
NAND2_X1 _10382_ ( .A1(_02768_ ), .A2(_02770_ ), .ZN(_02771_ ) );
OR2_X1 _10383_ ( .A1(_02436_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02772_ ) );
OAI211_X1 _10384_ ( .A(_02772_ ), .B(_02416_ ), .C1(fanout_net_20 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02773_ ) );
OR2_X1 _10385_ ( .A1(fanout_net_20 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02774_ ) );
OAI211_X1 _10386_ ( .A(_02774_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02422_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02775_ ) );
NAND3_X1 _10387_ ( .A1(_02773_ ), .A2(_02101_ ), .A3(_02775_ ), .ZN(_02776_ ) );
MUX2_X1 _10388_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02777_ ) );
MUX2_X1 _10389_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02778_ ) );
MUX2_X1 _10390_ ( .A(_02777_ ), .B(_02778_ ), .S(_02107_ ), .Z(_02779_ ) );
OAI211_X1 _10391_ ( .A(_02096_ ), .B(_02776_ ), .C1(_02779_ ), .C2(_02283_ ), .ZN(_02780_ ) );
OR2_X1 _10392_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02781_ ) );
OAI211_X1 _10393_ ( .A(_02781_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02422_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02782_ ) );
OR2_X1 _10394_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02783_ ) );
OAI211_X1 _10395_ ( .A(_02783_ ), .B(_02416_ ), .C1(_02422_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02784_ ) );
NAND3_X1 _10396_ ( .A1(_02782_ ), .A2(_02784_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02785_ ) );
MUX2_X1 _10397_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02786_ ) );
MUX2_X1 _10398_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02787_ ) );
MUX2_X1 _10399_ ( .A(_02786_ ), .B(_02787_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02788_ ) );
OAI211_X1 _10400_ ( .A(fanout_net_26 ), .B(_02785_ ), .C1(_02788_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02789_ ) );
OAI211_X1 _10401_ ( .A(_02780_ ), .B(_02789_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02790_ ) );
OR4_X1 _10402_ ( .A1(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02162_ ), .A3(_02147_ ), .A4(_02305_ ), .ZN(_02791_ ) );
NAND2_X2 _10403_ ( .A1(_02790_ ), .A2(_02791_ ), .ZN(_02792_ ) );
INV_X1 _10404_ ( .A(\ID_EX_imm [6] ), .ZN(_02793_ ) );
XNOR2_X1 _10405_ ( .A(_02792_ ), .B(_02793_ ), .ZN(_02794_ ) );
INV_X1 _10406_ ( .A(_02794_ ), .ZN(_02795_ ) );
OR2_X1 _10407_ ( .A1(_02436_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02796_ ) );
OAI211_X1 _10408_ ( .A(_02796_ ), .B(_02107_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02797_ ) );
OR2_X1 _10409_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02798_ ) );
OAI211_X1 _10410_ ( .A(_02798_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02422_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02799_ ) );
NAND3_X1 _10411_ ( .A1(_02797_ ), .A2(_02289_ ), .A3(_02799_ ), .ZN(_02800_ ) );
MUX2_X1 _10412_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02801_ ) );
MUX2_X1 _10413_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02802_ ) );
MUX2_X1 _10414_ ( .A(_02801_ ), .B(_02802_ ), .S(_02107_ ), .Z(_02803_ ) );
OAI211_X1 _10415_ ( .A(_02096_ ), .B(_02800_ ), .C1(_02803_ ), .C2(_02283_ ), .ZN(_02804_ ) );
OR2_X1 _10416_ ( .A1(_02436_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02805_ ) );
OAI211_X1 _10417_ ( .A(_02805_ ), .B(_02107_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02806_ ) );
OR2_X1 _10418_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02807_ ) );
OAI211_X1 _10419_ ( .A(_02807_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02422_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02808_ ) );
NAND3_X1 _10420_ ( .A1(_02806_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02808_ ), .ZN(_02809_ ) );
MUX2_X1 _10421_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02810_ ) );
MUX2_X1 _10422_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02811_ ) );
MUX2_X1 _10423_ ( .A(_02810_ ), .B(_02811_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02812_ ) );
OAI211_X1 _10424_ ( .A(fanout_net_26 ), .B(_02809_ ), .C1(_02812_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02813_ ) );
OAI211_X1 _10425_ ( .A(_02804_ ), .B(_02813_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02814_ ) );
OR4_X1 _10426_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02456_ ), .A3(_02165_ ), .A4(_02305_ ), .ZN(_02815_ ) );
NAND2_X2 _10427_ ( .A1(_02814_ ), .A2(_02815_ ), .ZN(_02816_ ) );
XNOR2_X1 _10428_ ( .A(_02816_ ), .B(\ID_EX_imm [7] ), .ZN(_02817_ ) );
NOR2_X1 _10429_ ( .A1(_02795_ ), .A2(_02817_ ), .ZN(_02818_ ) );
NAND2_X1 _10430_ ( .A1(_02148_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02819_ ) );
OR2_X1 _10431_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02820_ ) );
OAI211_X1 _10432_ ( .A(_02820_ ), .B(_02415_ ), .C1(_02319_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02821_ ) );
INV_X1 _10433_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02822_ ) );
NAND2_X1 _10434_ ( .A1(_02822_ ), .A2(fanout_net_21 ), .ZN(_02823_ ) );
OAI211_X1 _10435_ ( .A(_02823_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02824_ ) );
NAND3_X1 _10436_ ( .A1(_02821_ ), .A2(_02824_ ), .A3(_02100_ ), .ZN(_02825_ ) );
MUX2_X1 _10437_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02826_ ) );
MUX2_X1 _10438_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02827_ ) );
MUX2_X1 _10439_ ( .A(_02826_ ), .B(_02827_ ), .S(_02415_ ), .Z(_02828_ ) );
OAI211_X1 _10440_ ( .A(_02096_ ), .B(_02825_ ), .C1(_02828_ ), .C2(_02289_ ), .ZN(_02829_ ) );
OR2_X1 _10441_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02830_ ) );
OAI211_X1 _10442_ ( .A(_02830_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02319_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02831_ ) );
OR2_X1 _10443_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02832_ ) );
OAI211_X1 _10444_ ( .A(_02832_ ), .B(_02415_ ), .C1(_02319_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02833_ ) );
NAND3_X1 _10445_ ( .A1(_02831_ ), .A2(_02833_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02834_ ) );
MUX2_X1 _10446_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02835_ ) );
MUX2_X1 _10447_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02836_ ) );
MUX2_X1 _10448_ ( .A(_02835_ ), .B(_02836_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02837_ ) );
OAI211_X1 _10449_ ( .A(fanout_net_26 ), .B(_02834_ ), .C1(_02837_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02838_ ) );
NAND2_X1 _10450_ ( .A1(_02829_ ), .A2(_02838_ ), .ZN(_02839_ ) );
OAI21_X1 _10451_ ( .A(_02839_ ), .B1(_02166_ ), .B2(_02139_ ), .ZN(_02840_ ) );
AND2_X2 _10452_ ( .A1(_02819_ ), .A2(_02840_ ), .ZN(_02841_ ) );
XNOR2_X1 _10453_ ( .A(_02841_ ), .B(\ID_EX_imm [5] ), .ZN(_02842_ ) );
OR2_X1 _10454_ ( .A1(_02278_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02843_ ) );
OAI211_X1 _10455_ ( .A(_02843_ ), .B(_02277_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02844_ ) );
OR2_X1 _10456_ ( .A1(_02278_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02845_ ) );
OAI211_X1 _10457_ ( .A(_02845_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02846_ ) );
NAND3_X1 _10458_ ( .A1(_02844_ ), .A2(_02846_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02847_ ) );
MUX2_X1 _10459_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02848_ ) );
MUX2_X1 _10460_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02849_ ) );
MUX2_X1 _10461_ ( .A(_02848_ ), .B(_02849_ ), .S(_02287_ ), .Z(_02850_ ) );
OAI211_X1 _10462_ ( .A(_02097_ ), .B(_02847_ ), .C1(_02850_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02851_ ) );
NOR2_X1 _10463_ ( .A1(_02320_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02852_ ) );
OAI21_X1 _10464_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_21 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02853_ ) );
NOR2_X1 _10465_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02854_ ) );
OAI21_X1 _10466_ ( .A(_02287_ ), .B1(_02320_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02855_ ) );
OAI221_X1 _10467_ ( .A(_02101_ ), .B1(_02852_ ), .B2(_02853_ ), .C1(_02854_ ), .C2(_02855_ ), .ZN(_02856_ ) );
MUX2_X1 _10468_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02857_ ) );
MUX2_X1 _10469_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02858_ ) );
MUX2_X1 _10470_ ( .A(_02857_ ), .B(_02858_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02859_ ) );
OAI211_X1 _10471_ ( .A(fanout_net_26 ), .B(_02856_ ), .C1(_02859_ ), .C2(_02290_ ), .ZN(_02860_ ) );
OAI211_X1 _10472_ ( .A(_02851_ ), .B(_02860_ ), .C1(_02301_ ), .C2(_02355_ ), .ZN(_02861_ ) );
OR4_X1 _10473_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02304_ ), .A3(_02166_ ), .A4(_02305_ ), .ZN(_02862_ ) );
NAND2_X1 _10474_ ( .A1(_02861_ ), .A2(_02862_ ), .ZN(_02863_ ) );
BUF_X4 _10475_ ( .A(_02863_ ), .Z(_02864_ ) );
INV_X1 _10476_ ( .A(\ID_EX_imm [4] ), .ZN(_02865_ ) );
XNOR2_X1 _10477_ ( .A(_02864_ ), .B(_02865_ ), .ZN(_02866_ ) );
INV_X1 _10478_ ( .A(_02866_ ), .ZN(_02867_ ) );
NOR2_X1 _10479_ ( .A1(_02842_ ), .A2(_02867_ ), .ZN(_02868_ ) );
NAND3_X1 _10480_ ( .A1(_02771_ ), .A2(_02818_ ), .A3(_02868_ ), .ZN(_02869_ ) );
INV_X1 _10481_ ( .A(_02792_ ), .ZN(_02870_ ) );
NOR3_X1 _10482_ ( .A1(_02817_ ), .A2(_02793_ ), .A3(_02870_ ), .ZN(_02871_ ) );
AND2_X1 _10483_ ( .A1(_02864_ ), .A2(\ID_EX_imm [4] ), .ZN(_02872_ ) );
INV_X1 _10484_ ( .A(_02872_ ), .ZN(_02873_ ) );
OR2_X1 _10485_ ( .A1(_02842_ ), .A2(_02873_ ), .ZN(_02874_ ) );
INV_X1 _10486_ ( .A(_02841_ ), .ZN(_02875_ ) );
OAI21_X1 _10487_ ( .A(_02874_ ), .B1(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_02875_ ), .ZN(_02876_ ) );
AOI221_X4 _10488_ ( .A(_02871_ ), .B1(\ID_EX_imm [7] ), .B2(_02816_ ), .C1(_02876_ ), .C2(_02818_ ), .ZN(_02877_ ) );
AOI211_X1 _10489_ ( .A(_02578_ ), .B(_02674_ ), .C1(_02869_ ), .C2(_02877_ ), .ZN(_02878_ ) );
AND2_X1 _10490_ ( .A1(_02647_ ), .A2(\ID_EX_imm [10] ), .ZN(_02879_ ) );
AND2_X1 _10491_ ( .A1(_02672_ ), .A2(_02879_ ), .ZN(_02880_ ) );
AOI21_X1 _10492_ ( .A(_02880_ ), .B1(\ID_EX_imm [11] ), .B2(_02670_ ), .ZN(_02881_ ) );
NAND2_X1 _10493_ ( .A1(_02624_ ), .A2(\ID_EX_imm [9] ), .ZN(_02882_ ) );
NAND2_X1 _10494_ ( .A1(_02600_ ), .A2(\ID_EX_imm [8] ), .ZN(_02883_ ) );
OAI21_X1 _10495_ ( .A(_02882_ ), .B1(_02625_ ), .B2(_02883_ ), .ZN(_02884_ ) );
NAND2_X1 _10496_ ( .A1(_02673_ ), .A2(_02884_ ), .ZN(_02885_ ) );
AND2_X1 _10497_ ( .A1(_02881_ ), .A2(_02885_ ), .ZN(_02886_ ) );
OR2_X1 _10498_ ( .A1(_02886_ ), .A2(_02578_ ), .ZN(_02887_ ) );
NAND2_X1 _10499_ ( .A1(_02503_ ), .A2(\ID_EX_imm [15] ), .ZN(_02888_ ) );
NAND2_X1 _10500_ ( .A1(_02526_ ), .A2(\ID_EX_imm [14] ), .ZN(_02889_ ) );
OR2_X1 _10501_ ( .A1(_02504_ ), .A2(_02889_ ), .ZN(_02890_ ) );
NOR2_X1 _10502_ ( .A1(_02504_ ), .A2(_02529_ ), .ZN(_02891_ ) );
NAND2_X1 _10503_ ( .A1(_02552_ ), .A2(\ID_EX_imm [13] ), .ZN(_02892_ ) );
NAND2_X1 _10504_ ( .A1(_02574_ ), .A2(\ID_EX_imm [12] ), .ZN(_02893_ ) );
OAI21_X1 _10505_ ( .A(_02892_ ), .B1(_02553_ ), .B2(_02893_ ), .ZN(_02894_ ) );
NAND2_X1 _10506_ ( .A1(_02891_ ), .A2(_02894_ ), .ZN(_02895_ ) );
NAND4_X1 _10507_ ( .A1(_02887_ ), .A2(_02888_ ), .A3(_02890_ ), .A4(_02895_ ), .ZN(_02896_ ) );
OAI211_X1 _10508_ ( .A(_02385_ ), .B(_02483_ ), .C1(_02878_ ), .C2(_02896_ ), .ZN(_02897_ ) );
AND2_X1 _10509_ ( .A1(_02333_ ), .A2(\ID_EX_imm [22] ), .ZN(_02898_ ) );
NAND2_X1 _10510_ ( .A1(_02309_ ), .A2(_02898_ ), .ZN(_02899_ ) );
INV_X1 _10511_ ( .A(_02307_ ), .ZN(_02900_ ) );
OAI21_X1 _10512_ ( .A(_02899_ ), .B1(_02308_ ), .B2(_02900_ ), .ZN(_02901_ ) );
NAND2_X1 _10513_ ( .A1(_02382_ ), .A2(\ID_EX_imm [20] ), .ZN(_02902_ ) );
NOR3_X1 _10514_ ( .A1(_02902_ ), .A2(_02359_ ), .A3(_02360_ ), .ZN(_02903_ ) );
OR2_X1 _10515_ ( .A1(_02903_ ), .A2(_02360_ ), .ZN(_02904_ ) );
AND2_X1 _10516_ ( .A1(_02480_ ), .A2(\ID_EX_imm [16] ), .ZN(_02905_ ) );
AND2_X1 _10517_ ( .A1(_02459_ ), .A2(_02905_ ), .ZN(_02906_ ) );
AOI21_X1 _10518_ ( .A(_02906_ ), .B1(\ID_EX_imm [17] ), .B2(_02458_ ), .ZN(_02907_ ) );
INV_X1 _10519_ ( .A(_02407_ ), .ZN(_02908_ ) );
OR4_X1 _10520_ ( .A1(_02433_ ), .A2(_02907_ ), .A3(_02432_ ), .A4(_02908_ ), .ZN(_02909_ ) );
AND2_X1 _10521_ ( .A1(_02406_ ), .A2(\ID_EX_imm [18] ), .ZN(_02910_ ) );
AOI21_X1 _10522_ ( .A(_02433_ ), .B1(_02434_ ), .B2(_02910_ ), .ZN(_02911_ ) );
AND2_X1 _10523_ ( .A1(_02909_ ), .A2(_02911_ ), .ZN(_02912_ ) );
INV_X1 _10524_ ( .A(_02912_ ), .ZN(_02913_ ) );
AOI221_X4 _10525_ ( .A(_02901_ ), .B1(_02336_ ), .B2(_02904_ ), .C1(_02913_ ), .C2(_02385_ ), .ZN(_02914_ ) );
AOI21_X1 _10526_ ( .A(_02274_ ), .B1(_02897_ ), .B2(_02914_ ), .ZN(_02915_ ) );
AOI21_X1 _10527_ ( .A(_02272_ ), .B1(_02269_ ), .B2(_02270_ ), .ZN(_02916_ ) );
NOR2_X1 _10528_ ( .A1(_02915_ ), .A2(_02916_ ), .ZN(_02917_ ) );
OR2_X1 _10529_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02918_ ) );
OAI211_X1 _10530_ ( .A(_02918_ ), .B(_02109_ ), .C1(_02120_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02919_ ) );
INV_X1 _10531_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02920_ ) );
NAND2_X1 _10532_ ( .A1(_02920_ ), .A2(fanout_net_22 ), .ZN(_02921_ ) );
OAI211_X1 _10533_ ( .A(_02921_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02922_ ) );
NAND3_X1 _10534_ ( .A1(_02919_ ), .A2(_02922_ ), .A3(_02149_ ), .ZN(_02923_ ) );
MUX2_X1 _10535_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02924_ ) );
MUX2_X1 _10536_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02925_ ) );
MUX2_X1 _10537_ ( .A(_02924_ ), .B(_02925_ ), .S(_02109_ ), .Z(_02926_ ) );
OAI211_X1 _10538_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02923_ ), .C1(_02926_ ), .C2(_02149_ ), .ZN(_02927_ ) );
OR2_X1 _10539_ ( .A1(_02119_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02928_ ) );
OAI211_X1 _10540_ ( .A(_02928_ ), .B(_02109_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02929_ ) );
INV_X1 _10541_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02930_ ) );
NAND2_X1 _10542_ ( .A1(_02930_ ), .A2(fanout_net_22 ), .ZN(_02931_ ) );
OAI211_X1 _10543_ ( .A(_02931_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02932_ ) );
NAND3_X1 _10544_ ( .A1(_02929_ ), .A2(_02932_ ), .A3(_02102_ ), .ZN(_02933_ ) );
MUX2_X1 _10545_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02934_ ) );
MUX2_X1 _10546_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02935_ ) );
MUX2_X1 _10547_ ( .A(_02934_ ), .B(_02935_ ), .S(_02109_ ), .Z(_02936_ ) );
OAI211_X1 _10548_ ( .A(_02098_ ), .B(_02933_ ), .C1(_02936_ ), .C2(_02149_ ), .ZN(_02937_ ) );
OAI211_X1 _10549_ ( .A(_02927_ ), .B(_02937_ ), .C1(_02195_ ), .C2(_02168_ ), .ZN(_02938_ ) );
OR4_X1 _10550_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A2(_02197_ ), .A3(_02167_ ), .A4(_02170_ ), .ZN(_02939_ ) );
NAND2_X1 _10551_ ( .A1(_02938_ ), .A2(_02939_ ), .ZN(_02940_ ) );
NAND2_X1 _10552_ ( .A1(_02940_ ), .A2(\ID_EX_imm [25] ), .ZN(_02941_ ) );
NAND2_X1 _10553_ ( .A1(_02917_ ), .A2(_02941_ ), .ZN(_02942_ ) );
OR2_X1 _10554_ ( .A1(_02120_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02943_ ) );
OAI211_X1 _10555_ ( .A(_02943_ ), .B(_02110_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02944_ ) );
INV_X1 _10556_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02945_ ) );
INV_X1 _10557_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02946_ ) );
MUX2_X1 _10558_ ( .A(_02945_ ), .B(_02946_ ), .S(fanout_net_22 ), .Z(_02947_ ) );
OAI211_X1 _10559_ ( .A(_02944_ ), .B(_02113_ ), .C1(_02947_ ), .C2(_02110_ ), .ZN(_02948_ ) );
MUX2_X1 _10560_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02949_ ) );
MUX2_X1 _10561_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02950_ ) );
MUX2_X1 _10562_ ( .A(_02949_ ), .B(_02950_ ), .S(_02110_ ), .Z(_02951_ ) );
OAI211_X1 _10563_ ( .A(_02948_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .C1(_02951_ ), .C2(_02113_ ), .ZN(_02952_ ) );
OR2_X1 _10564_ ( .A1(_02120_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02953_ ) );
OAI211_X1 _10565_ ( .A(_02953_ ), .B(_02110_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02954_ ) );
OR2_X1 _10566_ ( .A1(_02120_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02955_ ) );
OAI211_X1 _10567_ ( .A(_02955_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02956_ ) );
NAND3_X1 _10568_ ( .A1(_02954_ ), .A2(_02956_ ), .A3(_02113_ ), .ZN(_02957_ ) );
MUX2_X1 _10569_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02958_ ) );
MUX2_X1 _10570_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02959_ ) );
MUX2_X1 _10571_ ( .A(_02958_ ), .B(_02959_ ), .S(_02110_ ), .Z(_02960_ ) );
OAI211_X1 _10572_ ( .A(_02098_ ), .B(_02957_ ), .C1(_02960_ ), .C2(_02113_ ), .ZN(_02961_ ) );
OAI211_X1 _10573_ ( .A(_02952_ ), .B(_02961_ ), .C1(_02195_ ), .C2(_02168_ ), .ZN(_02962_ ) );
OR4_X1 _10574_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A2(_02164_ ), .A3(_02168_ ), .A4(_02170_ ), .ZN(_02963_ ) );
NAND2_X1 _10575_ ( .A1(_02962_ ), .A2(_02963_ ), .ZN(_02964_ ) );
BUF_X4 _10576_ ( .A(_02964_ ), .Z(_02965_ ) );
INV_X1 _10577_ ( .A(\ID_EX_imm [26] ), .ZN(_02966_ ) );
XNOR2_X1 _10578_ ( .A(_02965_ ), .B(_02966_ ), .ZN(_02967_ ) );
INV_X1 _10579_ ( .A(\ID_EX_imm [25] ), .ZN(_02968_ ) );
NAND3_X1 _10580_ ( .A1(_02938_ ), .A2(_02939_ ), .A3(_02968_ ), .ZN(_02969_ ) );
AND4_X1 _10581_ ( .A1(_02250_ ), .A2(_02942_ ), .A3(_02967_ ), .A4(_02969_ ), .ZN(_02970_ ) );
AND2_X1 _10582_ ( .A1(_02965_ ), .A2(\ID_EX_imm [26] ), .ZN(_02971_ ) );
AND2_X1 _10583_ ( .A1(_02250_ ), .A2(_02971_ ), .ZN(_02972_ ) );
AOI21_X1 _10584_ ( .A(_02972_ ), .B1(\ID_EX_imm [27] ), .B2(_02248_ ), .ZN(_02973_ ) );
INV_X1 _10585_ ( .A(_02973_ ), .ZN(_02974_ ) );
OAI211_X1 _10586_ ( .A(_02201_ ), .B(_02228_ ), .C1(_02970_ ), .C2(_02974_ ), .ZN(_02975_ ) );
INV_X1 _10587_ ( .A(_02225_ ), .ZN(_02976_ ) );
NOR2_X1 _10588_ ( .A1(_02976_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02977_ ) );
INV_X1 _10589_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02978_ ) );
AOI22_X1 _10590_ ( .A1(_02977_ ), .A2(_02201_ ), .B1(_02978_ ), .B2(_02199_ ), .ZN(_02979_ ) );
AOI21_X1 _10591_ ( .A(_02174_ ), .B1(_02975_ ), .B2(_02979_ ), .ZN(_02980_ ) );
AOI21_X1 _10592_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02160_ ), .B2(_02171_ ), .ZN(_02981_ ) );
NOR2_X1 _10593_ ( .A1(_02980_ ), .A2(_02981_ ), .ZN(_02982_ ) );
OR2_X1 _10594_ ( .A1(_02120_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02983_ ) );
OAI211_X1 _10595_ ( .A(_02983_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02984_ ) );
OR2_X1 _10596_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02985_ ) );
OAI211_X1 _10597_ ( .A(_02985_ ), .B(_02125_ ), .C1(_02121_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02986_ ) );
NAND3_X1 _10598_ ( .A1(_02984_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02986_ ), .ZN(_02987_ ) );
MUX2_X1 _10599_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02988_ ) );
MUX2_X1 _10600_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02989_ ) );
MUX2_X1 _10601_ ( .A(_02988_ ), .B(_02989_ ), .S(_02125_ ), .Z(_02990_ ) );
OAI211_X1 _10602_ ( .A(_02098_ ), .B(_02987_ ), .C1(_02990_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02991_ ) );
NOR2_X1 _10603_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02992_ ) );
OAI21_X1 _10604_ ( .A(_02109_ ), .B1(_02121_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02993_ ) );
INV_X1 _10605_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02994_ ) );
INV_X1 _10606_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02995_ ) );
MUX2_X1 _10607_ ( .A(_02994_ ), .B(_02995_ ), .S(fanout_net_22 ), .Z(_02996_ ) );
OAI221_X1 _10608_ ( .A(_02149_ ), .B1(_02992_ ), .B2(_02993_ ), .C1(_02996_ ), .C2(_02110_ ), .ZN(_02997_ ) );
MUX2_X1 _10609_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02998_ ) );
MUX2_X1 _10610_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02999_ ) );
MUX2_X1 _10611_ ( .A(_02998_ ), .B(_02999_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03000_ ) );
OAI211_X1 _10612_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02997_ ), .C1(_03000_ ), .C2(_02113_ ), .ZN(_03001_ ) );
OAI211_X1 _10613_ ( .A(_02991_ ), .B(_03001_ ), .C1(_02195_ ), .C2(_02168_ ), .ZN(_03002_ ) );
OR4_X1 _10614_ ( .A1(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A2(_02197_ ), .A3(_02167_ ), .A4(_02170_ ), .ZN(_03003_ ) );
NAND2_X1 _10615_ ( .A1(_03002_ ), .A2(_03003_ ), .ZN(_03004_ ) );
BUF_X2 _10616_ ( .A(_03004_ ), .Z(_03005_ ) );
XNOR2_X1 _10617_ ( .A(_03005_ ), .B(\ID_EX_imm [31] ), .ZN(_03006_ ) );
XNOR2_X1 _10618_ ( .A(_02982_ ), .B(_03006_ ), .ZN(_03007_ ) );
AND2_X2 _10619_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_03008_ ) );
BUF_X4 _10620_ ( .A(_03008_ ), .Z(_03009_ ) );
NOR2_X1 _10621_ ( .A1(_03007_ ), .A2(_03009_ ), .ZN(_00097_ ) );
AND3_X1 _10622_ ( .A1(_02975_ ), .A2(_02979_ ), .A3(_02174_ ), .ZN(_03010_ ) );
NOR3_X1 _10623_ ( .A1(_03010_ ), .A2(_02980_ ), .A3(_03008_ ), .ZN(_00098_ ) );
OAI21_X1 _10624_ ( .A(_02483_ ), .B1(_02878_ ), .B2(_02896_ ), .ZN(_03011_ ) );
AND2_X1 _10625_ ( .A1(_03011_ ), .A2(_02912_ ), .ZN(_03012_ ) );
INV_X1 _10626_ ( .A(_02384_ ), .ZN(_03013_ ) );
OR2_X1 _10627_ ( .A1(_03012_ ), .A2(_03013_ ), .ZN(_03014_ ) );
NAND2_X1 _10628_ ( .A1(_03014_ ), .A2(_02902_ ), .ZN(_03015_ ) );
XNOR2_X1 _10629_ ( .A(_03015_ ), .B(_02361_ ), .ZN(_03016_ ) );
NOR2_X1 _10630_ ( .A1(_03016_ ), .A2(_03009_ ), .ZN(_00099_ ) );
XNOR2_X1 _10631_ ( .A(_03012_ ), .B(_02384_ ), .ZN(_03017_ ) );
INV_X1 _10632_ ( .A(_03008_ ), .ZN(_03018_ ) );
CLKBUF_X2 _10633_ ( .A(_03018_ ), .Z(_03019_ ) );
AND2_X1 _10634_ ( .A1(_03017_ ), .A2(_03019_ ), .ZN(_00100_ ) );
NOR2_X1 _10635_ ( .A1(_02878_ ), .A2(_02896_ ), .ZN(_03020_ ) );
NAND2_X1 _10636_ ( .A1(_02459_ ), .A2(_02482_ ), .ZN(_03021_ ) );
OR2_X1 _10637_ ( .A1(_03020_ ), .A2(_03021_ ), .ZN(_03022_ ) );
AOI21_X1 _10638_ ( .A(_02908_ ), .B1(_03022_ ), .B2(_02907_ ), .ZN(_03023_ ) );
OR2_X1 _10639_ ( .A1(_03023_ ), .A2(_02910_ ), .ZN(_03024_ ) );
XNOR2_X1 _10640_ ( .A(_03024_ ), .B(_02434_ ), .ZN(_03025_ ) );
NOR2_X1 _10641_ ( .A1(_03025_ ), .A2(_03009_ ), .ZN(_00101_ ) );
AND3_X1 _10642_ ( .A1(_03022_ ), .A2(_02908_ ), .A3(_02907_ ), .ZN(_03026_ ) );
NOR3_X1 _10643_ ( .A1(_03026_ ), .A2(_03023_ ), .A3(_03008_ ), .ZN(_00102_ ) );
AND3_X1 _10644_ ( .A1(_02478_ ), .A2(_02481_ ), .A3(_02479_ ), .ZN(_03027_ ) );
NOR3_X1 _10645_ ( .A1(_03020_ ), .A2(_02905_ ), .A3(_03027_ ), .ZN(_03028_ ) );
OR2_X1 _10646_ ( .A1(_03028_ ), .A2(_02905_ ), .ZN(_03029_ ) );
XNOR2_X1 _10647_ ( .A(_03029_ ), .B(_02459_ ), .ZN(_03030_ ) );
NOR2_X1 _10648_ ( .A1(_03030_ ), .A2(_03009_ ), .ZN(_00103_ ) );
XNOR2_X1 _10649_ ( .A(_03020_ ), .B(_02482_ ), .ZN(_03031_ ) );
AND2_X1 _10650_ ( .A1(_03031_ ), .A2(_03019_ ), .ZN(_00104_ ) );
AOI21_X1 _10651_ ( .A(_02674_ ), .B1(_02869_ ), .B2(_02877_ ), .ZN(_03032_ ) );
INV_X1 _10652_ ( .A(_02886_ ), .ZN(_03033_ ) );
NOR2_X1 _10653_ ( .A1(_03032_ ), .A2(_03033_ ), .ZN(_03034_ ) );
NOR3_X1 _10654_ ( .A1(_03034_ ), .A2(_02553_ ), .A3(_02577_ ), .ZN(_03035_ ) );
OAI21_X1 _10655_ ( .A(_02528_ ), .B1(_03035_ ), .B2(_02894_ ), .ZN(_03036_ ) );
AND2_X1 _10656_ ( .A1(_03036_ ), .A2(_02889_ ), .ZN(_03037_ ) );
XNOR2_X1 _10657_ ( .A(_03037_ ), .B(_02504_ ), .ZN(_03038_ ) );
NOR2_X1 _10658_ ( .A1(_03038_ ), .A2(_03009_ ), .ZN(_00105_ ) );
OR3_X1 _10659_ ( .A1(_03035_ ), .A2(_02528_ ), .A3(_02894_ ), .ZN(_03039_ ) );
AND3_X1 _10660_ ( .A1(_03039_ ), .A2(_03019_ ), .A3(_03036_ ), .ZN(_00106_ ) );
OAI21_X1 _10661_ ( .A(_02576_ ), .B1(_03032_ ), .B2(_03033_ ), .ZN(_03040_ ) );
AND2_X1 _10662_ ( .A1(_03040_ ), .A2(_02893_ ), .ZN(_03041_ ) );
XNOR2_X1 _10663_ ( .A(_03041_ ), .B(_02553_ ), .ZN(_03042_ ) );
NOR2_X1 _10664_ ( .A1(_03042_ ), .A2(_03009_ ), .ZN(_00107_ ) );
XNOR2_X1 _10665_ ( .A(_03034_ ), .B(_02576_ ), .ZN(_03043_ ) );
AND2_X1 _10666_ ( .A1(_03043_ ), .A2(_03019_ ), .ZN(_00108_ ) );
NOR2_X1 _10667_ ( .A1(_02970_ ), .A2(_02974_ ), .ZN(_03044_ ) );
NOR2_X1 _10668_ ( .A1(_03044_ ), .A2(_02227_ ), .ZN(_03045_ ) );
OR2_X1 _10669_ ( .A1(_03045_ ), .A2(_02977_ ), .ZN(_03046_ ) );
XNOR2_X1 _10670_ ( .A(_03046_ ), .B(_02201_ ), .ZN(_03047_ ) );
NOR2_X1 _10671_ ( .A1(_03047_ ), .A2(_03009_ ), .ZN(_00109_ ) );
XNOR2_X1 _10672_ ( .A(_03044_ ), .B(_02228_ ), .ZN(_03048_ ) );
AND2_X1 _10673_ ( .A1(_03048_ ), .A2(_03019_ ), .ZN(_00110_ ) );
AND3_X1 _10674_ ( .A1(_02942_ ), .A2(_02967_ ), .A3(_02969_ ), .ZN(_03049_ ) );
OR2_X1 _10675_ ( .A1(_03049_ ), .A2(_02971_ ), .ZN(_03050_ ) );
XNOR2_X1 _10676_ ( .A(_03050_ ), .B(_02250_ ), .ZN(_03051_ ) );
NOR2_X1 _10677_ ( .A1(_03051_ ), .A2(_03009_ ), .ZN(_00111_ ) );
AOI21_X1 _10678_ ( .A(_02967_ ), .B1(_02942_ ), .B2(_02969_ ), .ZN(_03052_ ) );
NOR3_X1 _10679_ ( .A1(_03049_ ), .A2(_03052_ ), .A3(_03008_ ), .ZN(_00112_ ) );
NAND2_X1 _10680_ ( .A1(_02941_ ), .A2(_02969_ ), .ZN(_03053_ ) );
XNOR2_X1 _10681_ ( .A(_02917_ ), .B(_03053_ ), .ZN(_03054_ ) );
NOR2_X1 _10682_ ( .A1(_03054_ ), .A2(_03009_ ), .ZN(_00113_ ) );
AND3_X1 _10683_ ( .A1(_02897_ ), .A2(_02914_ ), .A3(_02274_ ), .ZN(_03055_ ) );
NOR3_X1 _10684_ ( .A1(_03055_ ), .A2(_02915_ ), .A3(_03008_ ), .ZN(_00114_ ) );
NOR4_X1 _10685_ ( .A1(_03012_ ), .A2(_02359_ ), .A3(_02360_ ), .A4(_03013_ ), .ZN(_03056_ ) );
OR2_X1 _10686_ ( .A1(_03056_ ), .A2(_02904_ ), .ZN(_03057_ ) );
AND2_X1 _10687_ ( .A1(_03057_ ), .A2(_02335_ ), .ZN(_03058_ ) );
OR2_X1 _10688_ ( .A1(_03058_ ), .A2(_02898_ ), .ZN(_03059_ ) );
XNOR2_X1 _10689_ ( .A(_03059_ ), .B(_02309_ ), .ZN(_03060_ ) );
NOR2_X1 _10690_ ( .A1(_03060_ ), .A2(_03009_ ), .ZN(_00115_ ) );
XOR2_X1 _10691_ ( .A(_03057_ ), .B(_02335_ ), .Z(_03061_ ) );
AND2_X1 _10692_ ( .A1(_03061_ ), .A2(_03019_ ), .ZN(_00116_ ) );
INV_X1 _10693_ ( .A(\IF_ID_inst [6] ), .ZN(_03062_ ) );
NOR2_X1 _10694_ ( .A1(_03062_ ), .A2(\IF_ID_inst [12] ), .ZN(_03063_ ) );
AND2_X2 _10695_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03064_ ) );
AND3_X1 _10696_ ( .A1(_03063_ ), .A2(\IF_ID_inst [13] ), .A3(_03064_ ), .ZN(_03065_ ) );
AND2_X1 _10697_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_03066_ ) );
NOR2_X1 _10698_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_03067_ ) );
AND2_X1 _10699_ ( .A1(_03066_ ), .A2(_03067_ ), .ZN(_03068_ ) );
CLKBUF_X2 _10700_ ( .A(_03068_ ), .Z(_03069_ ) );
CLKBUF_X2 _10701_ ( .A(_03069_ ), .Z(_03070_ ) );
AND2_X1 _10702_ ( .A1(_03065_ ), .A2(_03070_ ), .ZN(_03071_ ) );
AND4_X1 _10703_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03072_ ) );
AND2_X1 _10704_ ( .A1(_03070_ ), .A2(_03072_ ), .ZN(_03073_ ) );
NOR2_X1 _10705_ ( .A1(_03071_ ), .A2(_03073_ ), .ZN(_03074_ ) );
BUF_X4 _10706_ ( .A(_03074_ ), .Z(_03075_ ) );
INV_X1 _10707_ ( .A(\IF_ID_inst [31] ), .ZN(_03076_ ) );
AND2_X1 _10708_ ( .A1(_02093_ ), .A2(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03077_ ) );
INV_X1 _10709_ ( .A(_03077_ ), .ZN(_03078_ ) );
BUF_X4 _10710_ ( .A(_03078_ ), .Z(_03079_ ) );
NOR3_X1 _10711_ ( .A1(_03075_ ), .A2(_03076_ ), .A3(_03079_ ), .ZN(_00195_ ) );
INV_X1 _10712_ ( .A(\IF_ID_inst [30] ), .ZN(_03080_ ) );
NOR3_X1 _10713_ ( .A1(_03075_ ), .A2(_03080_ ), .A3(_03079_ ), .ZN(_00196_ ) );
INV_X1 _10714_ ( .A(\IF_ID_inst [21] ), .ZN(_03081_ ) );
NOR3_X1 _10715_ ( .A1(_03075_ ), .A2(_03081_ ), .A3(_03079_ ), .ZN(_00197_ ) );
BUF_X4 _10716_ ( .A(_03078_ ), .Z(_03082_ ) );
INV_X1 _10717_ ( .A(_03074_ ), .ZN(_03083_ ) );
INV_X1 _10718_ ( .A(\IF_ID_inst [20] ), .ZN(_03084_ ) );
AOI21_X1 _10719_ ( .A(_03082_ ), .B1(_03083_ ), .B2(_03084_ ), .ZN(_00198_ ) );
INV_X1 _10720_ ( .A(\IF_ID_inst [29] ), .ZN(_03085_ ) );
AOI21_X1 _10721_ ( .A(_03082_ ), .B1(_03083_ ), .B2(_03085_ ), .ZN(_00199_ ) );
INV_X1 _10722_ ( .A(\IF_ID_inst [28] ), .ZN(_03086_ ) );
AOI21_X1 _10723_ ( .A(_03082_ ), .B1(_03083_ ), .B2(_03086_ ), .ZN(_00200_ ) );
INV_X1 _10724_ ( .A(\IF_ID_inst [27] ), .ZN(_03087_ ) );
NOR3_X1 _10725_ ( .A1(_03075_ ), .A2(_03087_ ), .A3(_03079_ ), .ZN(_00201_ ) );
INV_X1 _10726_ ( .A(\IF_ID_inst [26] ), .ZN(_03088_ ) );
AOI21_X1 _10727_ ( .A(_03082_ ), .B1(_03083_ ), .B2(_03088_ ), .ZN(_00202_ ) );
INV_X1 _10728_ ( .A(\IF_ID_inst [25] ), .ZN(_03089_ ) );
NOR3_X1 _10729_ ( .A1(_03075_ ), .A2(_03089_ ), .A3(_03079_ ), .ZN(_00203_ ) );
INV_X1 _10730_ ( .A(\IF_ID_inst [24] ), .ZN(_03090_ ) );
BUF_X4 _10731_ ( .A(_03078_ ), .Z(_03091_ ) );
NOR3_X1 _10732_ ( .A1(_03075_ ), .A2(_03090_ ), .A3(_03091_ ), .ZN(_00204_ ) );
INV_X1 _10733_ ( .A(\IF_ID_inst [23] ), .ZN(_03092_ ) );
NOR3_X1 _10734_ ( .A1(_03075_ ), .A2(_03092_ ), .A3(_03091_ ), .ZN(_00205_ ) );
INV_X1 _10735_ ( .A(\IF_ID_inst [22] ), .ZN(_03093_ ) );
NOR3_X1 _10736_ ( .A1(_03075_ ), .A2(_03093_ ), .A3(_03091_ ), .ZN(_00206_ ) );
AND4_X1 _10737_ ( .A1(_01535_ ), .A2(_02092_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .A4(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00207_ ) );
AND4_X1 _10738_ ( .A1(_01535_ ), .A2(_02092_ ), .A3(\myidu.state [2] ), .A4(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00208_ ) );
AND3_X1 _10739_ ( .A1(_03069_ ), .A2(\IF_ID_inst [12] ), .A3(\IF_ID_inst [6] ), .ZN(_03094_ ) );
INV_X1 _10740_ ( .A(\IF_ID_inst [5] ), .ZN(_03095_ ) );
NOR2_X1 _10741_ ( .A1(_03095_ ), .A2(\IF_ID_inst [4] ), .ZN(_03096_ ) );
AND2_X2 _10742_ ( .A1(_03094_ ), .A2(_03096_ ), .ZN(_03097_ ) );
AND2_X2 _10743_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03098_ ) );
NAND2_X1 _10744_ ( .A1(_03097_ ), .A2(_03098_ ), .ZN(_03099_ ) );
INV_X1 _10745_ ( .A(\IF_ID_inst [7] ), .ZN(_03100_ ) );
AND4_X1 _10746_ ( .A1(\IF_ID_inst [6] ), .A2(_03070_ ), .A3(_03100_ ), .A4(_03064_ ), .ZN(_03101_ ) );
OR3_X1 _10747_ ( .A1(\IF_ID_inst [11] ), .A2(\IF_ID_inst [10] ), .A3(\IF_ID_inst [9] ), .ZN(_03102_ ) );
NOR2_X1 _10748_ ( .A1(_03102_ ), .A2(\IF_ID_inst [8] ), .ZN(_03103_ ) );
NOR4_X1 _10749_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_03104_ ) );
AND3_X1 _10750_ ( .A1(_03101_ ), .A2(_03103_ ), .A3(_03104_ ), .ZN(_03105_ ) );
NOR2_X1 _10751_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_03106_ ) );
AND3_X1 _10752_ ( .A1(_03106_ ), .A2(\IF_ID_inst [21] ), .A3(_03084_ ), .ZN(_03107_ ) );
NOR2_X1 _10753_ ( .A1(\IF_ID_inst [18] ), .A2(\IF_ID_inst [17] ), .ZN(_03108_ ) );
NOR2_X1 _10754_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [16] ), .ZN(_03109_ ) );
AND2_X1 _10755_ ( .A1(_03108_ ), .A2(_03109_ ), .ZN(_03110_ ) );
AND2_X1 _10756_ ( .A1(_03107_ ), .A2(_03110_ ), .ZN(_03111_ ) );
NOR3_X1 _10757_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .A3(\IF_ID_inst [24] ), .ZN(_03112_ ) );
NAND2_X1 _10758_ ( .A1(_03080_ ), .A2(\IF_ID_inst [29] ), .ZN(_03113_ ) );
NOR3_X1 _10759_ ( .A1(_03113_ ), .A2(_03086_ ), .A3(\IF_ID_inst [31] ), .ZN(_03114_ ) );
AND4_X1 _10760_ ( .A1(_03087_ ), .A2(_03111_ ), .A3(_03112_ ), .A4(_03114_ ), .ZN(_03115_ ) );
NAND2_X1 _10761_ ( .A1(_03105_ ), .A2(_03115_ ), .ZN(_03116_ ) );
NAND4_X1 _10762_ ( .A1(_03110_ ), .A2(_03081_ ), .A3(\IF_ID_inst [20] ), .A4(_03106_ ), .ZN(_03117_ ) );
NAND2_X1 _10763_ ( .A1(_03112_ ), .A2(_03087_ ), .ZN(_03118_ ) );
NAND4_X1 _10764_ ( .A1(_03080_ ), .A2(_03085_ ), .A3(_03086_ ), .A4(_03076_ ), .ZN(_03119_ ) );
NOR3_X1 _10765_ ( .A1(_03117_ ), .A2(_03118_ ), .A3(_03119_ ), .ZN(_03120_ ) );
NAND2_X1 _10766_ ( .A1(_03105_ ), .A2(_03120_ ), .ZN(_03121_ ) );
AND3_X1 _10767_ ( .A1(_03066_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_03122_ ) );
CLKBUF_X2 _10768_ ( .A(_03122_ ), .Z(_03123_ ) );
NOR2_X1 _10769_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03124_ ) );
AND3_X1 _10770_ ( .A1(_03124_ ), .A2(\IF_ID_inst [12] ), .A3(_03062_ ), .ZN(_03125_ ) );
AND2_X1 _10771_ ( .A1(_03123_ ), .A2(_03125_ ), .ZN(_03126_ ) );
NOR2_X1 _10772_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03127_ ) );
BUF_X2 _10773_ ( .A(_03127_ ), .Z(_03128_ ) );
NAND2_X1 _10774_ ( .A1(_03126_ ), .A2(_03128_ ), .ZN(_03129_ ) );
AND4_X1 _10775_ ( .A1(_03099_ ), .A2(_03116_ ), .A3(_03121_ ), .A4(_03129_ ), .ZN(_03130_ ) );
INV_X1 _10776_ ( .A(\IF_ID_inst [14] ), .ZN(_03131_ ) );
NOR2_X1 _10777_ ( .A1(_03131_ ), .A2(\IF_ID_inst [13] ), .ZN(_03132_ ) );
AND2_X1 _10778_ ( .A1(_03063_ ), .A2(_03096_ ), .ZN(_03133_ ) );
AND2_X2 _10779_ ( .A1(_03133_ ), .A2(_03070_ ), .ZN(_03134_ ) );
AOI22_X1 _10780_ ( .A1(_03097_ ), .A2(_03132_ ), .B1(_03098_ ), .B2(_03134_ ), .ZN(_03135_ ) );
AOI22_X1 _10781_ ( .A1(_03097_ ), .A2(_03128_ ), .B1(_03132_ ), .B2(_03134_ ), .ZN(_03136_ ) );
NOR2_X1 _10782_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03137_ ) );
AND3_X1 _10783_ ( .A1(_03070_ ), .A2(_03096_ ), .A3(_03137_ ), .ZN(_03138_ ) );
INV_X1 _10784_ ( .A(\IF_ID_inst [13] ), .ZN(_03139_ ) );
NOR2_X1 _10785_ ( .A1(_03139_ ), .A2(\IF_ID_inst [14] ), .ZN(_03140_ ) );
AOI22_X1 _10786_ ( .A1(_03128_ ), .A2(_03134_ ), .B1(_03138_ ), .B2(_03140_ ), .ZN(_03141_ ) );
INV_X1 _10787_ ( .A(\IF_ID_inst [12] ), .ZN(_03142_ ) );
NOR2_X1 _10788_ ( .A1(_03142_ ), .A2(\IF_ID_inst [6] ), .ZN(_03143_ ) );
AND3_X1 _10789_ ( .A1(_03070_ ), .A2(_03096_ ), .A3(_03143_ ), .ZN(_03144_ ) );
NAND2_X1 _10790_ ( .A1(_03144_ ), .A2(_03128_ ), .ZN(_03145_ ) );
NAND2_X1 _10791_ ( .A1(_03138_ ), .A2(_03128_ ), .ZN(_03146_ ) );
AND2_X1 _10792_ ( .A1(_03145_ ), .A2(_03146_ ), .ZN(_03147_ ) );
AND4_X1 _10793_ ( .A1(_03135_ ), .A2(_03136_ ), .A3(_03141_ ), .A4(_03147_ ), .ZN(_03148_ ) );
CLKBUF_X2 _10794_ ( .A(_03077_ ), .Z(_03149_ ) );
AND4_X1 _10795_ ( .A1(\IF_ID_inst [11] ), .A2(_03130_ ), .A3(_03148_ ), .A4(_03149_ ), .ZN(_00209_ ) );
AND4_X1 _10796_ ( .A1(\IF_ID_inst [10] ), .A2(_03130_ ), .A3(_03148_ ), .A4(_03149_ ), .ZN(_00210_ ) );
AND4_X1 _10797_ ( .A1(\IF_ID_inst [9] ), .A2(_03130_ ), .A3(_03148_ ), .A4(_03149_ ), .ZN(_00211_ ) );
AND4_X1 _10798_ ( .A1(\IF_ID_inst [8] ), .A2(_03130_ ), .A3(_03148_ ), .A4(_03149_ ), .ZN(_00212_ ) );
AND4_X1 _10799_ ( .A1(\IF_ID_inst [7] ), .A2(_03130_ ), .A3(_03148_ ), .A4(_03149_ ), .ZN(_00213_ ) );
AND2_X1 _10800_ ( .A1(_03121_ ), .A2(_03129_ ), .ZN(_03150_ ) );
BUF_X2 _10801_ ( .A(_03149_ ), .Z(_03151_ ) );
NOR2_X1 _10802_ ( .A1(\IF_ID_inst [7] ), .A2(\IF_ID_inst [15] ), .ZN(_03152_ ) );
AND4_X1 _10803_ ( .A1(_03064_ ), .A2(_03063_ ), .A3(_03127_ ), .A4(_03152_ ), .ZN(_03153_ ) );
AND3_X1 _10804_ ( .A1(_03153_ ), .A2(_03070_ ), .A3(_03103_ ), .ZN(_03154_ ) );
NAND3_X1 _10805_ ( .A1(_03114_ ), .A2(_03107_ ), .A3(_03110_ ), .ZN(_03155_ ) );
NOR2_X1 _10806_ ( .A1(_03155_ ), .A2(_03118_ ), .ZN(_03156_ ) );
AND2_X1 _10807_ ( .A1(_03154_ ), .A2(_03156_ ), .ZN(_03157_ ) );
INV_X1 _10808_ ( .A(_03096_ ), .ZN(_03158_ ) );
NOR2_X1 _10809_ ( .A1(_03158_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03159_ ) );
AND2_X2 _10810_ ( .A1(_03159_ ), .A2(_03122_ ), .ZN(_03160_ ) );
BUF_X2 _10811_ ( .A(_03160_ ), .Z(_03161_ ) );
NAND3_X1 _10812_ ( .A1(\IF_ID_inst [2] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [1] ), .ZN(_03162_ ) );
NOR2_X1 _10813_ ( .A1(_03162_ ), .A2(\IF_ID_inst [3] ), .ZN(_03163_ ) );
INV_X1 _10814_ ( .A(\IF_ID_inst [4] ), .ZN(_03164_ ) );
NOR2_X1 _10815_ ( .A1(_03164_ ), .A2(\IF_ID_inst [6] ), .ZN(_03165_ ) );
AND2_X2 _10816_ ( .A1(_03163_ ), .A2(_03165_ ), .ZN(_03166_ ) );
NOR3_X1 _10817_ ( .A1(_03157_ ), .A2(_03161_ ), .A3(_03166_ ), .ZN(_03167_ ) );
AND4_X1 _10818_ ( .A1(\IF_ID_inst [19] ), .A2(_03150_ ), .A3(_03151_ ), .A4(_03167_ ), .ZN(_00214_ ) );
AND4_X1 _10819_ ( .A1(\IF_ID_inst [18] ), .A2(_03150_ ), .A3(_03151_ ), .A4(_03167_ ), .ZN(_00215_ ) );
AND4_X1 _10820_ ( .A1(\IF_ID_inst [17] ), .A2(_03150_ ), .A3(_03149_ ), .A4(_03167_ ), .ZN(_00216_ ) );
XNOR2_X1 _10821_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_03168_ ) );
XNOR2_X1 _10822_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_03169_ ) );
XNOR2_X1 _10823_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_03170_ ) );
XNOR2_X1 _10824_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_03171_ ) );
AND4_X1 _10825_ ( .A1(_03168_ ), .A2(_03169_ ), .A3(_03170_ ), .A4(_03171_ ), .ZN(_03172_ ) );
XNOR2_X1 _10826_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_03173_ ) );
XNOR2_X1 _10827_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_03174_ ) );
XNOR2_X1 _10828_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_03175_ ) );
XNOR2_X1 _10829_ ( .A(\IF_ID_pc [21] ), .B(\myexu.pc_jump [21] ), .ZN(_03176_ ) );
NAND4_X1 _10830_ ( .A1(_03173_ ), .A2(_03174_ ), .A3(_03175_ ), .A4(_03176_ ), .ZN(_03177_ ) );
XNOR2_X1 _10831_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_03178_ ) );
XNOR2_X1 _10832_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_03179_ ) );
XNOR2_X1 _10833_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_03180_ ) );
XNOR2_X1 _10834_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_03181_ ) );
NAND4_X1 _10835_ ( .A1(_03178_ ), .A2(_03179_ ), .A3(_03180_ ), .A4(_03181_ ), .ZN(_03182_ ) );
XNOR2_X1 _10836_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_03183_ ) );
XNOR2_X1 _10837_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_03184_ ) );
XNOR2_X1 _10838_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_03185_ ) );
XNOR2_X1 _10839_ ( .A(fanout_net_10 ), .B(\myexu.pc_jump [4] ), .ZN(_03186_ ) );
NAND4_X1 _10840_ ( .A1(_03183_ ), .A2(_03184_ ), .A3(_03185_ ), .A4(_03186_ ), .ZN(_03187_ ) );
XNOR2_X1 _10841_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_03188_ ) );
XNOR2_X1 _10842_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_03189_ ) );
XNOR2_X1 _10843_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_03190_ ) );
XNOR2_X1 _10844_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_03191_ ) );
NAND4_X1 _10845_ ( .A1(_03188_ ), .A2(_03189_ ), .A3(_03190_ ), .A4(_03191_ ), .ZN(_03192_ ) );
NOR4_X1 _10846_ ( .A1(_03177_ ), .A2(_03182_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03193_ ) );
XNOR2_X1 _10847_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_03194_ ) );
XNOR2_X1 _10848_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_03195_ ) );
XNOR2_X1 _10849_ ( .A(fanout_net_6 ), .B(\myexu.pc_jump [3] ), .ZN(_03196_ ) );
XNOR2_X1 _10850_ ( .A(\myexu.pc_jump [2] ), .B(\IF_ID_pc [2] ), .ZN(_03197_ ) );
AND4_X1 _10851_ ( .A1(_03194_ ), .A2(_03195_ ), .A3(_03196_ ), .A4(_03197_ ), .ZN(_03198_ ) );
XNOR2_X1 _10852_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_03199_ ) );
XNOR2_X1 _10853_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_03200_ ) );
XNOR2_X1 _10854_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_03201_ ) );
XNOR2_X1 _10855_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_03202_ ) );
NAND4_X1 _10856_ ( .A1(_03199_ ), .A2(_03200_ ), .A3(_03201_ ), .A4(_03202_ ), .ZN(_03203_ ) );
XNOR2_X1 _10857_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_03204_ ) );
XNOR2_X1 _10858_ ( .A(\IF_ID_pc [25] ), .B(\myexu.pc_jump [25] ), .ZN(_03205_ ) );
NAND2_X1 _10859_ ( .A1(_03204_ ), .A2(_03205_ ), .ZN(_03206_ ) );
XOR2_X1 _10860_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .Z(_03207_ ) );
XOR2_X1 _10861_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .Z(_03208_ ) );
NOR4_X1 _10862_ ( .A1(_03203_ ), .A2(_03206_ ), .A3(_03207_ ), .A4(_03208_ ), .ZN(_03209_ ) );
AND4_X2 _10863_ ( .A1(_03172_ ), .A2(_03193_ ), .A3(_03198_ ), .A4(_03209_ ), .ZN(_03210_ ) );
INV_X1 _10864_ ( .A(check_quest ), .ZN(_03211_ ) );
NOR2_X2 _10865_ ( .A1(_03210_ ), .A2(_03211_ ), .ZN(_03212_ ) );
INV_X1 _10866_ ( .A(\myifu.state [1] ), .ZN(_03213_ ) );
NOR2_X1 _10867_ ( .A1(_03213_ ), .A2(\myifu.to_reset ), .ZN(_03214_ ) );
INV_X1 _10868_ ( .A(_03214_ ), .ZN(_03215_ ) );
NOR2_X1 _10869_ ( .A1(_03212_ ), .A2(_03215_ ), .ZN(_03216_ ) );
AND2_X1 _10870_ ( .A1(_03216_ ), .A2(IDU_ready_IFU ), .ZN(_03217_ ) );
INV_X1 _10871_ ( .A(_03217_ ), .ZN(_03218_ ) );
BUF_X4 _10872_ ( .A(_03218_ ), .Z(_03219_ ) );
OAI21_X1 _10873_ ( .A(\IF_ID_inst [14] ), .B1(_03097_ ), .B2(_03134_ ), .ZN(_03220_ ) );
AND3_X1 _10874_ ( .A1(_03133_ ), .A2(_03069_ ), .A3(_03127_ ), .ZN(_03221_ ) );
AOI21_X1 _10875_ ( .A(_03221_ ), .B1(_03097_ ), .B2(_03127_ ), .ZN(_03222_ ) );
AND2_X1 _10876_ ( .A1(_03220_ ), .A2(_03222_ ), .ZN(_03223_ ) );
AND3_X1 _10877_ ( .A1(_03096_ ), .A2(_03143_ ), .A3(_03127_ ), .ZN(_03224_ ) );
AND3_X1 _10878_ ( .A1(_03224_ ), .A2(_03066_ ), .A3(_03067_ ), .ZN(_03225_ ) );
AND3_X1 _10879_ ( .A1(_03069_ ), .A2(_03096_ ), .A3(_03137_ ), .ZN(_03226_ ) );
AOI21_X1 _10880_ ( .A(_03225_ ), .B1(_03226_ ), .B2(_03127_ ), .ZN(_03227_ ) );
AND2_X1 _10881_ ( .A1(_03226_ ), .A2(_03140_ ), .ZN(_03228_ ) );
INV_X1 _10882_ ( .A(_03228_ ), .ZN(_03229_ ) );
AND2_X1 _10883_ ( .A1(_03227_ ), .A2(_03229_ ), .ZN(_03230_ ) );
AND2_X1 _10884_ ( .A1(_03223_ ), .A2(_03230_ ), .ZN(_03231_ ) );
INV_X1 _10885_ ( .A(_03231_ ), .ZN(_03232_ ) );
AND2_X2 _10886_ ( .A1(_03069_ ), .A2(_03137_ ), .ZN(_03233_ ) );
NOR3_X1 _10887_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_03234_ ) );
AND3_X1 _10888_ ( .A1(_03234_ ), .A2(_03087_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03235_ ) );
NOR2_X1 _10889_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_03236_ ) );
AND2_X1 _10890_ ( .A1(_03132_ ), .A2(_03236_ ), .ZN(_03237_ ) );
AND2_X1 _10891_ ( .A1(_03235_ ), .A2(_03237_ ), .ZN(_03238_ ) );
AND2_X1 _10892_ ( .A1(_03127_ ), .A2(_03236_ ), .ZN(_03239_ ) );
AND2_X1 _10893_ ( .A1(_03235_ ), .A2(_03239_ ), .ZN(_03240_ ) );
OAI211_X1 _10894_ ( .A(_03064_ ), .B(_03233_ ), .C1(_03238_ ), .C2(_03240_ ), .ZN(_03241_ ) );
AND2_X1 _10895_ ( .A1(_03234_ ), .A2(_03087_ ), .ZN(_03242_ ) );
AND4_X1 _10896_ ( .A1(_03131_ ), .A2(_03236_ ), .A3(\IF_ID_inst [13] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03243_ ) );
AND2_X1 _10897_ ( .A1(_03242_ ), .A2(_03243_ ), .ZN(_03244_ ) );
NOR3_X1 _10898_ ( .A1(_03238_ ), .A2(_03240_ ), .A3(_03244_ ), .ZN(_03245_ ) );
AND4_X1 _10899_ ( .A1(\IF_ID_inst [4] ), .A2(_03062_ ), .A3(\IF_ID_inst [5] ), .A4(\IF_ID_inst [12] ), .ZN(_03246_ ) );
AND2_X1 _10900_ ( .A1(_03069_ ), .A2(_03246_ ), .ZN(_03247_ ) );
INV_X1 _10901_ ( .A(_03247_ ), .ZN(_03248_ ) );
OAI21_X1 _10902_ ( .A(_03241_ ), .B1(_03245_ ), .B2(_03248_ ), .ZN(_03249_ ) );
NAND4_X1 _10903_ ( .A1(_03234_ ), .A2(_03087_ ), .A3(_03098_ ), .A4(_03236_ ), .ZN(_03250_ ) );
INV_X1 _10904_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03251_ ) );
NOR2_X1 _10905_ ( .A1(_03250_ ), .A2(_03251_ ), .ZN(_03252_ ) );
AND3_X1 _10906_ ( .A1(_03252_ ), .A2(_03233_ ), .A3(_03064_ ), .ZN(_03253_ ) );
AND2_X1 _10907_ ( .A1(_03252_ ), .A2(_03247_ ), .ZN(_03254_ ) );
OR2_X1 _10908_ ( .A1(_03253_ ), .A2(_03254_ ), .ZN(_03255_ ) );
NOR2_X1 _10909_ ( .A1(_03249_ ), .A2(_03255_ ), .ZN(_03256_ ) );
NAND3_X1 _10910_ ( .A1(_03086_ ), .A2(_03087_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03257_ ) );
NOR3_X1 _10911_ ( .A1(_03257_ ), .A2(_03080_ ), .A3(\IF_ID_inst [29] ), .ZN(_03258_ ) );
AND2_X1 _10912_ ( .A1(_03258_ ), .A2(_03237_ ), .ZN(_03259_ ) );
AND2_X1 _10913_ ( .A1(_03259_ ), .A2(_03247_ ), .ZN(_03260_ ) );
INV_X1 _10914_ ( .A(_03260_ ), .ZN(_03261_ ) );
NOR2_X1 _10915_ ( .A1(_03164_ ), .A2(\IF_ID_inst [5] ), .ZN(_03262_ ) );
AND3_X1 _10916_ ( .A1(_03262_ ), .A2(_03066_ ), .A3(_03067_ ), .ZN(_03263_ ) );
AND2_X1 _10917_ ( .A1(_03263_ ), .A2(_03143_ ), .ZN(_03264_ ) );
NAND2_X1 _10918_ ( .A1(_03240_ ), .A2(_03264_ ), .ZN(_03265_ ) );
NAND2_X1 _10919_ ( .A1(_03259_ ), .A2(_03264_ ), .ZN(_03266_ ) );
NAND4_X1 _10920_ ( .A1(_03235_ ), .A2(_03263_ ), .A3(_03143_ ), .A4(_03237_ ), .ZN(_03267_ ) );
NAND3_X1 _10921_ ( .A1(_03265_ ), .A2(_03266_ ), .A3(_03267_ ), .ZN(_03268_ ) );
AND2_X1 _10922_ ( .A1(_03233_ ), .A2(_03064_ ), .ZN(_03269_ ) );
AND2_X1 _10923_ ( .A1(_03258_ ), .A2(_03239_ ), .ZN(_03270_ ) );
OR2_X1 _10924_ ( .A1(_03270_ ), .A2(_03244_ ), .ZN(_03271_ ) );
AOI21_X1 _10925_ ( .A(_03268_ ), .B1(_03269_ ), .B2(_03271_ ), .ZN(_03272_ ) );
NAND3_X1 _10926_ ( .A1(_03256_ ), .A2(_03261_ ), .A3(_03272_ ), .ZN(_03273_ ) );
NOR2_X1 _10927_ ( .A1(_03232_ ), .A2(_03273_ ), .ZN(_03274_ ) );
AND2_X1 _10928_ ( .A1(_03233_ ), .A2(_03124_ ), .ZN(_03275_ ) );
AND2_X1 _10929_ ( .A1(_03275_ ), .A2(_03140_ ), .ZN(_03276_ ) );
AND3_X1 _10930_ ( .A1(_03063_ ), .A2(_03096_ ), .A3(_03127_ ), .ZN(_03277_ ) );
AND2_X1 _10931_ ( .A1(_03277_ ), .A2(_03163_ ), .ZN(_03278_ ) );
NOR2_X1 _10932_ ( .A1(_03276_ ), .A2(_03278_ ), .ZN(_03279_ ) );
NAND2_X1 _10933_ ( .A1(_03275_ ), .A2(_03139_ ), .ZN(_03280_ ) );
AND2_X1 _10934_ ( .A1(_03125_ ), .A2(_03069_ ), .ZN(_03281_ ) );
AND2_X1 _10935_ ( .A1(_03281_ ), .A2(_03132_ ), .ZN(_03282_ ) );
AND2_X1 _10936_ ( .A1(_03281_ ), .A2(_03127_ ), .ZN(_03283_ ) );
NOR2_X1 _10937_ ( .A1(_03282_ ), .A2(_03283_ ), .ZN(_03284_ ) );
NAND3_X1 _10938_ ( .A1(_03279_ ), .A2(_03280_ ), .A3(_03284_ ), .ZN(_03285_ ) );
AND2_X2 _10939_ ( .A1(_03233_ ), .A2(_03262_ ), .ZN(_03286_ ) );
AND4_X1 _10940_ ( .A1(\IF_ID_inst [4] ), .A2(_03095_ ), .A3(_03062_ ), .A4(\IF_ID_inst [12] ), .ZN(_03287_ ) );
AND2_X1 _10941_ ( .A1(_03069_ ), .A2(_03287_ ), .ZN(_03288_ ) );
AND2_X1 _10942_ ( .A1(_03288_ ), .A2(\IF_ID_inst [13] ), .ZN(_03289_ ) );
OR2_X1 _10943_ ( .A1(_03286_ ), .A2(_03289_ ), .ZN(_03290_ ) );
NOR2_X1 _10944_ ( .A1(_03285_ ), .A2(_03290_ ), .ZN(_03291_ ) );
AND2_X1 _10945_ ( .A1(_03291_ ), .A2(_03074_ ), .ZN(_03292_ ) );
AND2_X1 _10946_ ( .A1(_03274_ ), .A2(_03292_ ), .ZN(_03293_ ) );
AND2_X2 _10947_ ( .A1(_03150_ ), .A2(_03167_ ), .ZN(_03294_ ) );
AND2_X1 _10948_ ( .A1(_03293_ ), .A2(_03294_ ), .ZN(_03295_ ) );
BUF_X4 _10949_ ( .A(_03295_ ), .Z(_03296_ ) );
AOI211_X1 _10950_ ( .A(_03219_ ), .B(_03296_ ), .C1(\IF_ID_inst [18] ), .C2(_03294_ ), .ZN(_03297_ ) );
NOR2_X1 _10951_ ( .A1(_03295_ ), .A2(_03218_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _10952_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_03298_ ) );
AOI211_X1 _10953_ ( .A(_03091_ ), .B(_03297_ ), .C1(_02141_ ), .C2(_03298_ ), .ZN(_00217_ ) );
AND4_X1 _10954_ ( .A1(\IF_ID_inst [16] ), .A2(_03150_ ), .A3(_03149_ ), .A4(_03167_ ), .ZN(_00218_ ) );
AOI211_X1 _10955_ ( .A(_03219_ ), .B(_03296_ ), .C1(\IF_ID_inst [17] ), .C2(_03294_ ), .ZN(_03299_ ) );
OAI21_X1 _10956_ ( .A(_03151_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [2] ), .ZN(_03300_ ) );
NOR2_X1 _10957_ ( .A1(_03299_ ), .A2(_03300_ ), .ZN(_00219_ ) );
AND4_X1 _10958_ ( .A1(\IF_ID_inst [15] ), .A2(_03150_ ), .A3(_03149_ ), .A4(_03167_ ), .ZN(_00220_ ) );
AOI211_X1 _10959_ ( .A(_03219_ ), .B(_03296_ ), .C1(\IF_ID_inst [16] ), .C2(_03294_ ), .ZN(_03301_ ) );
OAI21_X1 _10960_ ( .A(_03151_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [1] ), .ZN(_03302_ ) );
NOR2_X1 _10961_ ( .A1(_03301_ ), .A2(_03302_ ), .ZN(_00221_ ) );
AOI221_X4 _10962_ ( .A(_03278_ ), .B1(_03286_ ), .B2(_03128_ ), .C1(_03140_ ), .C2(_03275_ ), .ZN(_03303_ ) );
AND4_X1 _10963_ ( .A1(\IF_ID_inst [12] ), .A2(_03127_ ), .A3(_03124_ ), .A4(_03062_ ), .ZN(_03304_ ) );
AND2_X1 _10964_ ( .A1(_03304_ ), .A2(_03123_ ), .ZN(_03305_ ) );
AOI21_X1 _10965_ ( .A(_03305_ ), .B1(_03154_ ), .B2(_03156_ ), .ZN(_03306_ ) );
AND3_X1 _10966_ ( .A1(_03108_ ), .A2(_03109_ ), .A3(_03106_ ), .ZN(_03307_ ) );
AND3_X1 _10967_ ( .A1(_03307_ ), .A2(_03081_ ), .A3(\IF_ID_inst [20] ), .ZN(_03308_ ) );
NOR2_X1 _10968_ ( .A1(_03118_ ), .A2(_03119_ ), .ZN(_03309_ ) );
NAND3_X1 _10969_ ( .A1(_03154_ ), .A2(_03308_ ), .A3(_03309_ ), .ZN(_03310_ ) );
INV_X1 _10970_ ( .A(_03160_ ), .ZN(_03311_ ) );
AND2_X1 _10971_ ( .A1(_03310_ ), .A2(_03311_ ), .ZN(_03312_ ) );
NAND4_X1 _10972_ ( .A1(_03303_ ), .A2(_03074_ ), .A3(_03306_ ), .A4(_03312_ ), .ZN(_03313_ ) );
AND2_X1 _10973_ ( .A1(_03284_ ), .A2(_03280_ ), .ZN(_03314_ ) );
AND2_X1 _10974_ ( .A1(_03286_ ), .A2(_03140_ ), .ZN(_03315_ ) );
NOR2_X1 _10975_ ( .A1(_03315_ ), .A2(_03166_ ), .ZN(_03316_ ) );
AND3_X1 _10976_ ( .A1(_03265_ ), .A2(_03266_ ), .A3(_03267_ ), .ZN(_03317_ ) );
AND3_X1 _10977_ ( .A1(_03263_ ), .A2(\IF_ID_inst [13] ), .A3(_03143_ ), .ZN(_03318_ ) );
AOI21_X1 _10978_ ( .A(_03318_ ), .B1(_03286_ ), .B2(\IF_ID_inst [14] ), .ZN(_03319_ ) );
NAND4_X1 _10979_ ( .A1(_03314_ ), .A2(_03316_ ), .A3(_03317_ ), .A4(_03319_ ), .ZN(_03320_ ) );
NOR4_X1 _10980_ ( .A1(_03313_ ), .A2(_03320_ ), .A3(_03090_ ), .A4(_03091_ ), .ZN(_00222_ ) );
AOI211_X1 _10981_ ( .A(_03219_ ), .B(_03296_ ), .C1(\IF_ID_inst [15] ), .C2(_03294_ ), .ZN(_03321_ ) );
OAI21_X1 _10982_ ( .A(_03151_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [0] ), .ZN(_03322_ ) );
NOR2_X1 _10983_ ( .A1(_03321_ ), .A2(_03322_ ), .ZN(_00223_ ) );
NOR4_X1 _10984_ ( .A1(_03313_ ), .A2(_03320_ ), .A3(_03092_ ), .A4(_03091_ ), .ZN(_00224_ ) );
NOR4_X1 _10985_ ( .A1(_03313_ ), .A2(_03320_ ), .A3(_03093_ ), .A4(_03091_ ), .ZN(_00225_ ) );
INV_X1 _10986_ ( .A(_03295_ ), .ZN(_03323_ ) );
NOR2_X1 _10987_ ( .A1(_03313_ ), .A2(_03320_ ), .ZN(_03324_ ) );
NAND4_X1 _10988_ ( .A1(_03323_ ), .A2(\IF_ID_inst [23] ), .A3(_03217_ ), .A4(_03324_ ), .ZN(_03325_ ) );
OAI21_X1 _10989_ ( .A(\ID_EX_rs2 [3] ), .B1(_03296_ ), .B2(_03219_ ), .ZN(_03326_ ) );
AOI21_X1 _10990_ ( .A(_03082_ ), .B1(_03325_ ), .B2(_03326_ ), .ZN(_00226_ ) );
NOR4_X1 _10991_ ( .A1(_03313_ ), .A2(_03320_ ), .A3(_03081_ ), .A4(_03091_ ), .ZN(_00227_ ) );
NAND4_X1 _10992_ ( .A1(_03323_ ), .A2(\IF_ID_inst [22] ), .A3(_03217_ ), .A4(_03324_ ), .ZN(_03327_ ) );
OAI21_X1 _10993_ ( .A(\ID_EX_rs2 [2] ), .B1(_03296_ ), .B2(_03219_ ), .ZN(_03328_ ) );
AOI21_X1 _10994_ ( .A(_03082_ ), .B1(_03327_ ), .B2(_03328_ ), .ZN(_00228_ ) );
NOR4_X1 _10995_ ( .A1(_03313_ ), .A2(_03320_ ), .A3(_03084_ ), .A4(_03078_ ), .ZN(_00229_ ) );
NAND4_X1 _10996_ ( .A1(_03323_ ), .A2(\IF_ID_inst [21] ), .A3(_03217_ ), .A4(_03324_ ), .ZN(_03329_ ) );
OAI21_X1 _10997_ ( .A(\ID_EX_rs2 [1] ), .B1(_03296_ ), .B2(_03219_ ), .ZN(_03330_ ) );
AOI21_X1 _10998_ ( .A(_03082_ ), .B1(_03329_ ), .B2(_03330_ ), .ZN(_00230_ ) );
INV_X1 _10999_ ( .A(IDU_valid_EXU ), .ZN(_03331_ ) );
AND4_X1 _11000_ ( .A1(_03331_ ), .A2(_03151_ ), .A3(_03123_ ), .A4(_03304_ ), .ZN(_00231_ ) );
OAI21_X1 _11001_ ( .A(_03151_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs2 [0] ), .ZN(_03332_ ) );
AOI221_X4 _11002_ ( .A(_03218_ ), .B1(\IF_ID_inst [20] ), .B2(_03324_ ), .C1(_03294_ ), .C2(_03293_ ), .ZN(_03333_ ) );
NOR2_X1 _11003_ ( .A1(_03332_ ), .A2(_03333_ ), .ZN(_00232_ ) );
INV_X1 _11004_ ( .A(_03292_ ), .ZN(_03334_ ) );
XNOR2_X1 _11005_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_03335_ ) );
XNOR2_X1 _11006_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_03336_ ) );
XNOR2_X1 _11007_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_03337_ ) );
XNOR2_X1 _11008_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_03338_ ) );
NAND4_X1 _11009_ ( .A1(_03335_ ), .A2(_03336_ ), .A3(_03337_ ), .A4(_03338_ ), .ZN(_03339_ ) );
XOR2_X1 _11010_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .Z(_03340_ ) );
NOR2_X1 _11011_ ( .A1(_03339_ ), .A2(_03340_ ), .ZN(_03341_ ) );
AND2_X1 _11012_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03342_ ) );
INV_X1 _11013_ ( .A(\ID_EX_typ [7] ), .ZN(_03343_ ) );
AND2_X1 _11014_ ( .A1(_03342_ ), .A2(_03343_ ), .ZN(_03344_ ) );
AND2_X1 _11015_ ( .A1(_03341_ ), .A2(_03344_ ), .ZN(_03345_ ) );
INV_X1 _11016_ ( .A(_03345_ ), .ZN(_03346_ ) );
XNOR2_X1 _11017_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_03347_ ) );
XNOR2_X1 _11018_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_03348_ ) );
XNOR2_X1 _11019_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_03349_ ) );
XNOR2_X1 _11020_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_03350_ ) );
AND4_X1 _11021_ ( .A1(_03347_ ), .A2(_03348_ ), .A3(_03349_ ), .A4(_03350_ ), .ZN(_03351_ ) );
XNOR2_X1 _11022_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_03352_ ) );
NAND3_X1 _11023_ ( .A1(_03351_ ), .A2(_03344_ ), .A3(_03352_ ), .ZN(_03353_ ) );
AND2_X1 _11024_ ( .A1(_03346_ ), .A2(_03353_ ), .ZN(_03354_ ) );
INV_X1 _11025_ ( .A(_03354_ ), .ZN(_03355_ ) );
AND3_X1 _11026_ ( .A1(_03355_ ), .A2(_03150_ ), .A3(_03167_ ), .ZN(_03356_ ) );
OAI211_X1 _11027_ ( .A(IDU_ready_IFU ), .B(_03149_ ), .C1(_03334_ ), .C2(_03356_ ), .ZN(_03357_ ) );
AOI21_X1 _11028_ ( .A(_03357_ ), .B1(_03334_ ), .B2(_03346_ ), .ZN(_00233_ ) );
AND4_X1 _11029_ ( .A1(_03064_ ), .A2(_03063_ ), .A3(_03128_ ), .A4(_03152_ ), .ZN(_03358_ ) );
AND3_X1 _11030_ ( .A1(_03358_ ), .A2(_03070_ ), .A3(_03103_ ), .ZN(_03359_ ) );
AND3_X1 _11031_ ( .A1(_03307_ ), .A2(_03081_ ), .A3(_03084_ ), .ZN(_03360_ ) );
NAND3_X1 _11032_ ( .A1(_03359_ ), .A2(_03309_ ), .A3(_03360_ ), .ZN(_03361_ ) );
AND2_X1 _11033_ ( .A1(_03361_ ), .A2(_03074_ ), .ZN(_03362_ ) );
NOR2_X1 _11034_ ( .A1(_03161_ ), .A2(_03278_ ), .ZN(_03363_ ) );
AND4_X1 _11035_ ( .A1(_03116_ ), .A2(_03362_ ), .A3(_03129_ ), .A4(_03363_ ), .ZN(_03364_ ) );
AOI21_X1 _11036_ ( .A(_03082_ ), .B1(_03364_ ), .B2(_03223_ ), .ZN(_00234_ ) );
OAI21_X1 _11037_ ( .A(_03128_ ), .B1(_03226_ ), .B2(_03144_ ), .ZN(_03365_ ) );
AND2_X1 _11038_ ( .A1(_03229_ ), .A2(_03365_ ), .ZN(_03366_ ) );
INV_X1 _11039_ ( .A(_03276_ ), .ZN(_03367_ ) );
AND4_X1 _11040_ ( .A1(_03366_ ), .A2(_03367_ ), .A3(_03280_ ), .A4(_03284_ ), .ZN(_03368_ ) );
AOI21_X1 _11041_ ( .A(_03082_ ), .B1(_03368_ ), .B2(_03362_ ), .ZN(_00235_ ) );
AND2_X1 _11042_ ( .A1(_03269_ ), .A2(_03238_ ), .ZN(_03369_ ) );
INV_X1 _11043_ ( .A(_03369_ ), .ZN(_03370_ ) );
AND3_X1 _11044_ ( .A1(_03098_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03236_ ), .ZN(_03371_ ) );
OAI211_X1 _11045_ ( .A(_03242_ ), .B(_03371_ ), .C1(_03269_ ), .C2(_03247_ ), .ZN(_03372_ ) );
NAND2_X1 _11046_ ( .A1(_03370_ ), .A2(_03372_ ), .ZN(_03373_ ) );
NOR2_X1 _11047_ ( .A1(_03245_ ), .A2(_03248_ ), .ZN(_03374_ ) );
AND3_X1 _11048_ ( .A1(_03240_ ), .A2(_03064_ ), .A3(_03233_ ), .ZN(_03375_ ) );
NOR3_X1 _11049_ ( .A1(_03373_ ), .A2(_03374_ ), .A3(_03375_ ), .ZN(_03376_ ) );
NAND2_X1 _11050_ ( .A1(_03286_ ), .A2(_03128_ ), .ZN(_03377_ ) );
AND3_X1 _11051_ ( .A1(_03359_ ), .A2(_03309_ ), .A3(_03360_ ), .ZN(_03378_ ) );
NOR3_X1 _11052_ ( .A1(_03276_ ), .A2(_03378_ ), .A3(_03260_ ), .ZN(_03379_ ) );
NAND3_X1 _11053_ ( .A1(_03244_ ), .A2(_03064_ ), .A3(_03233_ ), .ZN(_03380_ ) );
NAND4_X1 _11054_ ( .A1(_03233_ ), .A2(_03064_ ), .A3(_03258_ ), .A4(_03239_ ), .ZN(_03381_ ) );
AND2_X1 _11055_ ( .A1(_03380_ ), .A2(_03381_ ), .ZN(_03382_ ) );
AND4_X1 _11056_ ( .A1(_03377_ ), .A2(_03379_ ), .A3(_03382_ ), .A4(_03319_ ), .ZN(_03383_ ) );
AND4_X1 _11057_ ( .A1(_03376_ ), .A2(_03383_ ), .A3(_03314_ ), .A4(_03363_ ), .ZN(_03384_ ) );
OAI21_X1 _11058_ ( .A(_03288_ ), .B1(_03238_ ), .B2(_03259_ ), .ZN(_03385_ ) );
NAND3_X1 _11059_ ( .A1(_03288_ ), .A2(_03235_ ), .A3(_03239_ ), .ZN(_03386_ ) );
AND2_X1 _11060_ ( .A1(_03385_ ), .A2(_03386_ ), .ZN(_03387_ ) );
AND2_X1 _11061_ ( .A1(_03316_ ), .A2(_03387_ ), .ZN(_03388_ ) );
AOI21_X1 _11062_ ( .A(_03082_ ), .B1(_03384_ ), .B2(_03388_ ), .ZN(_00236_ ) );
INV_X1 _11063_ ( .A(_03305_ ), .ZN(_03389_ ) );
AND3_X1 _11064_ ( .A1(_03319_ ), .A2(_03389_ ), .A3(_03377_ ), .ZN(_03390_ ) );
AOI21_X1 _11065_ ( .A(_03079_ ), .B1(_03388_ ), .B2(_03390_ ), .ZN(_00237_ ) );
AND2_X1 _11066_ ( .A1(_03114_ ), .A2(_03107_ ), .ZN(_03391_ ) );
AND4_X1 _11067_ ( .A1(_03087_ ), .A2(_03391_ ), .A3(_03110_ ), .A4(_03112_ ), .ZN(_03392_ ) );
NAND2_X1 _11068_ ( .A1(_03392_ ), .A2(_03359_ ), .ZN(_03393_ ) );
AND3_X1 _11069_ ( .A1(_03382_ ), .A2(_03229_ ), .A3(_03393_ ), .ZN(_03394_ ) );
AOI21_X1 _11070_ ( .A(_03079_ ), .B1(_03394_ ), .B2(_03316_ ), .ZN(_00238_ ) );
NOR2_X1 _11071_ ( .A1(_03374_ ), .A2(_03260_ ), .ZN(_03395_ ) );
INV_X1 _11072_ ( .A(_03166_ ), .ZN(_03396_ ) );
OAI21_X1 _11073_ ( .A(_03140_ ), .B1(_03275_ ), .B2(_03264_ ), .ZN(_03397_ ) );
AND4_X1 _11074_ ( .A1(_03229_ ), .A2(_03395_ ), .A3(_03396_ ), .A4(_03397_ ), .ZN(_03398_ ) );
AOI221_X4 _11075_ ( .A(_03268_ ), .B1(\IF_ID_inst [14] ), .B2(_03097_ ), .C1(\IF_ID_inst [13] ), .C2(_03073_ ), .ZN(_03399_ ) );
AOI21_X1 _11076_ ( .A(_03079_ ), .B1(_03398_ ), .B2(_03399_ ), .ZN(_00239_ ) );
NAND2_X1 _11077_ ( .A1(_03266_ ), .A2(_03267_ ), .ZN(_03400_ ) );
AOI211_X1 _11078_ ( .A(_03071_ ), .B(_03400_ ), .C1(\IF_ID_inst [14] ), .C2(_03286_ ), .ZN(_03401_ ) );
OAI21_X1 _11079_ ( .A(_03237_ ), .B1(_03235_ ), .B2(_03258_ ), .ZN(_03402_ ) );
NOR2_X1 _11080_ ( .A1(_03402_ ), .A2(_03248_ ), .ZN(_03403_ ) );
AND3_X1 _11081_ ( .A1(_03062_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_03404_ ) );
AOI21_X1 _11082_ ( .A(_03403_ ), .B1(_03163_ ), .B2(_03404_ ), .ZN(_03405_ ) );
AOI221_X4 _11083_ ( .A(_03225_ ), .B1(_03281_ ), .B2(_03132_ ), .C1(\IF_ID_inst [14] ), .C2(_03134_ ), .ZN(_03406_ ) );
AND4_X1 _11084_ ( .A1(_03370_ ), .A2(_03401_ ), .A3(_03405_ ), .A4(_03406_ ), .ZN(_03407_ ) );
NOR3_X1 _11085_ ( .A1(_03253_ ), .A2(_03228_ ), .A3(_03283_ ), .ZN(_03408_ ) );
AOI21_X1 _11086_ ( .A(_03079_ ), .B1(_03407_ ), .B2(_03408_ ), .ZN(_00240_ ) );
AOI22_X1 _11087_ ( .A1(_03269_ ), .A2(_03238_ ), .B1(_03247_ ), .B2(_03252_ ), .ZN(_03409_ ) );
NAND3_X1 _11088_ ( .A1(_03263_ ), .A2(_03098_ ), .A3(_03143_ ), .ZN(_03410_ ) );
OAI21_X1 _11089_ ( .A(_03098_ ), .B1(_03134_ ), .B2(_03073_ ), .ZN(_03411_ ) );
AND3_X1 _11090_ ( .A1(_03409_ ), .A2(_03410_ ), .A3(_03411_ ), .ZN(_03412_ ) );
OAI21_X1 _11091_ ( .A(_03247_ ), .B1(_03240_ ), .B2(_03259_ ), .ZN(_03413_ ) );
NAND3_X1 _11092_ ( .A1(_03413_ ), .A2(_03380_ ), .A3(_03265_ ), .ZN(_03414_ ) );
AOI21_X1 _11093_ ( .A(_03414_ ), .B1(_03132_ ), .B2(_03286_ ), .ZN(_03415_ ) );
AOI22_X1 _11094_ ( .A1(_03097_ ), .A2(_03128_ ), .B1(_03140_ ), .B2(_03226_ ), .ZN(_03416_ ) );
NAND3_X1 _11095_ ( .A1(_03070_ ), .A2(_03072_ ), .A3(_03132_ ), .ZN(_03417_ ) );
NAND2_X1 _11096_ ( .A1(_03275_ ), .A2(_03132_ ), .ZN(_03418_ ) );
INV_X1 _11097_ ( .A(_03282_ ), .ZN(_03419_ ) );
NAND3_X1 _11098_ ( .A1(_03065_ ), .A2(\IF_ID_inst [14] ), .A3(_03070_ ), .ZN(_03420_ ) );
AND4_X1 _11099_ ( .A1(_03417_ ), .A2(_03418_ ), .A3(_03419_ ), .A4(_03420_ ), .ZN(_03421_ ) );
AND4_X1 _11100_ ( .A1(_03412_ ), .A2(_03415_ ), .A3(_03416_ ), .A4(_03421_ ), .ZN(_03422_ ) );
AOI21_X1 _11101_ ( .A(_03278_ ), .B1(_03097_ ), .B2(_03098_ ), .ZN(_03423_ ) );
AND4_X1 _11102_ ( .A1(_03310_ ), .A2(_03423_ ), .A3(_03227_ ), .A4(_03266_ ), .ZN(_03424_ ) );
AOI21_X1 _11103_ ( .A(_03079_ ), .B1(_03422_ ), .B2(_03424_ ), .ZN(_00241_ ) );
INV_X1 _11104_ ( .A(_03210_ ), .ZN(_03425_ ) );
INV_X1 _11105_ ( .A(\myifu.to_reset ), .ZN(_03426_ ) );
BUF_X4 _11106_ ( .A(_03426_ ), .Z(_03427_ ) );
NAND4_X1 _11107_ ( .A1(_03425_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_03427_ ), .ZN(_03428_ ) );
NAND2_X1 _11108_ ( .A1(\mtvec [0] ), .A2(\myifu.to_reset ), .ZN(_03429_ ) );
AOI21_X1 _11109_ ( .A(fanout_net_2 ), .B1(_03428_ ), .B2(_03429_ ), .ZN(_00245_ ) );
NOR4_X1 _11110_ ( .A1(_03076_ ), .A2(_03095_ ), .A3(\IF_ID_inst [4] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03430_ ) );
AND2_X1 _11111_ ( .A1(_03430_ ), .A2(_03069_ ), .ZN(_03431_ ) );
AND2_X1 _11112_ ( .A1(_03431_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03432_ ) );
OAI211_X1 _11113_ ( .A(_03159_ ), .B(\IF_ID_inst [31] ), .C1(_03069_ ), .C2(_03123_ ), .ZN(_03433_ ) );
NOR2_X1 _11114_ ( .A1(_03432_ ), .A2(_03433_ ), .ZN(_03434_ ) );
BUF_X4 _11115_ ( .A(_03434_ ), .Z(_03435_ ) );
XNOR2_X1 _11116_ ( .A(_03435_ ), .B(_01757_ ), .ZN(_03436_ ) );
AND2_X1 _11117_ ( .A1(_03160_ ), .A2(\IF_ID_inst [20] ), .ZN(_03437_ ) );
INV_X1 _11118_ ( .A(_03437_ ), .ZN(_03438_ ) );
INV_X1 _11119_ ( .A(_03431_ ), .ZN(_03439_ ) );
OAI21_X1 _11120_ ( .A(_03438_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03439_ ), .ZN(_03440_ ) );
XNOR2_X1 _11121_ ( .A(_03440_ ), .B(_01782_ ), .ZN(_03441_ ) );
OAI21_X1 _11122_ ( .A(_03439_ ), .B1(_03311_ ), .B2(_03142_ ), .ZN(_03442_ ) );
INV_X1 _11123_ ( .A(_03432_ ), .ZN(_03443_ ) );
NAND2_X1 _11124_ ( .A1(_03442_ ), .A2(_03443_ ), .ZN(_03444_ ) );
XNOR2_X1 _11125_ ( .A(_03444_ ), .B(\IF_ID_pc [12] ), .ZN(_03445_ ) );
AND2_X1 _11126_ ( .A1(_03441_ ), .A2(_03445_ ), .ZN(_03446_ ) );
AND2_X1 _11127_ ( .A1(_03160_ ), .A2(\IF_ID_inst [29] ), .ZN(_03447_ ) );
INV_X1 _11128_ ( .A(_03447_ ), .ZN(_03448_ ) );
OAI21_X1 _11129_ ( .A(_03448_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03439_ ), .ZN(_03449_ ) );
INV_X1 _11130_ ( .A(\IF_ID_pc [9] ), .ZN(_03450_ ) );
XNOR2_X1 _11131_ ( .A(_03449_ ), .B(_03450_ ), .ZN(_03451_ ) );
AND2_X1 _11132_ ( .A1(_03160_ ), .A2(\IF_ID_inst [30] ), .ZN(_03452_ ) );
INV_X1 _11133_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03453_ ) );
BUF_X4 _11134_ ( .A(_03431_ ), .Z(_03454_ ) );
AOI21_X1 _11135_ ( .A(_03452_ ), .B1(_03453_ ), .B2(_03454_ ), .ZN(_03455_ ) );
XNOR2_X1 _11136_ ( .A(_03455_ ), .B(\IF_ID_pc [10] ), .ZN(_03456_ ) );
AND3_X1 _11137_ ( .A1(_03446_ ), .A2(_03451_ ), .A3(_03456_ ), .ZN(_03457_ ) );
NAND3_X1 _11138_ ( .A1(_03159_ ), .A2(\IF_ID_inst [16] ), .A3(_03123_ ), .ZN(_03458_ ) );
AOI21_X1 _11139_ ( .A(_03432_ ), .B1(_03439_ ), .B2(_03458_ ), .ZN(_03459_ ) );
XOR2_X1 _11140_ ( .A(_03459_ ), .B(\IF_ID_pc [16] ), .Z(_03460_ ) );
AND3_X1 _11141_ ( .A1(_03159_ ), .A2(\IF_ID_inst [15] ), .A3(_03122_ ), .ZN(_03461_ ) );
MUX2_X1 _11142_ ( .A(_03461_ ), .B(_03251_ ), .S(_03454_ ), .Z(_03462_ ) );
INV_X1 _11143_ ( .A(\IF_ID_pc [15] ), .ZN(_03463_ ) );
XNOR2_X1 _11144_ ( .A(_03462_ ), .B(_03463_ ), .ZN(_03464_ ) );
AND2_X1 _11145_ ( .A1(_03460_ ), .A2(_03464_ ), .ZN(_03465_ ) );
OAI21_X1 _11146_ ( .A(_03439_ ), .B1(_03311_ ), .B2(_03131_ ), .ZN(_03466_ ) );
AND3_X1 _11147_ ( .A1(_03466_ ), .A2(\IF_ID_pc [14] ), .A3(_03443_ ), .ZN(_03467_ ) );
AOI21_X1 _11148_ ( .A(\IF_ID_pc [14] ), .B1(_03466_ ), .B2(_03443_ ), .ZN(_03468_ ) );
NOR2_X1 _11149_ ( .A1(_03467_ ), .A2(_03468_ ), .ZN(_03469_ ) );
NAND3_X1 _11150_ ( .A1(_03159_ ), .A2(\IF_ID_inst [13] ), .A3(_03123_ ), .ZN(_03470_ ) );
MUX2_X1 _11151_ ( .A(_03470_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .S(_03454_ ), .Z(_03471_ ) );
XNOR2_X1 _11152_ ( .A(_03471_ ), .B(\IF_ID_pc [13] ), .ZN(_03472_ ) );
AND2_X1 _11153_ ( .A1(_03469_ ), .A2(_03472_ ), .ZN(_03473_ ) );
NAND3_X1 _11154_ ( .A1(_03457_ ), .A2(_03465_ ), .A3(_03473_ ), .ZN(_03474_ ) );
AND2_X1 _11155_ ( .A1(_03160_ ), .A2(\IF_ID_inst [26] ), .ZN(_03475_ ) );
INV_X1 _11156_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03476_ ) );
AOI21_X1 _11157_ ( .A(_03475_ ), .B1(_03476_ ), .B2(_03454_ ), .ZN(_03477_ ) );
INV_X1 _11158_ ( .A(\IF_ID_pc [6] ), .ZN(_03478_ ) );
OR2_X1 _11159_ ( .A1(_03477_ ), .A2(_03478_ ), .ZN(_03479_ ) );
AND2_X1 _11160_ ( .A1(_03160_ ), .A2(\IF_ID_inst [25] ), .ZN(_03480_ ) );
NOR2_X1 _11161_ ( .A1(_03439_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03481_ ) );
NOR2_X1 _11162_ ( .A1(_03480_ ), .A2(_03481_ ), .ZN(_03482_ ) );
AND3_X1 _11163_ ( .A1(_03159_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .A3(_03122_ ), .ZN(_03483_ ) );
AND3_X1 _11164_ ( .A1(_03430_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_03068_ ), .ZN(_03484_ ) );
NOR2_X1 _11165_ ( .A1(_03483_ ), .A2(_03484_ ), .ZN(_03485_ ) );
INV_X1 _11166_ ( .A(\IF_ID_pc [2] ), .ZN(_03486_ ) );
XNOR2_X1 _11167_ ( .A(_03485_ ), .B(_03486_ ), .ZN(_03487_ ) );
AND2_X1 _11168_ ( .A1(_03160_ ), .A2(\IF_ID_inst [21] ), .ZN(_03488_ ) );
INV_X1 _11169_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03489_ ) );
AND3_X1 _11170_ ( .A1(_03430_ ), .A2(_03489_ ), .A3(_03068_ ), .ZN(_03490_ ) );
NOR2_X1 _11171_ ( .A1(_03488_ ), .A2(_03490_ ), .ZN(_03491_ ) );
INV_X1 _11172_ ( .A(\IF_ID_pc [1] ), .ZN(_03492_ ) );
NOR2_X1 _11173_ ( .A1(_03491_ ), .A2(_03492_ ), .ZN(_03493_ ) );
AND2_X1 _11174_ ( .A1(_03487_ ), .A2(_03493_ ), .ZN(_03494_ ) );
NOR3_X1 _11175_ ( .A1(_03483_ ), .A2(_03486_ ), .A3(_03484_ ), .ZN(_03495_ ) );
NOR2_X1 _11176_ ( .A1(_03494_ ), .A2(_03495_ ), .ZN(_03496_ ) );
AND2_X1 _11177_ ( .A1(_03160_ ), .A2(\IF_ID_inst [23] ), .ZN(_03497_ ) );
INV_X1 _11178_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03498_ ) );
AND3_X1 _11179_ ( .A1(_03430_ ), .A2(_03498_ ), .A3(_03068_ ), .ZN(_03499_ ) );
NOR2_X1 _11180_ ( .A1(_03497_ ), .A2(_03499_ ), .ZN(_03500_ ) );
INV_X1 _11181_ ( .A(fanout_net_6 ), .ZN(_03501_ ) );
XNOR2_X1 _11182_ ( .A(_03500_ ), .B(_03501_ ), .ZN(_03502_ ) );
OR2_X1 _11183_ ( .A1(_03496_ ), .A2(_03502_ ), .ZN(_03503_ ) );
OR2_X1 _11184_ ( .A1(_03500_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03504_ ) );
INV_X1 _11185_ ( .A(fanout_net_10 ), .ZN(_03505_ ) );
AND2_X1 _11186_ ( .A1(_03160_ ), .A2(\IF_ID_inst [24] ), .ZN(_03506_ ) );
INV_X1 _11187_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03507_ ) );
AOI21_X1 _11188_ ( .A(_03506_ ), .B1(_03507_ ), .B2(_03454_ ), .ZN(_03508_ ) );
AOI22_X1 _11189_ ( .A1(_03503_ ), .A2(_03504_ ), .B1(_03505_ ), .B2(_03508_ ), .ZN(_03509_ ) );
NOR2_X1 _11190_ ( .A1(_03508_ ), .A2(_03505_ ), .ZN(_03510_ ) );
NOR2_X1 _11191_ ( .A1(_03509_ ), .A2(_03510_ ), .ZN(_03511_ ) );
INV_X1 _11192_ ( .A(\IF_ID_pc [5] ), .ZN(_03512_ ) );
XNOR2_X1 _11193_ ( .A(_03482_ ), .B(_03512_ ), .ZN(_03513_ ) );
OAI221_X1 _11194_ ( .A(_03479_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_03482_ ), .C1(_03511_ ), .C2(_03513_ ), .ZN(_03514_ ) );
AND2_X1 _11195_ ( .A1(_03161_ ), .A2(\IF_ID_inst [27] ), .ZN(_03515_ ) );
INV_X1 _11196_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03516_ ) );
AOI21_X1 _11197_ ( .A(_03515_ ), .B1(_03516_ ), .B2(_03454_ ), .ZN(_03517_ ) );
XNOR2_X1 _11198_ ( .A(_03517_ ), .B(\IF_ID_pc [7] ), .ZN(_03518_ ) );
NAND2_X1 _11199_ ( .A1(_03477_ ), .A2(_03478_ ), .ZN(_03519_ ) );
AND3_X1 _11200_ ( .A1(_03514_ ), .A2(_03518_ ), .A3(_03519_ ), .ZN(_03520_ ) );
NOR2_X1 _11201_ ( .A1(_03517_ ), .A2(_01852_ ), .ZN(_03521_ ) );
AND2_X1 _11202_ ( .A1(_03161_ ), .A2(\IF_ID_inst [28] ), .ZN(_03522_ ) );
INV_X1 _11203_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03523_ ) );
AOI21_X1 _11204_ ( .A(_03522_ ), .B1(_03523_ ), .B2(_03454_ ), .ZN(_03524_ ) );
INV_X1 _11205_ ( .A(_03524_ ), .ZN(_03525_ ) );
OAI22_X1 _11206_ ( .A1(_03520_ ), .A2(_03521_ ), .B1(\IF_ID_pc [8] ), .B2(_03525_ ), .ZN(_03526_ ) );
OR2_X1 _11207_ ( .A1(_03524_ ), .A2(_01803_ ), .ZN(_03527_ ) );
AOI21_X1 _11208_ ( .A(_03474_ ), .B1(_03526_ ), .B2(_03527_ ), .ZN(_03528_ ) );
INV_X1 _11209_ ( .A(_03446_ ), .ZN(_03529_ ) );
INV_X1 _11210_ ( .A(\IF_ID_pc [10] ), .ZN(_03530_ ) );
NOR2_X1 _11211_ ( .A1(_03455_ ), .A2(_03530_ ), .ZN(_03531_ ) );
AND2_X1 _11212_ ( .A1(_03455_ ), .A2(_03530_ ), .ZN(_03532_ ) );
INV_X1 _11213_ ( .A(_03532_ ), .ZN(_03533_ ) );
AND2_X1 _11214_ ( .A1(_03449_ ), .A2(\IF_ID_pc [9] ), .ZN(_03534_ ) );
AOI21_X1 _11215_ ( .A(_03531_ ), .B1(_03533_ ), .B2(_03534_ ), .ZN(_03535_ ) );
NOR2_X1 _11216_ ( .A1(_03529_ ), .A2(_03535_ ), .ZN(_03536_ ) );
AND3_X1 _11217_ ( .A1(_03442_ ), .A2(\IF_ID_pc [12] ), .A3(_03443_ ), .ZN(_03537_ ) );
AND2_X1 _11218_ ( .A1(_03440_ ), .A2(\IF_ID_pc [11] ), .ZN(_03538_ ) );
AND2_X1 _11219_ ( .A1(_03445_ ), .A2(_03538_ ), .ZN(_03539_ ) );
OR3_X1 _11220_ ( .A1(_03536_ ), .A2(_03537_ ), .A3(_03539_ ), .ZN(_03540_ ) );
NAND3_X1 _11221_ ( .A1(_03540_ ), .A2(_03465_ ), .A3(_03473_ ), .ZN(_03541_ ) );
INV_X1 _11222_ ( .A(\IF_ID_pc [13] ), .ZN(_03542_ ) );
NOR2_X1 _11223_ ( .A1(_03471_ ), .A2(_03542_ ), .ZN(_03543_ ) );
INV_X1 _11224_ ( .A(_03543_ ), .ZN(_03544_ ) );
NOR3_X1 _11225_ ( .A1(_03544_ ), .A2(_03467_ ), .A3(_03468_ ), .ZN(_03545_ ) );
OAI21_X1 _11226_ ( .A(_03465_ ), .B1(_03467_ ), .B2(_03545_ ), .ZN(_03546_ ) );
AND2_X1 _11227_ ( .A1(_03462_ ), .A2(\IF_ID_pc [15] ), .ZN(_03547_ ) );
AND2_X1 _11228_ ( .A1(_03460_ ), .A2(_03547_ ), .ZN(_03548_ ) );
AOI21_X1 _11229_ ( .A(_03548_ ), .B1(\IF_ID_pc [16] ), .B2(_03459_ ), .ZN(_03549_ ) );
NAND3_X1 _11230_ ( .A1(_03541_ ), .A2(_03546_ ), .A3(_03549_ ), .ZN(_03550_ ) );
NOR2_X1 _11231_ ( .A1(_03528_ ), .A2(_03550_ ), .ZN(_03551_ ) );
XNOR2_X1 _11232_ ( .A(_03434_ ), .B(_01797_ ), .ZN(_03552_ ) );
INV_X1 _11233_ ( .A(_03552_ ), .ZN(_03553_ ) );
AND3_X1 _11234_ ( .A1(_03159_ ), .A2(\IF_ID_inst [19] ), .A3(_03123_ ), .ZN(_03554_ ) );
MUX2_X1 _11235_ ( .A(_03554_ ), .B(_03251_ ), .S(_03454_ ), .Z(_03555_ ) );
XNOR2_X1 _11236_ ( .A(_03555_ ), .B(_01772_ ), .ZN(_03556_ ) );
INV_X1 _11237_ ( .A(_03556_ ), .ZN(_03557_ ) );
AND3_X1 _11238_ ( .A1(_03159_ ), .A2(\IF_ID_inst [18] ), .A3(_03123_ ), .ZN(_03558_ ) );
MUX2_X1 _11239_ ( .A(_03558_ ), .B(_03251_ ), .S(_03454_ ), .Z(_03559_ ) );
XNOR2_X1 _11240_ ( .A(_03559_ ), .B(_01985_ ), .ZN(_03560_ ) );
AND3_X1 _11241_ ( .A1(_03159_ ), .A2(\IF_ID_inst [17] ), .A3(_03123_ ), .ZN(_03561_ ) );
MUX2_X1 _11242_ ( .A(_03561_ ), .B(_03251_ ), .S(_03454_ ), .Z(_03562_ ) );
XNOR2_X1 _11243_ ( .A(_03562_ ), .B(_01957_ ), .ZN(_03563_ ) );
NAND2_X1 _11244_ ( .A1(_03560_ ), .A2(_03563_ ), .ZN(_03564_ ) );
NOR4_X1 _11245_ ( .A1(_03551_ ), .A2(_03553_ ), .A3(_03557_ ), .A4(_03564_ ), .ZN(_03565_ ) );
AND2_X1 _11246_ ( .A1(_03559_ ), .A2(\IF_ID_pc [18] ), .ZN(_03566_ ) );
AND2_X1 _11247_ ( .A1(_03562_ ), .A2(\IF_ID_pc [17] ), .ZN(_03567_ ) );
OR2_X1 _11248_ ( .A1(_03566_ ), .A2(_03567_ ), .ZN(_03568_ ) );
NOR2_X1 _11249_ ( .A1(_03559_ ), .A2(\IF_ID_pc [18] ), .ZN(_03569_ ) );
INV_X1 _11250_ ( .A(_03569_ ), .ZN(_03570_ ) );
AND4_X1 _11251_ ( .A1(_03552_ ), .A2(_03568_ ), .A3(_03556_ ), .A4(_03570_ ), .ZN(_03571_ ) );
NOR3_X1 _11252_ ( .A1(_03432_ ), .A2(_01797_ ), .A3(_03433_ ), .ZN(_03572_ ) );
AND2_X1 _11253_ ( .A1(_03555_ ), .A2(\IF_ID_pc [19] ), .ZN(_03573_ ) );
AND2_X1 _11254_ ( .A1(_03552_ ), .A2(_03573_ ), .ZN(_03574_ ) );
OR3_X1 _11255_ ( .A1(_03571_ ), .A2(_03572_ ), .A3(_03574_ ), .ZN(_03575_ ) );
OR2_X1 _11256_ ( .A1(_03565_ ), .A2(_03575_ ), .ZN(_03576_ ) );
XNOR2_X1 _11257_ ( .A(_03434_ ), .B(_01759_ ), .ZN(_03577_ ) );
XNOR2_X1 _11258_ ( .A(_03434_ ), .B(_01952_ ), .ZN(_03578_ ) );
AND2_X1 _11259_ ( .A1(_03577_ ), .A2(_03578_ ), .ZN(_03579_ ) );
XNOR2_X1 _11260_ ( .A(_03434_ ), .B(\IF_ID_pc [21] ), .ZN(_03580_ ) );
XNOR2_X1 _11261_ ( .A(_03434_ ), .B(\IF_ID_pc [22] ), .ZN(_03581_ ) );
NOR2_X1 _11262_ ( .A1(_03580_ ), .A2(_03581_ ), .ZN(_03582_ ) );
AND3_X1 _11263_ ( .A1(_03576_ ), .A2(_03579_ ), .A3(_03582_ ), .ZN(_03583_ ) );
AND2_X1 _11264_ ( .A1(_03435_ ), .A2(\IF_ID_pc [22] ), .ZN(_03584_ ) );
AND2_X1 _11265_ ( .A1(_03435_ ), .A2(\IF_ID_pc [21] ), .ZN(_03585_ ) );
OAI21_X1 _11266_ ( .A(_03579_ ), .B1(_03584_ ), .B2(_03585_ ), .ZN(_03586_ ) );
NAND2_X1 _11267_ ( .A1(_03435_ ), .A2(\IF_ID_pc [24] ), .ZN(_03587_ ) );
NAND2_X1 _11268_ ( .A1(_03435_ ), .A2(\IF_ID_pc [23] ), .ZN(_03588_ ) );
NAND3_X1 _11269_ ( .A1(_03586_ ), .A2(_03587_ ), .A3(_03588_ ), .ZN(_03589_ ) );
OAI21_X1 _11270_ ( .A(_03436_ ), .B1(_03583_ ), .B2(_03589_ ), .ZN(_03590_ ) );
BUF_X4 _11271_ ( .A(_03435_ ), .Z(_03591_ ) );
XNOR2_X1 _11272_ ( .A(_03591_ ), .B(_01899_ ), .ZN(_03592_ ) );
INV_X1 _11273_ ( .A(_03592_ ), .ZN(_03593_ ) );
NOR2_X1 _11274_ ( .A1(_03590_ ), .A2(_03593_ ), .ZN(_03594_ ) );
XOR2_X1 _11275_ ( .A(_03435_ ), .B(\IF_ID_pc [27] ), .Z(_03595_ ) );
XNOR2_X1 _11276_ ( .A(_03435_ ), .B(_01787_ ), .ZN(_03596_ ) );
AND2_X1 _11277_ ( .A1(_03595_ ), .A2(_03596_ ), .ZN(_03597_ ) );
NAND2_X1 _11278_ ( .A1(_03594_ ), .A2(_03597_ ), .ZN(_03598_ ) );
AND2_X1 _11279_ ( .A1(_03435_ ), .A2(\IF_ID_pc [27] ), .ZN(_03599_ ) );
OAI21_X1 _11280_ ( .A(_03435_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_03600_ ) );
INV_X1 _11281_ ( .A(_03600_ ), .ZN(_03601_ ) );
AOI221_X4 _11282_ ( .A(_03599_ ), .B1(\IF_ID_pc [28] ), .B2(_03591_ ), .C1(_03597_ ), .C2(_03601_ ), .ZN(_03602_ ) );
NAND2_X1 _11283_ ( .A1(_03598_ ), .A2(_03602_ ), .ZN(_03603_ ) );
XNOR2_X1 _11284_ ( .A(_03591_ ), .B(_01875_ ), .ZN(_03604_ ) );
NAND2_X1 _11285_ ( .A1(_03603_ ), .A2(_03604_ ), .ZN(_03605_ ) );
NAND2_X1 _11286_ ( .A1(_03591_ ), .A2(\IF_ID_pc [29] ), .ZN(_03606_ ) );
AND2_X1 _11287_ ( .A1(_03605_ ), .A2(_03606_ ), .ZN(_03607_ ) );
XNOR2_X1 _11288_ ( .A(_03591_ ), .B(\IF_ID_pc [30] ), .ZN(_03608_ ) );
OR2_X1 _11289_ ( .A1(_03607_ ), .A2(_03608_ ), .ZN(_03609_ ) );
AOI21_X1 _11290_ ( .A(_03212_ ), .B1(_03607_ ), .B2(_03608_ ), .ZN(_03610_ ) );
AOI221_X4 _11291_ ( .A(\myifu.to_reset ), .B1(\myexu.pc_jump [30] ), .B2(_03212_ ), .C1(_03609_ ), .C2(_03610_ ), .ZN(_03611_ ) );
BUF_X4 _11292_ ( .A(_03427_ ), .Z(_03612_ ) );
NOR2_X1 _11293_ ( .A1(_03612_ ), .A2(\mtvec [30] ), .ZN(_03613_ ) );
NOR3_X1 _11294_ ( .A1(_03611_ ), .A2(fanout_net_2 ), .A3(_03613_ ), .ZN(_00246_ ) );
BUF_X4 _11295_ ( .A(_03427_ ), .Z(_03614_ ) );
OR3_X1 _11296_ ( .A1(_03210_ ), .A2(_03211_ ), .A3(\myexu.pc_jump [21] ), .ZN(_03615_ ) );
XNOR2_X1 _11297_ ( .A(_03576_ ), .B(_03580_ ), .ZN(_03616_ ) );
BUF_X4 _11298_ ( .A(_03212_ ), .Z(_03617_ ) );
BUF_X4 _11299_ ( .A(_03617_ ), .Z(_03618_ ) );
OAI211_X1 _11300_ ( .A(_03614_ ), .B(_03615_ ), .C1(_03616_ ), .C2(_03618_ ), .ZN(_03619_ ) );
NAND2_X1 _11301_ ( .A1(\mtvec [21] ), .A2(\myifu.to_reset ), .ZN(_03620_ ) );
AOI21_X1 _11302_ ( .A(fanout_net_2 ), .B1(_03619_ ), .B2(_03620_ ), .ZN(_00247_ ) );
NOR2_X1 _11303_ ( .A1(_03427_ ), .A2(\mtvec [20] ), .ZN(_03621_ ) );
NOR2_X1 _11304_ ( .A1(_03551_ ), .A2(_03564_ ), .ZN(_03622_ ) );
INV_X1 _11305_ ( .A(_03622_ ), .ZN(_03623_ ) );
NAND2_X1 _11306_ ( .A1(_03568_ ), .A2(_03570_ ), .ZN(_03624_ ) );
AOI21_X1 _11307_ ( .A(_03557_ ), .B1(_03623_ ), .B2(_03624_ ), .ZN(_03625_ ) );
OR3_X1 _11308_ ( .A1(_03625_ ), .A2(_03573_ ), .A3(_03552_ ), .ZN(_03626_ ) );
INV_X1 _11309_ ( .A(_03212_ ), .ZN(_03627_ ) );
BUF_X4 _11310_ ( .A(_03627_ ), .Z(_03628_ ) );
BUF_X4 _11311_ ( .A(_03628_ ), .Z(_03629_ ) );
BUF_X4 _11312_ ( .A(_03629_ ), .Z(_03630_ ) );
OAI21_X1 _11313_ ( .A(_03552_ ), .B1(_03625_ ), .B2(_03573_ ), .ZN(_03631_ ) );
NAND3_X1 _11314_ ( .A1(_03626_ ), .A2(_03630_ ), .A3(_03631_ ), .ZN(_03632_ ) );
AOI21_X1 _11315_ ( .A(\myifu.to_reset ), .B1(_03618_ ), .B2(\myexu.pc_jump [20] ), .ZN(_03633_ ) );
AOI211_X1 _11316_ ( .A(fanout_net_2 ), .B(_03621_ ), .C1(_03632_ ), .C2(_03633_ ), .ZN(_00248_ ) );
AND2_X1 _11317_ ( .A1(_03623_ ), .A2(_03624_ ), .ZN(_03634_ ) );
XNOR2_X1 _11318_ ( .A(_03634_ ), .B(_03556_ ), .ZN(_03635_ ) );
MUX2_X1 _11319_ ( .A(\myexu.pc_jump [19] ), .B(_03635_ ), .S(_03628_ ), .Z(_03636_ ) );
MUX2_X1 _11320_ ( .A(\mtvec [19] ), .B(_03636_ ), .S(_03427_ ), .Z(_03637_ ) );
AND2_X1 _11321_ ( .A1(_03637_ ), .A2(_01570_ ), .ZN(_00249_ ) );
INV_X1 _11322_ ( .A(_03560_ ), .ZN(_03638_ ) );
INV_X1 _11323_ ( .A(_03457_ ), .ZN(_03639_ ) );
AOI21_X1 _11324_ ( .A(_03639_ ), .B1(_03526_ ), .B2(_03527_ ), .ZN(_03640_ ) );
NOR2_X1 _11325_ ( .A1(_03640_ ), .A2(_03540_ ), .ZN(_03641_ ) );
NAND3_X1 _11326_ ( .A1(_03473_ ), .A2(_03460_ ), .A3(_03464_ ), .ZN(_03642_ ) );
NOR2_X1 _11327_ ( .A1(_03641_ ), .A2(_03642_ ), .ZN(_03643_ ) );
AND2_X1 _11328_ ( .A1(_03459_ ), .A2(\IF_ID_pc [16] ), .ZN(_03644_ ) );
INV_X1 _11329_ ( .A(_03644_ ), .ZN(_03645_ ) );
OAI21_X1 _11330_ ( .A(_03547_ ), .B1(\IF_ID_pc [16] ), .B2(_03459_ ), .ZN(_03646_ ) );
NAND3_X1 _11331_ ( .A1(_03546_ ), .A2(_03645_ ), .A3(_03646_ ), .ZN(_03647_ ) );
OAI21_X1 _11332_ ( .A(_03563_ ), .B1(_03643_ ), .B2(_03647_ ), .ZN(_03648_ ) );
INV_X1 _11333_ ( .A(_03567_ ), .ZN(_03649_ ) );
AOI21_X1 _11334_ ( .A(_03638_ ), .B1(_03648_ ), .B2(_03649_ ), .ZN(_03650_ ) );
OR2_X1 _11335_ ( .A1(_03641_ ), .A2(_03642_ ), .ZN(_03651_ ) );
OR2_X1 _11336_ ( .A1(_03545_ ), .A2(_03467_ ), .ZN(_03652_ ) );
AOI22_X1 _11337_ ( .A1(_03652_ ), .A2(_03465_ ), .B1(\IF_ID_pc [16] ), .B2(_03459_ ), .ZN(_03653_ ) );
NAND3_X1 _11338_ ( .A1(_03651_ ), .A2(_03646_ ), .A3(_03653_ ), .ZN(_03654_ ) );
AOI211_X1 _11339_ ( .A(_03560_ ), .B(_03567_ ), .C1(_03654_ ), .C2(_03563_ ), .ZN(_03655_ ) );
NOR3_X1 _11340_ ( .A1(_03650_ ), .A2(_03655_ ), .A3(_03617_ ), .ZN(_03656_ ) );
AOI211_X1 _11341_ ( .A(\myifu.to_reset ), .B(_03656_ ), .C1(\myexu.pc_jump [18] ), .C2(_03618_ ), .ZN(_03657_ ) );
NOR2_X1 _11342_ ( .A1(_03612_ ), .A2(\mtvec [18] ), .ZN(_03658_ ) );
NOR3_X1 _11343_ ( .A1(_03657_ ), .A2(fanout_net_2 ), .A3(_03658_ ), .ZN(_00250_ ) );
XOR2_X1 _11344_ ( .A(_03551_ ), .B(_03563_ ), .Z(_03659_ ) );
NAND2_X1 _11345_ ( .A1(_03659_ ), .A2(_03629_ ), .ZN(_03660_ ) );
OAI211_X1 _11346_ ( .A(_03660_ ), .B(_03614_ ), .C1(\myexu.pc_jump [17] ), .C2(_03630_ ), .ZN(_03661_ ) );
NAND2_X1 _11347_ ( .A1(\mtvec [17] ), .A2(\myifu.to_reset ), .ZN(_03662_ ) );
AOI21_X1 _11348_ ( .A(fanout_net_2 ), .B1(_03661_ ), .B2(_03662_ ), .ZN(_00251_ ) );
NOR2_X1 _11349_ ( .A1(_03427_ ), .A2(\mtvec [16] ), .ZN(_03663_ ) );
OAI21_X1 _11350_ ( .A(_03473_ ), .B1(_03640_ ), .B2(_03540_ ), .ZN(_03664_ ) );
AOI21_X1 _11351_ ( .A(_03467_ ), .B1(_03469_ ), .B2(_03543_ ), .ZN(_03665_ ) );
NAND2_X1 _11352_ ( .A1(_03664_ ), .A2(_03665_ ), .ZN(_03666_ ) );
AND2_X1 _11353_ ( .A1(_03666_ ), .A2(_03464_ ), .ZN(_03667_ ) );
OR3_X1 _11354_ ( .A1(_03667_ ), .A2(_03460_ ), .A3(_03547_ ), .ZN(_03668_ ) );
OAI21_X1 _11355_ ( .A(_03460_ ), .B1(_03667_ ), .B2(_03547_ ), .ZN(_03669_ ) );
NAND3_X1 _11356_ ( .A1(_03668_ ), .A2(_03630_ ), .A3(_03669_ ), .ZN(_03670_ ) );
AOI21_X1 _11357_ ( .A(\myifu.to_reset ), .B1(_03618_ ), .B2(\myexu.pc_jump [16] ), .ZN(_03671_ ) );
AOI211_X1 _11358_ ( .A(fanout_net_2 ), .B(_03663_ ), .C1(_03670_ ), .C2(_03671_ ), .ZN(_00252_ ) );
NOR2_X1 _11359_ ( .A1(_03666_ ), .A2(_03464_ ), .ZN(_03672_ ) );
OAI21_X1 _11360_ ( .A(_03629_ ), .B1(_03667_ ), .B2(_03672_ ), .ZN(_03673_ ) );
OAI211_X1 _11361_ ( .A(_03673_ ), .B(_03614_ ), .C1(\myexu.pc_jump [15] ), .C2(_03630_ ), .ZN(_03674_ ) );
NAND2_X1 _11362_ ( .A1(\mtvec [15] ), .A2(\myifu.to_reset ), .ZN(_03675_ ) );
AOI21_X1 _11363_ ( .A(fanout_net_2 ), .B1(_03674_ ), .B2(_03675_ ), .ZN(_00253_ ) );
OAI21_X1 _11364_ ( .A(_03472_ ), .B1(_03640_ ), .B2(_03540_ ), .ZN(_03676_ ) );
AND2_X1 _11365_ ( .A1(_03676_ ), .A2(_03544_ ), .ZN(_03677_ ) );
XNOR2_X1 _11366_ ( .A(_03677_ ), .B(_03469_ ), .ZN(_03678_ ) );
MUX2_X1 _11367_ ( .A(\myexu.pc_jump [14] ), .B(_03678_ ), .S(_03628_ ), .Z(_03679_ ) );
MUX2_X1 _11368_ ( .A(\mtvec [14] ), .B(_03679_ ), .S(_03426_ ), .Z(_03680_ ) );
AND2_X1 _11369_ ( .A1(_03680_ ), .A2(_01570_ ), .ZN(_00254_ ) );
XOR2_X1 _11370_ ( .A(_03641_ ), .B(_03472_ ), .Z(_03681_ ) );
NAND2_X1 _11371_ ( .A1(_03681_ ), .A2(_03629_ ), .ZN(_03682_ ) );
OAI211_X1 _11372_ ( .A(_03682_ ), .B(_03614_ ), .C1(\myexu.pc_jump [13] ), .C2(_03630_ ), .ZN(_03683_ ) );
NAND2_X1 _11373_ ( .A1(\mtvec [13] ), .A2(\myifu.to_reset ), .ZN(_03684_ ) );
AOI21_X1 _11374_ ( .A(fanout_net_2 ), .B1(_03683_ ), .B2(_03684_ ), .ZN(_00255_ ) );
NOR2_X1 _11375_ ( .A1(_03427_ ), .A2(\mtvec [12] ), .ZN(_03685_ ) );
INV_X1 _11376_ ( .A(_03451_ ), .ZN(_03686_ ) );
AOI21_X1 _11377_ ( .A(_03686_ ), .B1(_03526_ ), .B2(_03527_ ), .ZN(_03687_ ) );
NOR2_X1 _11378_ ( .A1(_03687_ ), .A2(_03534_ ), .ZN(_03688_ ) );
OAI21_X1 _11379_ ( .A(_03688_ ), .B1(_03530_ ), .B2(_03455_ ), .ZN(_03689_ ) );
AND3_X1 _11380_ ( .A1(_03689_ ), .A2(_03441_ ), .A3(_03533_ ), .ZN(_03690_ ) );
OAI21_X1 _11381_ ( .A(_03445_ ), .B1(_03690_ ), .B2(_03538_ ), .ZN(_03691_ ) );
OR3_X1 _11382_ ( .A1(_03690_ ), .A2(_03538_ ), .A3(_03445_ ), .ZN(_03692_ ) );
NAND3_X1 _11383_ ( .A1(_03691_ ), .A2(_03630_ ), .A3(_03692_ ), .ZN(_03693_ ) );
AOI21_X1 _11384_ ( .A(\myifu.to_reset ), .B1(_03618_ ), .B2(\myexu.pc_jump [12] ), .ZN(_03694_ ) );
AOI211_X1 _11385_ ( .A(fanout_net_2 ), .B(_03685_ ), .C1(_03693_ ), .C2(_03694_ ), .ZN(_00256_ ) );
OR2_X1 _11386_ ( .A1(_03603_ ), .A2(_03604_ ), .ZN(_03695_ ) );
AND3_X1 _11387_ ( .A1(_03695_ ), .A2(_03628_ ), .A3(_03605_ ), .ZN(_03696_ ) );
AOI211_X1 _11388_ ( .A(\myifu.to_reset ), .B(_03696_ ), .C1(\myexu.pc_jump [29] ), .C2(_03618_ ), .ZN(_03697_ ) );
NOR2_X1 _11389_ ( .A1(_03612_ ), .A2(\mtvec [29] ), .ZN(_03698_ ) );
NOR3_X1 _11390_ ( .A1(_03697_ ), .A2(fanout_net_2 ), .A3(_03698_ ), .ZN(_00257_ ) );
AOI21_X1 _11391_ ( .A(_03441_ ), .B1(_03689_ ), .B2(_03533_ ), .ZN(_03699_ ) );
NOR3_X1 _11392_ ( .A1(_03690_ ), .A2(_03699_ ), .A3(_03617_ ), .ZN(_03700_ ) );
AOI211_X1 _11393_ ( .A(\myifu.to_reset ), .B(_03700_ ), .C1(\myexu.pc_jump [11] ), .C2(_03618_ ), .ZN(_03701_ ) );
NOR2_X1 _11394_ ( .A1(_03612_ ), .A2(\mtvec [11] ), .ZN(_03702_ ) );
NOR3_X1 _11395_ ( .A1(_03701_ ), .A2(fanout_net_2 ), .A3(_03702_ ), .ZN(_00258_ ) );
INV_X1 _11396_ ( .A(_03688_ ), .ZN(_03703_ ) );
OAI21_X1 _11397_ ( .A(_03628_ ), .B1(_03703_ ), .B2(_03456_ ), .ZN(_03704_ ) );
AOI21_X1 _11398_ ( .A(_03704_ ), .B1(_03703_ ), .B2(_03456_ ), .ZN(_03705_ ) );
AOI211_X1 _11399_ ( .A(\myifu.to_reset ), .B(_03705_ ), .C1(\myexu.pc_jump [10] ), .C2(_03617_ ), .ZN(_03706_ ) );
NOR2_X1 _11400_ ( .A1(_03612_ ), .A2(\mtvec [10] ), .ZN(_03707_ ) );
NOR3_X1 _11401_ ( .A1(_03706_ ), .A2(fanout_net_2 ), .A3(_03707_ ), .ZN(_00259_ ) );
AND3_X1 _11402_ ( .A1(_03526_ ), .A2(_03527_ ), .A3(_03686_ ), .ZN(_03708_ ) );
NOR3_X1 _11403_ ( .A1(_03708_ ), .A2(_03687_ ), .A3(_03212_ ), .ZN(_03709_ ) );
AOI211_X1 _11404_ ( .A(\myifu.to_reset ), .B(_03709_ ), .C1(\myexu.pc_jump [9] ), .C2(_03617_ ), .ZN(_03710_ ) );
NOR2_X1 _11405_ ( .A1(_03612_ ), .A2(\mtvec [9] ), .ZN(_03711_ ) );
NOR3_X1 _11406_ ( .A1(_03710_ ), .A2(fanout_net_2 ), .A3(_03711_ ), .ZN(_00260_ ) );
NOR2_X1 _11407_ ( .A1(_03520_ ), .A2(_03521_ ), .ZN(_03712_ ) );
XNOR2_X1 _11408_ ( .A(_03524_ ), .B(_01803_ ), .ZN(_03713_ ) );
OR2_X1 _11409_ ( .A1(_03712_ ), .A2(_03713_ ), .ZN(_03714_ ) );
AOI21_X1 _11410_ ( .A(_03212_ ), .B1(_03712_ ), .B2(_03713_ ), .ZN(_03715_ ) );
AOI221_X4 _11411_ ( .A(\myifu.to_reset ), .B1(\myexu.pc_jump [8] ), .B2(_03212_ ), .C1(_03714_ ), .C2(_03715_ ), .ZN(_03716_ ) );
NOR2_X1 _11412_ ( .A1(_03612_ ), .A2(\mtvec [8] ), .ZN(_03717_ ) );
NOR3_X1 _11413_ ( .A1(_03716_ ), .A2(fanout_net_2 ), .A3(_03717_ ), .ZN(_00261_ ) );
AOI21_X1 _11414_ ( .A(_03518_ ), .B1(_03514_ ), .B2(_03519_ ), .ZN(_03718_ ) );
NOR3_X1 _11415_ ( .A1(_03520_ ), .A2(_03718_ ), .A3(_03212_ ), .ZN(_03719_ ) );
AOI211_X1 _11416_ ( .A(\myifu.to_reset ), .B(_03719_ ), .C1(\myexu.pc_jump [7] ), .C2(_03617_ ), .ZN(_03720_ ) );
NOR2_X1 _11417_ ( .A1(_03612_ ), .A2(\mtvec [7] ), .ZN(_03721_ ) );
NOR3_X1 _11418_ ( .A1(_03720_ ), .A2(fanout_net_2 ), .A3(_03721_ ), .ZN(_00262_ ) );
NOR2_X1 _11419_ ( .A1(_03511_ ), .A2(_03513_ ), .ZN(_03722_ ) );
NOR2_X1 _11420_ ( .A1(_03482_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03723_ ) );
XNOR2_X1 _11421_ ( .A(_03477_ ), .B(_03478_ ), .ZN(_03724_ ) );
OR3_X1 _11422_ ( .A1(_03722_ ), .A2(_03723_ ), .A3(_03724_ ), .ZN(_03725_ ) );
OAI21_X1 _11423_ ( .A(_03724_ ), .B1(_03722_ ), .B2(_03723_ ), .ZN(_03726_ ) );
AOI21_X1 _11424_ ( .A(_03617_ ), .B1(_03725_ ), .B2(_03726_ ), .ZN(_03727_ ) );
AOI211_X1 _11425_ ( .A(\myifu.to_reset ), .B(_03727_ ), .C1(\myexu.pc_jump [6] ), .C2(_03617_ ), .ZN(_03728_ ) );
NOR2_X1 _11426_ ( .A1(_03612_ ), .A2(\mtvec [6] ), .ZN(_03729_ ) );
NOR3_X1 _11427_ ( .A1(_03728_ ), .A2(fanout_net_2 ), .A3(_03729_ ), .ZN(_00263_ ) );
AND2_X1 _11428_ ( .A1(_03511_ ), .A2(_03513_ ), .ZN(_03730_ ) );
NOR3_X1 _11429_ ( .A1(_03730_ ), .A2(_03722_ ), .A3(_03212_ ), .ZN(_03731_ ) );
AOI211_X1 _11430_ ( .A(\myifu.to_reset ), .B(_03731_ ), .C1(\myexu.pc_jump [5] ), .C2(_03617_ ), .ZN(_03732_ ) );
NOR2_X1 _11431_ ( .A1(_03614_ ), .A2(\mtvec [5] ), .ZN(_03733_ ) );
NOR3_X1 _11432_ ( .A1(_03732_ ), .A2(fanout_net_2 ), .A3(_03733_ ), .ZN(_00264_ ) );
NAND2_X1 _11433_ ( .A1(_03503_ ), .A2(_03504_ ), .ZN(_03734_ ) );
XNOR2_X1 _11434_ ( .A(_03508_ ), .B(_03505_ ), .ZN(_03735_ ) );
XOR2_X1 _11435_ ( .A(_03734_ ), .B(_03735_ ), .Z(_03736_ ) );
NAND2_X1 _11436_ ( .A1(_03736_ ), .A2(_03628_ ), .ZN(_03737_ ) );
OAI211_X1 _11437_ ( .A(_03737_ ), .B(_03426_ ), .C1(\myexu.pc_jump [4] ), .C2(_03628_ ), .ZN(_03738_ ) );
NAND2_X1 _11438_ ( .A1(\mtvec [4] ), .A2(\myifu.to_reset ), .ZN(_03739_ ) );
AOI21_X1 _11439_ ( .A(fanout_net_2 ), .B1(_03738_ ), .B2(_03739_ ), .ZN(_00265_ ) );
AND2_X1 _11440_ ( .A1(\mtvec [3] ), .A2(\myifu.to_reset ), .ZN(_03740_ ) );
XOR2_X1 _11441_ ( .A(_03496_ ), .B(_03502_ ), .Z(_03741_ ) );
MUX2_X1 _11442_ ( .A(\myexu.pc_jump [3] ), .B(_03741_ ), .S(_03628_ ), .Z(_03742_ ) );
AOI21_X1 _11443_ ( .A(_03740_ ), .B1(_03742_ ), .B2(_03612_ ), .ZN(_03743_ ) );
NOR2_X1 _11444_ ( .A1(_03743_ ), .A2(fanout_net_2 ), .ZN(_00266_ ) );
AND2_X1 _11445_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
NOR2_X1 _11446_ ( .A1(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A2(fanout_net_2 ), .ZN(_03744_ ) );
NOR2_X1 _11447_ ( .A1(_00265_ ), .A2(_03744_ ), .ZN(_03745_ ) );
BUF_X4 _11448_ ( .A(_03505_ ), .Z(_03746_ ) );
BUF_X4 _11449_ ( .A(_03746_ ), .Z(_03747_ ) );
BUF_X2 _11450_ ( .A(_03747_ ), .Z(_03748_ ) );
INV_X1 _11451_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_03749_ ) );
AOI21_X1 _11452_ ( .A(_03745_ ), .B1(_03748_ ), .B2(_03749_ ), .ZN(_00267_ ) );
NOR2_X1 _11453_ ( .A1(_03487_ ), .A2(_03493_ ), .ZN(_03750_ ) );
OAI22_X1 _11454_ ( .A1(_03494_ ), .A2(_03750_ ), .B1(_03211_ ), .B2(_03210_ ), .ZN(_03751_ ) );
OAI211_X1 _11455_ ( .A(_03751_ ), .B(_03614_ ), .C1(\myexu.pc_jump [2] ), .C2(_03630_ ), .ZN(_03752_ ) );
NAND2_X1 _11456_ ( .A1(\mtvec [2] ), .A2(\myifu.to_reset ), .ZN(_03753_ ) );
AOI21_X1 _11457_ ( .A(reset ), .B1(_03752_ ), .B2(_03753_ ), .ZN(_00268_ ) );
AOI211_X1 _11458_ ( .A(_03740_ ), .B(_03749_ ), .C1(_03742_ ), .C2(_03427_ ), .ZN(_03754_ ) );
BUF_X4 _11459_ ( .A(_03501_ ), .Z(_03755_ ) );
BUF_X2 _11460_ ( .A(_03755_ ), .Z(_03756_ ) );
AOI211_X1 _11461_ ( .A(reset ), .B(_03754_ ), .C1(_03756_ ), .C2(_03749_ ), .ZN(_00269_ ) );
OAI21_X1 _11462_ ( .A(_03595_ ), .B1(_03594_ ), .B2(_03601_ ), .ZN(_03757_ ) );
INV_X1 _11463_ ( .A(_03599_ ), .ZN(_03758_ ) );
AND2_X1 _11464_ ( .A1(_03757_ ), .A2(_03758_ ), .ZN(_03759_ ) );
XNOR2_X1 _11465_ ( .A(_03759_ ), .B(_03596_ ), .ZN(_03760_ ) );
MUX2_X1 _11466_ ( .A(\myexu.pc_jump [28] ), .B(_03760_ ), .S(_03628_ ), .Z(_03761_ ) );
MUX2_X1 _11467_ ( .A(\mtvec [28] ), .B(_03761_ ), .S(_03426_ ), .Z(_03762_ ) );
AND2_X1 _11468_ ( .A1(_03762_ ), .A2(_01570_ ), .ZN(_00270_ ) );
XNOR2_X1 _11469_ ( .A(_03491_ ), .B(_03492_ ), .ZN(_03763_ ) );
OAI21_X1 _11470_ ( .A(_03763_ ), .B1(_03210_ ), .B2(_03211_ ), .ZN(_03764_ ) );
OAI211_X1 _11471_ ( .A(_03764_ ), .B(_03614_ ), .C1(_03630_ ), .C2(\myexu.pc_jump [1] ), .ZN(_03765_ ) );
NAND2_X1 _11472_ ( .A1(\mtvec [1] ), .A2(\myifu.to_reset ), .ZN(_03766_ ) );
AOI21_X1 _11473_ ( .A(reset ), .B1(_03765_ ), .B2(_03766_ ), .ZN(_00271_ ) );
NOR2_X1 _11474_ ( .A1(_03594_ ), .A2(_03601_ ), .ZN(_03767_ ) );
XOR2_X1 _11475_ ( .A(_03767_ ), .B(_03595_ ), .Z(_03768_ ) );
NAND2_X1 _11476_ ( .A1(_03768_ ), .A2(_03629_ ), .ZN(_03769_ ) );
OAI211_X1 _11477_ ( .A(_03769_ ), .B(_03614_ ), .C1(\myexu.pc_jump [27] ), .C2(_03629_ ), .ZN(_03770_ ) );
NAND2_X1 _11478_ ( .A1(\mtvec [27] ), .A2(\myifu.to_reset ), .ZN(_03771_ ) );
AOI21_X1 _11479_ ( .A(reset ), .B1(_03770_ ), .B2(_03771_ ), .ZN(_00272_ ) );
OR3_X1 _11480_ ( .A1(_03210_ ), .A2(_03211_ ), .A3(\myexu.pc_jump [26] ), .ZN(_03772_ ) );
NAND2_X1 _11481_ ( .A1(_03591_ ), .A2(\IF_ID_pc [25] ), .ZN(_03773_ ) );
NAND2_X1 _11482_ ( .A1(_03590_ ), .A2(_03773_ ), .ZN(_03774_ ) );
XNOR2_X1 _11483_ ( .A(_03774_ ), .B(_03593_ ), .ZN(_03775_ ) );
OAI211_X1 _11484_ ( .A(_03614_ ), .B(_03772_ ), .C1(_03775_ ), .C2(_03618_ ), .ZN(_03776_ ) );
NAND2_X1 _11485_ ( .A1(\mtvec [26] ), .A2(\myifu.to_reset ), .ZN(_03777_ ) );
AOI21_X1 _11486_ ( .A(reset ), .B1(_03776_ ), .B2(_03777_ ), .ZN(_00273_ ) );
INV_X1 _11487_ ( .A(_03590_ ), .ZN(_03778_ ) );
NOR3_X1 _11488_ ( .A1(_03583_ ), .A2(_03589_ ), .A3(_03436_ ), .ZN(_03779_ ) );
OAI21_X1 _11489_ ( .A(_03629_ ), .B1(_03778_ ), .B2(_03779_ ), .ZN(_03780_ ) );
OAI211_X1 _11490_ ( .A(_03780_ ), .B(_03614_ ), .C1(\myexu.pc_jump [25] ), .C2(_03629_ ), .ZN(_03781_ ) );
NAND2_X1 _11491_ ( .A1(\mtvec [25] ), .A2(\myifu.to_reset ), .ZN(_03782_ ) );
AOI21_X1 _11492_ ( .A(reset ), .B1(_03781_ ), .B2(_03782_ ), .ZN(_00274_ ) );
OAI21_X1 _11493_ ( .A(_03582_ ), .B1(_03565_ ), .B2(_03575_ ), .ZN(_03783_ ) );
OAI21_X1 _11494_ ( .A(_03591_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_03784_ ) );
NAND2_X1 _11495_ ( .A1(_03783_ ), .A2(_03784_ ), .ZN(_03785_ ) );
NAND2_X1 _11496_ ( .A1(_03785_ ), .A2(_03578_ ), .ZN(_03786_ ) );
AND2_X1 _11497_ ( .A1(_03786_ ), .A2(_03588_ ), .ZN(_03787_ ) );
XNOR2_X1 _11498_ ( .A(_03787_ ), .B(_03577_ ), .ZN(_03788_ ) );
MUX2_X1 _11499_ ( .A(\myexu.pc_jump [24] ), .B(_03788_ ), .S(_03628_ ), .Z(_03789_ ) );
MUX2_X1 _11500_ ( .A(\mtvec [24] ), .B(_03789_ ), .S(_03426_ ), .Z(_03790_ ) );
AND2_X1 _11501_ ( .A1(_03790_ ), .A2(_01570_ ), .ZN(_00275_ ) );
XNOR2_X1 _11502_ ( .A(_03785_ ), .B(_03578_ ), .ZN(_03791_ ) );
NAND2_X1 _11503_ ( .A1(_03791_ ), .A2(_03629_ ), .ZN(_03792_ ) );
OAI211_X1 _11504_ ( .A(_03792_ ), .B(_03427_ ), .C1(\myexu.pc_jump [23] ), .C2(_03629_ ), .ZN(_03793_ ) );
NAND2_X1 _11505_ ( .A1(\mtvec [23] ), .A2(\myifu.to_reset ), .ZN(_03794_ ) );
AOI21_X1 _11506_ ( .A(reset ), .B1(_03793_ ), .B2(_03794_ ), .ZN(_00276_ ) );
INV_X1 _11507_ ( .A(_03576_ ), .ZN(_03795_ ) );
NOR2_X1 _11508_ ( .A1(_03795_ ), .A2(_03580_ ), .ZN(_03796_ ) );
NOR2_X1 _11509_ ( .A1(_03796_ ), .A2(_03585_ ), .ZN(_03797_ ) );
XOR2_X1 _11510_ ( .A(_03797_ ), .B(_03581_ ), .Z(_03798_ ) );
MUX2_X1 _11511_ ( .A(\myexu.pc_jump [22] ), .B(_03798_ ), .S(_03627_ ), .Z(_03799_ ) );
MUX2_X1 _11512_ ( .A(\mtvec [22] ), .B(_03799_ ), .S(_03426_ ), .Z(_03800_ ) );
AND2_X1 _11513_ ( .A1(_03800_ ), .A2(_01570_ ), .ZN(_00277_ ) );
NAND2_X1 _11514_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_03801_ ) );
AND2_X1 _11515_ ( .A1(_03591_ ), .A2(\IF_ID_pc [30] ), .ZN(_03802_ ) );
INV_X1 _11516_ ( .A(_03802_ ), .ZN(_03803_ ) );
OAI21_X1 _11517_ ( .A(_01866_ ), .B1(_03432_ ), .B2(_03433_ ), .ZN(_03804_ ) );
NAND4_X1 _11518_ ( .A1(_03603_ ), .A2(_03604_ ), .A3(_03803_ ), .A4(_03804_ ), .ZN(_03805_ ) );
NAND3_X1 _11519_ ( .A1(_03591_ ), .A2(_01866_ ), .A3(\IF_ID_pc [29] ), .ZN(_03806_ ) );
AND3_X1 _11520_ ( .A1(_03805_ ), .A2(_03803_ ), .A3(_03806_ ), .ZN(_03807_ ) );
XNOR2_X1 _11521_ ( .A(_03591_ ), .B(_01837_ ), .ZN(_03808_ ) );
OR2_X1 _11522_ ( .A1(_03807_ ), .A2(_03808_ ), .ZN(_03809_ ) );
AOI21_X1 _11523_ ( .A(_03617_ ), .B1(_03807_ ), .B2(_03808_ ), .ZN(_03810_ ) );
AND2_X1 _11524_ ( .A1(_03809_ ), .A2(_03810_ ), .ZN(_03811_ ) );
OAI21_X1 _11525_ ( .A(_03427_ ), .B1(_03630_ ), .B2(\myexu.pc_jump [31] ), .ZN(_03812_ ) );
OAI211_X1 _11526_ ( .A(_01570_ ), .B(_03801_ ), .C1(_03811_ ), .C2(_03812_ ), .ZN(_00278_ ) );
NOR2_X1 _11527_ ( .A1(_01986_ ), .A2(_02022_ ), .ZN(_03813_ ) );
INV_X1 _11528_ ( .A(_03813_ ), .ZN(_03814_ ) );
NOR2_X1 _11529_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_03815_ ) );
NOR2_X1 _11530_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_03816_ ) );
INV_X1 _11531_ ( .A(\io_master_rid [1] ), .ZN(_03817_ ) );
NAND4_X1 _11532_ ( .A1(_03815_ ), .A2(_03816_ ), .A3(_03817_ ), .A4(\io_master_rid [0] ), .ZN(_03818_ ) );
AOI21_X1 _11533_ ( .A(_01954_ ), .B1(_03814_ ), .B2(_03818_ ), .ZN(_03819_ ) );
NOR2_X1 _11534_ ( .A1(_02072_ ), .A2(io_master_rlast ), .ZN(_03820_ ) );
INV_X1 _11535_ ( .A(_03820_ ), .ZN(_03821_ ) );
INV_X1 _11536_ ( .A(_01999_ ), .ZN(\io_master_araddr [21] ) );
INV_X1 _11537_ ( .A(_02016_ ), .ZN(\io_master_araddr [22] ) );
NOR4_X4 _11538_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [22] ), .A3(\io_master_araddr [23] ), .A4(\io_master_araddr [20] ), .ZN(_03822_ ) );
INV_X1 _11539_ ( .A(_02003_ ), .ZN(\io_master_araddr [19] ) );
INV_X2 _11540_ ( .A(_02020_ ), .ZN(\io_master_araddr [16] ) );
NOR4_X4 _11541_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [16] ), .A3(\io_master_araddr [17] ), .A4(\io_master_araddr [18] ), .ZN(_03823_ ) );
AND2_X4 _11542_ ( .A1(_03822_ ), .A2(_03823_ ), .ZN(_03824_ ) );
NAND4_X2 _11543_ ( .A1(\io_master_araddr [25] ), .A2(_01979_ ), .A3(_01995_ ), .A4(_02012_ ), .ZN(_03825_ ) );
NAND4_X2 _11544_ ( .A1(_01970_ ), .A2(_01974_ ), .A3(_01991_ ), .A4(_02008_ ), .ZN(_03826_ ) );
NOR2_X2 _11545_ ( .A1(_03825_ ), .A2(_03826_ ), .ZN(_03827_ ) );
AOI21_X1 _11546_ ( .A(io_master_rvalid ), .B1(_03824_ ), .B2(_03827_ ), .ZN(_03828_ ) );
AND4_X1 _11547_ ( .A1(\myclint.state_r_$_NOT__A_Y ), .A2(_03822_ ), .A3(_03823_ ), .A4(_03827_ ), .ZN(_03829_ ) );
NOR2_X1 _11548_ ( .A1(_03828_ ), .A2(_03829_ ), .ZN(_03830_ ) );
NAND3_X1 _11549_ ( .A1(_03819_ ), .A2(_03821_ ), .A3(_03830_ ), .ZN(_03831_ ) );
INV_X1 _11550_ ( .A(\myifu.tmp_offset [2] ), .ZN(_03832_ ) );
AND3_X1 _11551_ ( .A1(_03831_ ), .A2(_01536_ ), .A3(_03832_ ), .ZN(_00279_ ) );
NOR3_X1 _11552_ ( .A1(reset ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00280_ ) );
AND3_X1 _11553_ ( .A1(_02092_ ), .A2(_03213_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_03833_ ) );
INV_X1 _11554_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_03834_ ) );
MUX2_X1 _11555_ ( .A(_02092_ ), .B(_03834_ ), .S(\myifu.to_reset ), .Z(_03835_ ) );
AOI211_X1 _11556_ ( .A(reset ), .B(_03833_ ), .C1(_03835_ ), .C2(\myifu.state [1] ), .ZN(_00281_ ) );
INV_X1 _11557_ ( .A(_02051_ ), .ZN(_03836_ ) );
NOR2_X2 _11558_ ( .A1(_02059_ ), .A2(_03836_ ), .ZN(_03837_ ) );
INV_X2 _11559_ ( .A(_03837_ ), .ZN(_03838_ ) );
BUF_X2 _11560_ ( .A(_03838_ ), .Z(_03839_ ) );
BUF_X4 _11561_ ( .A(_02128_ ), .Z(_03840_ ) );
BUF_X4 _11562_ ( .A(_03840_ ), .Z(_03841_ ) );
MUX2_X1 _11563_ ( .A(\LS_WB_waddr_csreg [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_03841_ ), .Z(_03842_ ) );
NOR2_X1 _11564_ ( .A1(\EX_LS_flag [2] ), .A2(\EX_LS_flag [1] ), .ZN(_03843_ ) );
NOR2_X1 _11565_ ( .A1(_02050_ ), .A2(_03843_ ), .ZN(_03844_ ) );
NOR2_X1 _11566_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_03845_ ) );
AND2_X2 _11567_ ( .A1(_03845_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_03846_ ) );
NOR2_X1 _11568_ ( .A1(_03844_ ), .A2(_03846_ ), .ZN(_03847_ ) );
BUF_X4 _11569_ ( .A(_03847_ ), .Z(_03848_ ) );
BUF_X2 _11570_ ( .A(_03848_ ), .Z(_03849_ ) );
AND3_X1 _11571_ ( .A1(_03839_ ), .A2(_03842_ ), .A3(_03849_ ), .ZN(_00284_ ) );
NOR2_X1 _11572_ ( .A1(_03837_ ), .A2(_03846_ ), .ZN(_03850_ ) );
AND2_X1 _11573_ ( .A1(_03850_ ), .A2(_02040_ ), .ZN(_03851_ ) );
INV_X1 _11574_ ( .A(_03851_ ), .ZN(_03852_ ) );
BUF_X2 _11575_ ( .A(_02050_ ), .Z(_03853_ ) );
NAND3_X1 _11576_ ( .A1(_03853_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_03854_ ) );
BUF_X4 _11577_ ( .A(_01941_ ), .Z(_03855_ ) );
NAND2_X1 _11578_ ( .A1(_03855_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03856_ ) );
AOI21_X1 _11579_ ( .A(_03852_ ), .B1(_03854_ ), .B2(_03856_ ), .ZN(_00285_ ) );
NAND3_X1 _11580_ ( .A1(_03853_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_03857_ ) );
NAND2_X1 _11581_ ( .A1(_03855_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_03858_ ) );
AOI21_X1 _11582_ ( .A(_03852_ ), .B1(_03857_ ), .B2(_03858_ ), .ZN(_00286_ ) );
NAND3_X1 _11583_ ( .A1(_03853_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_03859_ ) );
NAND2_X1 _11584_ ( .A1(_03855_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_03860_ ) );
AOI21_X1 _11585_ ( .A(_03852_ ), .B1(_03859_ ), .B2(_03860_ ), .ZN(_00287_ ) );
NAND3_X1 _11586_ ( .A1(_03853_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_03861_ ) );
NAND2_X1 _11587_ ( .A1(_03855_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03862_ ) );
AOI21_X1 _11588_ ( .A(_03852_ ), .B1(_03861_ ), .B2(_03862_ ), .ZN(_00288_ ) );
NAND3_X1 _11589_ ( .A1(_03853_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_03863_ ) );
NAND2_X1 _11590_ ( .A1(_03855_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_03864_ ) );
AOI21_X1 _11591_ ( .A(_03852_ ), .B1(_03863_ ), .B2(_03864_ ), .ZN(_00289_ ) );
NAND3_X1 _11592_ ( .A1(_03853_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_03865_ ) );
NAND2_X1 _11593_ ( .A1(_03855_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_03866_ ) );
AOI21_X1 _11594_ ( .A(_03852_ ), .B1(_03865_ ), .B2(_03866_ ), .ZN(_00290_ ) );
NAND3_X1 _11595_ ( .A1(_03853_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_flag [2] ), .ZN(_03867_ ) );
NAND2_X1 _11596_ ( .A1(_03855_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_03868_ ) );
AOI21_X1 _11597_ ( .A(_03852_ ), .B1(_03867_ ), .B2(_03868_ ), .ZN(_00291_ ) );
INV_X1 _11598_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_03869_ ) );
INV_X1 _11599_ ( .A(\EX_LS_flag [0] ), .ZN(_03870_ ) );
AND4_X1 _11600_ ( .A1(_03869_ ), .A2(_03870_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03871_ ) );
NOR2_X1 _11601_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_03872_ ) );
OAI211_X1 _11602_ ( .A(_03850_ ), .B(_02040_ ), .C1(_03871_ ), .C2(_03872_ ), .ZN(_00292_ ) );
INV_X1 _11603_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_03873_ ) );
AND4_X1 _11604_ ( .A1(_03873_ ), .A2(_03870_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03874_ ) );
NOR2_X1 _11605_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_03875_ ) );
OAI211_X1 _11606_ ( .A(_03850_ ), .B(_02040_ ), .C1(_03874_ ), .C2(_03875_ ), .ZN(_00293_ ) );
INV_X1 _11607_ ( .A(\EX_LS_dest_csreg_mem [6] ), .ZN(_03876_ ) );
AND4_X1 _11608_ ( .A1(_03876_ ), .A2(_03870_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03877_ ) );
NOR2_X1 _11609_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_03878_ ) );
OAI211_X1 _11610_ ( .A(_03850_ ), .B(_02040_ ), .C1(_03877_ ), .C2(_03878_ ), .ZN(_00294_ ) );
INV_X1 _11611_ ( .A(fanout_net_3 ), .ZN(_03879_ ) );
AND4_X1 _11612_ ( .A1(_03879_ ), .A2(_03870_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03880_ ) );
NOR2_X1 _11613_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_03881_ ) );
OAI211_X1 _11614_ ( .A(_03850_ ), .B(_02040_ ), .C1(_03880_ ), .C2(_03881_ ), .ZN(_00295_ ) );
INV_X1 _11615_ ( .A(\mysc.state [2] ), .ZN(_03882_ ) );
NOR2_X1 _11616_ ( .A1(_03882_ ), .A2(reset ), .ZN(_00303_ ) );
NOR2_X1 _11617_ ( .A1(_03331_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _11618_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_03883_ ) );
NOR2_X1 _11619_ ( .A1(_03343_ ), .A2(\ID_EX_typ [6] ), .ZN(_03884_ ) );
AND2_X2 _11620_ ( .A1(_03884_ ), .A2(\ID_EX_typ [5] ), .ZN(_03885_ ) );
INV_X1 _11621_ ( .A(fanout_net_4 ), .ZN(_03886_ ) );
AND2_X2 _11622_ ( .A1(_03885_ ), .A2(_03886_ ), .ZN(_03887_ ) );
INV_X1 _11623_ ( .A(_03887_ ), .ZN(_03888_ ) );
INV_X1 _11624_ ( .A(\ID_EX_typ [5] ), .ZN(_03889_ ) );
INV_X1 _11625_ ( .A(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_03890_ ) );
NAND3_X1 _11626_ ( .A1(_03884_ ), .A2(_03889_ ), .A3(_03890_ ), .ZN(_03891_ ) );
AOI21_X1 _11627_ ( .A(_03883_ ), .B1(_03888_ ), .B2(_03891_ ), .ZN(_03892_ ) );
INV_X1 _11628_ ( .A(\myec.state [1] ), .ZN(_03893_ ) );
NAND2_X1 _11629_ ( .A1(_03893_ ), .A2(\myec.state [0] ), .ZN(_03894_ ) );
NOR2_X1 _11630_ ( .A1(reset ), .A2(excp_written ), .ZN(_03895_ ) );
AND2_X1 _11631_ ( .A1(_03894_ ), .A2(_03895_ ), .ZN(_03896_ ) );
BUF_X4 _11632_ ( .A(_03896_ ), .Z(_03897_ ) );
INV_X1 _11633_ ( .A(\ID_EX_typ [6] ), .ZN(_03898_ ) );
INV_X1 _11634_ ( .A(EXU_valid_LSU ), .ZN(_03899_ ) );
AND4_X1 _11635_ ( .A1(\ID_EX_typ [7] ), .A2(_03898_ ), .A3(_03899_ ), .A4(IDU_valid_EXU ), .ZN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _11636_ ( .A1(_03211_ ), .A2(check_assert ), .ZN(_03900_ ) );
OAI21_X1 _11637_ ( .A(_03897_ ), .B1(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(_03900_ ), .ZN(_03901_ ) );
NOR2_X1 _11638_ ( .A1(_03892_ ), .A2(_03901_ ), .ZN(_00096_ ) );
CLKBUF_X2 _11639_ ( .A(_03894_ ), .Z(_03902_ ) );
CLKBUF_X2 _11640_ ( .A(_03902_ ), .Z(_03903_ ) );
CLKBUF_X2 _11641_ ( .A(_03895_ ), .Z(_03904_ ) );
CLKBUF_X2 _11642_ ( .A(_03904_ ), .Z(_03905_ ) );
AND3_X1 _11643_ ( .A1(_03903_ ), .A2(\ID_EX_rd [4] ), .A3(_03905_ ), .ZN(_00117_ ) );
AND3_X1 _11644_ ( .A1(_03903_ ), .A2(\ID_EX_rd [3] ), .A3(_03905_ ), .ZN(_00118_ ) );
AND3_X1 _11645_ ( .A1(_03903_ ), .A2(\ID_EX_rd [2] ), .A3(_03905_ ), .ZN(_00119_ ) );
AND3_X1 _11646_ ( .A1(_03903_ ), .A2(\ID_EX_rd [1] ), .A3(_03905_ ), .ZN(_00120_ ) );
AND3_X1 _11647_ ( .A1(_03903_ ), .A2(\ID_EX_rd [0] ), .A3(_03905_ ), .ZN(_00121_ ) );
INV_X2 _11648_ ( .A(_03897_ ), .ZN(_03906_ ) );
BUF_X4 _11649_ ( .A(_03906_ ), .Z(_03907_ ) );
AND2_X1 _11650_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_03908_ ) );
AND2_X1 _11651_ ( .A1(_03908_ ), .A2(\ID_EX_pc [4] ), .ZN(_03909_ ) );
AND2_X1 _11652_ ( .A1(_03909_ ), .A2(\ID_EX_pc [5] ), .ZN(_03910_ ) );
AND2_X1 _11653_ ( .A1(_03910_ ), .A2(\ID_EX_pc [6] ), .ZN(_03911_ ) );
AND2_X1 _11654_ ( .A1(_03911_ ), .A2(\ID_EX_pc [7] ), .ZN(_03912_ ) );
AND2_X1 _11655_ ( .A1(_03912_ ), .A2(\ID_EX_pc [8] ), .ZN(_03913_ ) );
AND2_X2 _11656_ ( .A1(_03913_ ), .A2(\ID_EX_pc [9] ), .ZN(_03914_ ) );
AND2_X1 _11657_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_03915_ ) );
AND2_X1 _11658_ ( .A1(_03914_ ), .A2(_03915_ ), .ZN(_03916_ ) );
AND3_X1 _11659_ ( .A1(_03916_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_03917_ ) );
AND3_X1 _11660_ ( .A1(_03917_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_03918_ ) );
AND3_X1 _11661_ ( .A1(_03918_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_03919_ ) );
AND3_X1 _11662_ ( .A1(_03919_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_03920_ ) );
AND3_X1 _11663_ ( .A1(_03920_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_03921_ ) );
AND3_X1 _11664_ ( .A1(_03921_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_03922_ ) );
AND3_X1 _11665_ ( .A1(_03922_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_03923_ ) );
AND3_X1 _11666_ ( .A1(_03923_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_03924_ ) );
NAND3_X1 _11667_ ( .A1(_03924_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_03925_ ) );
XNOR2_X1 _11668_ ( .A(_03925_ ), .B(\ID_EX_pc [30] ), .ZN(_03926_ ) );
XOR2_X1 _11669_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_03927_ ) );
XOR2_X1 _11670_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_03928_ ) );
XOR2_X1 _11671_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_03929_ ) );
XOR2_X1 _11672_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_03930_ ) );
AND2_X1 _11673_ ( .A1(_03929_ ), .A2(_03930_ ), .ZN(_03931_ ) );
XOR2_X1 _11674_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_03932_ ) );
XOR2_X1 _11675_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_03933_ ) );
AND2_X1 _11676_ ( .A1(_03932_ ), .A2(_03933_ ), .ZN(_03934_ ) );
AND2_X1 _11677_ ( .A1(_03931_ ), .A2(_03934_ ), .ZN(_03935_ ) );
XOR2_X1 _11678_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_03936_ ) );
XOR2_X1 _11679_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_03937_ ) );
AND2_X1 _11680_ ( .A1(_03936_ ), .A2(_03937_ ), .ZN(_03938_ ) );
XOR2_X1 _11681_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_03939_ ) );
XOR2_X1 _11682_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_03940_ ) );
AND3_X1 _11683_ ( .A1(_03938_ ), .A2(_03939_ ), .A3(_03940_ ), .ZN(_03941_ ) );
XOR2_X1 _11684_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_03942_ ) );
XOR2_X1 _11685_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_03943_ ) );
AND2_X1 _11686_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_03944_ ) );
AND2_X1 _11687_ ( .A1(_03943_ ), .A2(_03944_ ), .ZN(_03945_ ) );
AND2_X1 _11688_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_03946_ ) );
OAI21_X1 _11689_ ( .A(_03942_ ), .B1(_03945_ ), .B2(_03946_ ), .ZN(_03947_ ) );
INV_X1 _11690_ ( .A(_03947_ ), .ZN(_03948_ ) );
AND2_X1 _11691_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_03949_ ) );
NOR2_X1 _11692_ ( .A1(_03948_ ), .A2(_03949_ ), .ZN(_03950_ ) );
NOR2_X1 _11693_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03951_ ) );
NOR2_X1 _11694_ ( .A1(_03950_ ), .A2(_03951_ ), .ZN(_03952_ ) );
AND2_X1 _11695_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03953_ ) );
NOR2_X1 _11696_ ( .A1(_03952_ ), .A2(_03953_ ), .ZN(_03954_ ) );
AND2_X1 _11697_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03955_ ) );
NOR2_X1 _11698_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03956_ ) );
NOR3_X1 _11699_ ( .A1(_03954_ ), .A2(_03955_ ), .A3(_03956_ ), .ZN(_03957_ ) );
NOR2_X1 _11700_ ( .A1(_03957_ ), .A2(_03955_ ), .ZN(_03958_ ) );
NOR2_X1 _11701_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03959_ ) );
NOR2_X1 _11702_ ( .A1(_03958_ ), .A2(_03959_ ), .ZN(_03960_ ) );
AND2_X1 _11703_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03961_ ) );
NOR2_X1 _11704_ ( .A1(_03960_ ), .A2(_03961_ ), .ZN(_03962_ ) );
AND2_X1 _11705_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03963_ ) );
NOR2_X1 _11706_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03964_ ) );
NOR3_X1 _11707_ ( .A1(_03962_ ), .A2(_03963_ ), .A3(_03964_ ), .ZN(_03965_ ) );
NOR2_X1 _11708_ ( .A1(_03965_ ), .A2(_03963_ ), .ZN(_03966_ ) );
NOR2_X1 _11709_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03967_ ) );
NOR2_X1 _11710_ ( .A1(_03966_ ), .A2(_03967_ ), .ZN(_03968_ ) );
AND2_X1 _11711_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03969_ ) );
NOR2_X1 _11712_ ( .A1(_03968_ ), .A2(_03969_ ), .ZN(_03970_ ) );
INV_X1 _11713_ ( .A(_03970_ ), .ZN(_03971_ ) );
XOR2_X1 _11714_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_03972_ ) );
XOR2_X1 _11715_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_03973_ ) );
AND2_X1 _11716_ ( .A1(_03972_ ), .A2(_03973_ ), .ZN(_03974_ ) );
XOR2_X1 _11717_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_03975_ ) );
XOR2_X1 _11718_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .Z(_03976_ ) );
AND2_X1 _11719_ ( .A1(_03975_ ), .A2(_03976_ ), .ZN(_03977_ ) );
AND2_X1 _11720_ ( .A1(_03974_ ), .A2(_03977_ ), .ZN(_03978_ ) );
XOR2_X1 _11721_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_03979_ ) );
XOR2_X1 _11722_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_03980_ ) );
AND2_X1 _11723_ ( .A1(_03979_ ), .A2(_03980_ ), .ZN(_03981_ ) );
XOR2_X1 _11724_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_03982_ ) );
XOR2_X1 _11725_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_03983_ ) );
AND2_X1 _11726_ ( .A1(_03982_ ), .A2(_03983_ ), .ZN(_03984_ ) );
AND2_X1 _11727_ ( .A1(_03981_ ), .A2(_03984_ ), .ZN(_03985_ ) );
AND3_X1 _11728_ ( .A1(_03971_ ), .A2(_03978_ ), .A3(_03985_ ), .ZN(_03986_ ) );
AND2_X1 _11729_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_03987_ ) );
AND2_X1 _11730_ ( .A1(_03979_ ), .A2(_03987_ ), .ZN(_03988_ ) );
AOI21_X1 _11731_ ( .A(_03988_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_03989_ ) );
AND2_X1 _11732_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_03990_ ) );
AND2_X1 _11733_ ( .A1(_03983_ ), .A2(_03990_ ), .ZN(_03991_ ) );
AOI21_X1 _11734_ ( .A(_03991_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_03992_ ) );
INV_X1 _11735_ ( .A(_03981_ ), .ZN(_03993_ ) );
OAI21_X1 _11736_ ( .A(_03989_ ), .B1(_03992_ ), .B2(_03993_ ), .ZN(_03994_ ) );
NAND2_X1 _11737_ ( .A1(_03994_ ), .A2(_03978_ ), .ZN(_03995_ ) );
AND2_X1 _11738_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_imm [13] ), .ZN(_03996_ ) );
AND2_X1 _11739_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_03997_ ) );
AOI21_X1 _11740_ ( .A(_03996_ ), .B1(_03976_ ), .B2(_03997_ ), .ZN(_03998_ ) );
INV_X1 _11741_ ( .A(_03998_ ), .ZN(_03999_ ) );
NAND2_X1 _11742_ ( .A1(_03999_ ), .A2(_03974_ ), .ZN(_04000_ ) );
AND2_X1 _11743_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04001_ ) );
AND2_X1 _11744_ ( .A1(_03972_ ), .A2(_04001_ ), .ZN(_04002_ ) );
AOI21_X1 _11745_ ( .A(_04002_ ), .B1(\ID_EX_pc [15] ), .B2(\ID_EX_imm [15] ), .ZN(_04003_ ) );
AND3_X1 _11746_ ( .A1(_03995_ ), .A2(_04000_ ), .A3(_04003_ ), .ZN(_04004_ ) );
INV_X1 _11747_ ( .A(_04004_ ), .ZN(_04005_ ) );
OAI211_X1 _11748_ ( .A(_03935_ ), .B(_03941_ ), .C1(_03986_ ), .C2(_04005_ ), .ZN(_04006_ ) );
NAND3_X1 _11749_ ( .A1(_03929_ ), .A2(\ID_EX_pc [22] ), .A3(\ID_EX_imm [22] ), .ZN(_04007_ ) );
INV_X1 _11750_ ( .A(\ID_EX_pc [23] ), .ZN(_04008_ ) );
NAND3_X1 _11751_ ( .A1(_03936_ ), .A2(\ID_EX_pc [18] ), .A3(\ID_EX_imm [18] ), .ZN(_04009_ ) );
INV_X1 _11752_ ( .A(\ID_EX_pc [19] ), .ZN(_04010_ ) );
OAI21_X1 _11753_ ( .A(_04009_ ), .B1(_04010_ ), .B2(_02430_ ), .ZN(_04011_ ) );
AND2_X1 _11754_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_04012_ ) );
AND2_X1 _11755_ ( .A1(_03939_ ), .A2(_04012_ ), .ZN(_04013_ ) );
AOI21_X1 _11756_ ( .A(_04013_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_04014_ ) );
INV_X1 _11757_ ( .A(_04014_ ), .ZN(_04015_ ) );
AOI21_X1 _11758_ ( .A(_04011_ ), .B1(_04015_ ), .B2(_03938_ ), .ZN(_04016_ ) );
INV_X1 _11759_ ( .A(_03935_ ), .ZN(_04017_ ) );
OAI221_X1 _11760_ ( .A(_04007_ ), .B1(_04008_ ), .B2(_02308_ ), .C1(_04016_ ), .C2(_04017_ ), .ZN(_04018_ ) );
AND2_X1 _11761_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_04019_ ) );
AND2_X1 _11762_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_04020_ ) );
AOI21_X1 _11763_ ( .A(_04019_ ), .B1(_03933_ ), .B2(_04020_ ), .ZN(_04021_ ) );
INV_X1 _11764_ ( .A(_04021_ ), .ZN(_04022_ ) );
AOI21_X1 _11765_ ( .A(_04018_ ), .B1(_03931_ ), .B2(_04022_ ), .ZN(_04023_ ) );
NAND2_X1 _11766_ ( .A1(_04006_ ), .A2(_04023_ ), .ZN(_04024_ ) );
XOR2_X1 _11767_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_04025_ ) );
NAND2_X1 _11768_ ( .A1(_04024_ ), .A2(_04025_ ), .ZN(_04026_ ) );
NAND2_X1 _11769_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_04027_ ) );
INV_X1 _11770_ ( .A(\ID_EX_pc [25] ), .ZN(_04028_ ) );
AOI22_X1 _11771_ ( .A1(_04026_ ), .A2(_04027_ ), .B1(_04028_ ), .B2(_02968_ ), .ZN(_04029_ ) );
AND2_X1 _11772_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_04030_ ) );
OAI211_X1 _11773_ ( .A(_03927_ ), .B(_03928_ ), .C1(_04029_ ), .C2(_04030_ ), .ZN(_04031_ ) );
AND2_X1 _11774_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_04032_ ) );
AND2_X1 _11775_ ( .A1(_03927_ ), .A2(_04032_ ), .ZN(_04033_ ) );
AOI21_X1 _11776_ ( .A(_04033_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_04034_ ) );
NAND2_X1 _11777_ ( .A1(_04031_ ), .A2(_04034_ ), .ZN(_04035_ ) );
XOR2_X1 _11778_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_04036_ ) );
NAND2_X1 _11779_ ( .A1(_04035_ ), .A2(_04036_ ), .ZN(_04037_ ) );
NAND2_X1 _11780_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_04038_ ) );
INV_X1 _11781_ ( .A(\ID_EX_pc [29] ), .ZN(_04039_ ) );
AOI22_X1 _11782_ ( .A1(_04037_ ), .A2(_04038_ ), .B1(_04039_ ), .B2(_02200_ ), .ZN(_04040_ ) );
AND2_X1 _11783_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_04041_ ) );
OR2_X1 _11784_ ( .A1(_04040_ ), .A2(_04041_ ), .ZN(_04042_ ) );
XOR2_X1 _11785_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_04043_ ) );
XOR2_X1 _11786_ ( .A(_04042_ ), .B(_04043_ ), .Z(_04044_ ) );
NOR2_X1 _11787_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_4 ), .ZN(_04045_ ) );
AND2_X1 _11788_ ( .A1(_04045_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04046_ ) );
INV_X1 _11789_ ( .A(fanout_net_39 ), .ZN(_04047_ ) );
BUF_X4 _11790_ ( .A(_04047_ ), .Z(_04048_ ) );
BUF_X4 _11791_ ( .A(_04048_ ), .Z(_04049_ ) );
BUF_X4 _11792_ ( .A(_04049_ ), .Z(_04050_ ) );
INV_X1 _11793_ ( .A(fanout_net_27 ), .ZN(_04051_ ) );
CLKBUF_X2 _11794_ ( .A(_04051_ ), .Z(_04052_ ) );
CLKBUF_X2 _11795_ ( .A(_04052_ ), .Z(_04053_ ) );
BUF_X2 _11796_ ( .A(_04053_ ), .Z(_04054_ ) );
BUF_X2 _11797_ ( .A(_04054_ ), .Z(_04055_ ) );
OR2_X1 _11798_ ( .A1(_04055_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04056_ ) );
OAI211_X1 _11799_ ( .A(_04056_ ), .B(fanout_net_36 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04057_ ) );
INV_X1 _11800_ ( .A(fanout_net_38 ), .ZN(_04058_ ) );
BUF_X4 _11801_ ( .A(_04058_ ), .Z(_04059_ ) );
BUF_X4 _11802_ ( .A(_04059_ ), .Z(_04060_ ) );
BUF_X4 _11803_ ( .A(_04060_ ), .Z(_04061_ ) );
NAND2_X1 _11804_ ( .A1(_02154_ ), .A2(fanout_net_27 ), .ZN(_04062_ ) );
INV_X2 _11805_ ( .A(fanout_net_36 ), .ZN(_04063_ ) );
BUF_X4 _11806_ ( .A(_04063_ ), .Z(_04064_ ) );
BUF_X4 _11807_ ( .A(_04064_ ), .Z(_04065_ ) );
BUF_X4 _11808_ ( .A(_04065_ ), .Z(_04066_ ) );
BUF_X4 _11809_ ( .A(_04066_ ), .Z(_04067_ ) );
OAI211_X1 _11810_ ( .A(_04062_ ), .B(_04067_ ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04068_ ) );
NAND3_X1 _11811_ ( .A1(_04057_ ), .A2(_04061_ ), .A3(_04068_ ), .ZN(_04069_ ) );
MUX2_X1 _11812_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04070_ ) );
MUX2_X1 _11813_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04071_ ) );
MUX2_X1 _11814_ ( .A(_04070_ ), .B(_04071_ ), .S(_04067_ ), .Z(_04072_ ) );
BUF_X4 _11815_ ( .A(_04061_ ), .Z(_04073_ ) );
OAI211_X1 _11816_ ( .A(_04050_ ), .B(_04069_ ), .C1(_04072_ ), .C2(_04073_ ), .ZN(_04074_ ) );
OR2_X1 _11817_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04075_ ) );
BUF_X2 _11818_ ( .A(_04055_ ), .Z(_04076_ ) );
OAI211_X1 _11819_ ( .A(_04075_ ), .B(fanout_net_36 ), .C1(_04076_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04077_ ) );
OR2_X1 _11820_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04078_ ) );
OAI211_X1 _11821_ ( .A(_04078_ ), .B(_04067_ ), .C1(_04076_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04079_ ) );
NAND3_X1 _11822_ ( .A1(_04077_ ), .A2(_04079_ ), .A3(fanout_net_38 ), .ZN(_04080_ ) );
MUX2_X1 _11823_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04081_ ) );
MUX2_X1 _11824_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04082_ ) );
MUX2_X1 _11825_ ( .A(_04081_ ), .B(_04082_ ), .S(fanout_net_36 ), .Z(_04083_ ) );
OAI211_X1 _11826_ ( .A(fanout_net_39 ), .B(_04080_ ), .C1(_04083_ ), .C2(fanout_net_38 ), .ZN(_04084_ ) );
NAND2_X1 _11827_ ( .A1(_04074_ ), .A2(_04084_ ), .ZN(_04085_ ) );
XNOR2_X1 _11828_ ( .A(\EX_LS_dest_reg [3] ), .B(\ID_EX_rs2 [3] ), .ZN(_04086_ ) );
XNOR2_X1 _11829_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_04087_ ) );
XNOR2_X1 _11830_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_04088_ ) );
XNOR2_X1 _11831_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_04089_ ) );
AND4_X1 _11832_ ( .A1(_04086_ ), .A2(_04087_ ), .A3(_04088_ ), .A4(_04089_ ), .ZN(_04090_ ) );
OAI21_X1 _11833_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02133_ ), .B2(\ID_EX_rs2 [1] ), .ZN(_04091_ ) );
AOI21_X1 _11834_ ( .A(_04091_ ), .B1(_02133_ ), .B2(\ID_EX_rs2 [1] ), .ZN(_04092_ ) );
OAI211_X1 _11835_ ( .A(_04090_ ), .B(_04092_ ), .C1(_02136_ ), .C2(_02135_ ), .ZN(_04093_ ) );
BUF_X2 _11836_ ( .A(_04093_ ), .Z(_04094_ ) );
CLKBUF_X2 _11837_ ( .A(_04094_ ), .Z(_04095_ ) );
BUF_X2 _11838_ ( .A(_04095_ ), .Z(_04096_ ) );
BUF_X2 _11839_ ( .A(_04096_ ), .Z(_04097_ ) );
OAI21_X1 _11840_ ( .A(_04085_ ), .B1(_02197_ ), .B2(_04097_ ), .ZN(_04098_ ) );
NOR2_X1 _11841_ ( .A1(_04094_ ), .A2(_02161_ ), .ZN(_04099_ ) );
NAND2_X1 _11842_ ( .A1(_04099_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_04100_ ) );
AND2_X1 _11843_ ( .A1(_04098_ ), .A2(_04100_ ), .ZN(_04101_ ) );
INV_X1 _11844_ ( .A(_04101_ ), .ZN(_04102_ ) );
XNOR2_X1 _11845_ ( .A(_02172_ ), .B(_04102_ ), .ZN(_04103_ ) );
OR2_X1 _11846_ ( .A1(_04076_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04104_ ) );
BUF_X4 _11847_ ( .A(_04067_ ), .Z(_04105_ ) );
OAI211_X1 _11848_ ( .A(_04104_ ), .B(_04105_ ), .C1(fanout_net_27 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04106_ ) );
OR2_X1 _11849_ ( .A1(fanout_net_27 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04107_ ) );
BUF_X4 _11850_ ( .A(_04076_ ), .Z(_04108_ ) );
OAI211_X1 _11851_ ( .A(_04107_ ), .B(fanout_net_36 ), .C1(_04108_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04109_ ) );
NAND3_X1 _11852_ ( .A1(_04106_ ), .A2(fanout_net_38 ), .A3(_04109_ ), .ZN(_04110_ ) );
MUX2_X1 _11853_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04111_ ) );
MUX2_X1 _11854_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04112_ ) );
MUX2_X1 _11855_ ( .A(_04111_ ), .B(_04112_ ), .S(_04105_ ), .Z(_04113_ ) );
OAI211_X1 _11856_ ( .A(_04050_ ), .B(_04110_ ), .C1(_04113_ ), .C2(fanout_net_38 ), .ZN(_04114_ ) );
NOR2_X1 _11857_ ( .A1(fanout_net_27 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04115_ ) );
BUF_X4 _11858_ ( .A(_04067_ ), .Z(_04116_ ) );
OAI21_X1 _11859_ ( .A(_04116_ ), .B1(_04108_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04117_ ) );
MUX2_X1 _11860_ ( .A(_02994_ ), .B(_02995_ ), .S(fanout_net_27 ), .Z(_04118_ ) );
OAI221_X1 _11861_ ( .A(_04073_ ), .B1(_04115_ ), .B2(_04117_ ), .C1(_04118_ ), .C2(_04105_ ), .ZN(_04119_ ) );
MUX2_X1 _11862_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04120_ ) );
MUX2_X1 _11863_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04121_ ) );
MUX2_X1 _11864_ ( .A(_04120_ ), .B(_04121_ ), .S(fanout_net_36 ), .Z(_04122_ ) );
BUF_X4 _11865_ ( .A(_04073_ ), .Z(_04123_ ) );
OAI211_X1 _11866_ ( .A(fanout_net_39 ), .B(_04119_ ), .C1(_04122_ ), .C2(_04123_ ), .ZN(_04124_ ) );
OAI211_X1 _11867_ ( .A(_04114_ ), .B(_04124_ ), .C1(_04097_ ), .C2(_02164_ ), .ZN(_04125_ ) );
OR3_X1 _11868_ ( .A1(_04097_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02164_ ), .ZN(_04126_ ) );
NAND2_X1 _11869_ ( .A1(_04125_ ), .A2(_04126_ ), .ZN(_04127_ ) );
XNOR2_X1 _11870_ ( .A(_03004_ ), .B(_04127_ ), .ZN(_04128_ ) );
AND2_X1 _11871_ ( .A1(_04103_ ), .A2(_04128_ ), .ZN(_04129_ ) );
OR2_X1 _11872_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04130_ ) );
OAI211_X1 _11873_ ( .A(_04130_ ), .B(fanout_net_36 ), .C1(_04055_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04131_ ) );
NAND2_X1 _11874_ ( .A1(_02205_ ), .A2(fanout_net_27 ), .ZN(_04132_ ) );
OAI211_X1 _11875_ ( .A(_04132_ ), .B(_04067_ ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04133_ ) );
NAND3_X1 _11876_ ( .A1(_04131_ ), .A2(_04133_ ), .A3(_04061_ ), .ZN(_04134_ ) );
MUX2_X1 _11877_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04135_ ) );
MUX2_X1 _11878_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04136_ ) );
MUX2_X1 _11879_ ( .A(_04135_ ), .B(_04136_ ), .S(_04066_ ), .Z(_04137_ ) );
OAI211_X1 _11880_ ( .A(_04050_ ), .B(_04134_ ), .C1(_04137_ ), .C2(_04061_ ), .ZN(_04138_ ) );
OR2_X1 _11881_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04139_ ) );
OAI211_X1 _11882_ ( .A(_04139_ ), .B(_04067_ ), .C1(_04055_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04140_ ) );
NAND2_X1 _11883_ ( .A1(_02215_ ), .A2(fanout_net_27 ), .ZN(_04141_ ) );
OAI211_X1 _11884_ ( .A(_04141_ ), .B(fanout_net_36 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04142_ ) );
NAND3_X1 _11885_ ( .A1(_04140_ ), .A2(_04142_ ), .A3(fanout_net_38 ), .ZN(_04143_ ) );
MUX2_X1 _11886_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04144_ ) );
MUX2_X1 _11887_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04145_ ) );
MUX2_X1 _11888_ ( .A(_04144_ ), .B(_04145_ ), .S(fanout_net_36 ), .Z(_04146_ ) );
OAI211_X1 _11889_ ( .A(fanout_net_39 ), .B(_04143_ ), .C1(_04146_ ), .C2(fanout_net_38 ), .ZN(_04147_ ) );
NAND2_X1 _11890_ ( .A1(_04138_ ), .A2(_04147_ ), .ZN(_04148_ ) );
OAI21_X1 _11891_ ( .A(_04148_ ), .B1(_02197_ ), .B2(_04096_ ), .ZN(_04149_ ) );
NAND2_X1 _11892_ ( .A1(_04099_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_04150_ ) );
AND2_X1 _11893_ ( .A1(_04149_ ), .A2(_04150_ ), .ZN(_04151_ ) );
XNOR2_X1 _11894_ ( .A(_02225_ ), .B(_04151_ ), .ZN(_04152_ ) );
OR2_X1 _11895_ ( .A1(fanout_net_27 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04153_ ) );
OAI211_X1 _11896_ ( .A(_04153_ ), .B(fanout_net_36 ), .C1(_04076_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04154_ ) );
NAND2_X1 _11897_ ( .A1(_02177_ ), .A2(fanout_net_27 ), .ZN(_04155_ ) );
OAI211_X1 _11898_ ( .A(_04155_ ), .B(_04116_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04156_ ) );
NAND3_X1 _11899_ ( .A1(_04154_ ), .A2(_04156_ ), .A3(_04073_ ), .ZN(_04157_ ) );
MUX2_X1 _11900_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04158_ ) );
MUX2_X1 _11901_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04159_ ) );
MUX2_X1 _11902_ ( .A(_04158_ ), .B(_04159_ ), .S(_04116_ ), .Z(_04160_ ) );
OAI211_X1 _11903_ ( .A(fanout_net_39 ), .B(_04157_ ), .C1(_04160_ ), .C2(_04123_ ), .ZN(_04161_ ) );
OR2_X1 _11904_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04162_ ) );
OAI211_X1 _11905_ ( .A(_04162_ ), .B(_04116_ ), .C1(_04076_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04163_ ) );
NAND2_X1 _11906_ ( .A1(_02187_ ), .A2(fanout_net_28 ), .ZN(_04164_ ) );
OAI211_X1 _11907_ ( .A(_04164_ ), .B(fanout_net_36 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04165_ ) );
NAND3_X1 _11908_ ( .A1(_04163_ ), .A2(_04165_ ), .A3(_04073_ ), .ZN(_04166_ ) );
MUX2_X1 _11909_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04167_ ) );
MUX2_X1 _11910_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04168_ ) );
MUX2_X1 _11911_ ( .A(_04167_ ), .B(_04168_ ), .S(_04116_ ), .Z(_04169_ ) );
OAI211_X1 _11912_ ( .A(_04050_ ), .B(_04166_ ), .C1(_04169_ ), .C2(_04123_ ), .ZN(_04170_ ) );
OAI211_X1 _11913_ ( .A(_04161_ ), .B(_04170_ ), .C1(_04097_ ), .C2(_02164_ ), .ZN(_04171_ ) );
OR3_X1 _11914_ ( .A1(_04096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02197_ ), .ZN(_04172_ ) );
NAND2_X1 _11915_ ( .A1(_04171_ ), .A2(_04172_ ), .ZN(_04173_ ) );
AND3_X1 _11916_ ( .A1(_04173_ ), .A2(_02196_ ), .A3(_02198_ ), .ZN(_04174_ ) );
AOI21_X1 _11917_ ( .A(_04173_ ), .B1(_02196_ ), .B2(_02198_ ), .ZN(_04175_ ) );
NOR2_X1 _11918_ ( .A1(_04174_ ), .A2(_04175_ ), .ZN(_04176_ ) );
NAND3_X1 _11919_ ( .A1(_04129_ ), .A2(_04152_ ), .A3(_04176_ ), .ZN(_04177_ ) );
OR2_X1 _11920_ ( .A1(_04076_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04178_ ) );
OAI211_X1 _11921_ ( .A(_04178_ ), .B(fanout_net_36 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04179_ ) );
OR2_X1 _11922_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04180_ ) );
OAI211_X1 _11923_ ( .A(_04180_ ), .B(_04105_ ), .C1(_04108_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04181_ ) );
NAND3_X1 _11924_ ( .A1(_04179_ ), .A2(_04123_ ), .A3(_04181_ ), .ZN(_04182_ ) );
MUX2_X1 _11925_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04183_ ) );
MUX2_X1 _11926_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04184_ ) );
MUX2_X1 _11927_ ( .A(_04183_ ), .B(_04184_ ), .S(_04116_ ), .Z(_04185_ ) );
OAI211_X1 _11928_ ( .A(fanout_net_39 ), .B(_04182_ ), .C1(_04185_ ), .C2(_04123_ ), .ZN(_04186_ ) );
OR2_X1 _11929_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04187_ ) );
OAI211_X1 _11930_ ( .A(_04187_ ), .B(_04116_ ), .C1(_04108_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04188_ ) );
NOR2_X1 _11931_ ( .A1(_04108_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04189_ ) );
OAI21_X1 _11932_ ( .A(fanout_net_36 ), .B1(fanout_net_28 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04190_ ) );
OAI211_X1 _11933_ ( .A(_04188_ ), .B(_04073_ ), .C1(_04189_ ), .C2(_04190_ ), .ZN(_04191_ ) );
MUX2_X1 _11934_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04192_ ) );
MUX2_X1 _11935_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04193_ ) );
MUX2_X1 _11936_ ( .A(_04192_ ), .B(_04193_ ), .S(_04116_ ), .Z(_04194_ ) );
OAI211_X1 _11937_ ( .A(_04050_ ), .B(_04191_ ), .C1(_04194_ ), .C2(_04123_ ), .ZN(_04195_ ) );
OAI211_X1 _11938_ ( .A(_04186_ ), .B(_04195_ ), .C1(_04097_ ), .C2(_02164_ ), .ZN(_04196_ ) );
INV_X1 _11939_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04197_ ) );
OR3_X1 _11940_ ( .A1(_04097_ ), .A2(_04197_ ), .A3(_02164_ ), .ZN(_04198_ ) );
NAND2_X1 _11941_ ( .A1(_04196_ ), .A2(_04198_ ), .ZN(_04199_ ) );
INV_X1 _11942_ ( .A(_04199_ ), .ZN(_04200_ ) );
NAND2_X1 _11943_ ( .A1(_02248_ ), .A2(_04200_ ), .ZN(_04201_ ) );
NAND3_X1 _11944_ ( .A1(_02246_ ), .A2(_02247_ ), .A3(_04199_ ), .ZN(_04202_ ) );
AND2_X1 _11945_ ( .A1(_04201_ ), .A2(_04202_ ), .ZN(_04203_ ) );
OR2_X1 _11946_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04204_ ) );
OAI211_X1 _11947_ ( .A(_04204_ ), .B(_04105_ ), .C1(_04108_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04205_ ) );
OR2_X1 _11948_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04206_ ) );
OAI211_X1 _11949_ ( .A(_04206_ ), .B(fanout_net_36 ), .C1(_04108_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04207_ ) );
NAND3_X1 _11950_ ( .A1(_04205_ ), .A2(_04207_ ), .A3(fanout_net_38 ), .ZN(_04208_ ) );
MUX2_X1 _11951_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04209_ ) );
MUX2_X1 _11952_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04210_ ) );
MUX2_X1 _11953_ ( .A(_04209_ ), .B(_04210_ ), .S(_04105_ ), .Z(_04211_ ) );
OAI211_X1 _11954_ ( .A(_04050_ ), .B(_04208_ ), .C1(_04211_ ), .C2(fanout_net_38 ), .ZN(_04212_ ) );
NOR2_X1 _11955_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04213_ ) );
OAI21_X1 _11956_ ( .A(_04116_ ), .B1(_04108_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04214_ ) );
MUX2_X1 _11957_ ( .A(_02945_ ), .B(_02946_ ), .S(fanout_net_28 ), .Z(_04215_ ) );
OAI221_X1 _11958_ ( .A(_04123_ ), .B1(_04213_ ), .B2(_04214_ ), .C1(_04215_ ), .C2(_04105_ ), .ZN(_04216_ ) );
MUX2_X1 _11959_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04217_ ) );
MUX2_X1 _11960_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04218_ ) );
MUX2_X1 _11961_ ( .A(_04217_ ), .B(_04218_ ), .S(fanout_net_36 ), .Z(_04219_ ) );
OAI211_X1 _11962_ ( .A(fanout_net_39 ), .B(_04216_ ), .C1(_04219_ ), .C2(_04123_ ), .ZN(_04220_ ) );
OAI211_X1 _11963_ ( .A(_04212_ ), .B(_04220_ ), .C1(_04097_ ), .C2(_02164_ ), .ZN(_04221_ ) );
INV_X1 _11964_ ( .A(\EX_LS_result_reg [26] ), .ZN(_04222_ ) );
OR3_X1 _11965_ ( .A1(_04097_ ), .A2(_04222_ ), .A3(_02164_ ), .ZN(_04223_ ) );
NAND2_X1 _11966_ ( .A1(_04221_ ), .A2(_04223_ ), .ZN(_04224_ ) );
XNOR2_X1 _11967_ ( .A(_02965_ ), .B(_04224_ ), .ZN(_04225_ ) );
AND2_X1 _11968_ ( .A1(_04203_ ), .A2(_04225_ ), .ZN(_04226_ ) );
OR2_X1 _11969_ ( .A1(_04055_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04227_ ) );
OAI211_X1 _11970_ ( .A(_04227_ ), .B(_04116_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04228_ ) );
NAND2_X1 _11971_ ( .A1(_02920_ ), .A2(fanout_net_28 ), .ZN(_04229_ ) );
OAI211_X1 _11972_ ( .A(_04229_ ), .B(fanout_net_36 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04230_ ) );
NAND3_X1 _11973_ ( .A1(_04228_ ), .A2(_04073_ ), .A3(_04230_ ), .ZN(_04231_ ) );
MUX2_X1 _11974_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04232_ ) );
MUX2_X1 _11975_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04233_ ) );
MUX2_X1 _11976_ ( .A(_04232_ ), .B(_04233_ ), .S(_04067_ ), .Z(_04234_ ) );
OAI211_X1 _11977_ ( .A(fanout_net_39 ), .B(_04231_ ), .C1(_04234_ ), .C2(_04073_ ), .ZN(_04235_ ) );
OR2_X1 _11978_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04236_ ) );
OAI211_X1 _11979_ ( .A(_04236_ ), .B(_04067_ ), .C1(_04076_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04237_ ) );
NAND2_X1 _11980_ ( .A1(_02930_ ), .A2(fanout_net_29 ), .ZN(_04238_ ) );
OAI211_X1 _11981_ ( .A(_04238_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04239_ ) );
NAND3_X1 _11982_ ( .A1(_04237_ ), .A2(_04239_ ), .A3(_04073_ ), .ZN(_04240_ ) );
MUX2_X1 _11983_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04241_ ) );
MUX2_X1 _11984_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04242_ ) );
MUX2_X1 _11985_ ( .A(_04241_ ), .B(_04242_ ), .S(_04067_ ), .Z(_04243_ ) );
OAI211_X1 _11986_ ( .A(_04050_ ), .B(_04240_ ), .C1(_04243_ ), .C2(_04073_ ), .ZN(_04244_ ) );
OAI211_X1 _11987_ ( .A(_04235_ ), .B(_04244_ ), .C1(_04097_ ), .C2(_02197_ ), .ZN(_04245_ ) );
INV_X1 _11988_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04246_ ) );
OR3_X1 _11989_ ( .A1(_04096_ ), .A2(_04246_ ), .A3(_02197_ ), .ZN(_04247_ ) );
NAND2_X1 _11990_ ( .A1(_04245_ ), .A2(_04247_ ), .ZN(_04248_ ) );
XNOR2_X1 _11991_ ( .A(_02940_ ), .B(_04248_ ), .ZN(_04249_ ) );
NAND2_X1 _11992_ ( .A1(_04099_ ), .A2(\EX_LS_result_reg [24] ), .ZN(_04250_ ) );
OR2_X1 _11993_ ( .A1(_04076_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04251_ ) );
OAI211_X1 _11994_ ( .A(_04251_ ), .B(_04105_ ), .C1(fanout_net_29 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04252_ ) );
OR2_X1 _11995_ ( .A1(_04076_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04253_ ) );
OAI211_X1 _11996_ ( .A(_04253_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04254_ ) );
NAND3_X1 _11997_ ( .A1(_04252_ ), .A2(_04254_ ), .A3(fanout_net_38 ), .ZN(_04255_ ) );
MUX2_X1 _11998_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04256_ ) );
MUX2_X1 _11999_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04257_ ) );
MUX2_X1 _12000_ ( .A(_04256_ ), .B(_04257_ ), .S(_04105_ ), .Z(_04258_ ) );
OAI211_X1 _12001_ ( .A(_04050_ ), .B(_04255_ ), .C1(_04258_ ), .C2(fanout_net_38 ), .ZN(_04259_ ) );
NOR2_X1 _12002_ ( .A1(_04108_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04260_ ) );
OAI21_X1 _12003_ ( .A(fanout_net_36 ), .B1(fanout_net_29 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04261_ ) );
NOR2_X1 _12004_ ( .A1(fanout_net_29 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04262_ ) );
OAI21_X1 _12005_ ( .A(_04105_ ), .B1(_04108_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04263_ ) );
OAI221_X1 _12006_ ( .A(_04123_ ), .B1(_04260_ ), .B2(_04261_ ), .C1(_04262_ ), .C2(_04263_ ), .ZN(_04264_ ) );
MUX2_X1 _12007_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04265_ ) );
MUX2_X1 _12008_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04266_ ) );
MUX2_X1 _12009_ ( .A(_04265_ ), .B(_04266_ ), .S(fanout_net_36 ), .Z(_04267_ ) );
OAI211_X1 _12010_ ( .A(fanout_net_39 ), .B(_04264_ ), .C1(_04267_ ), .C2(_04123_ ), .ZN(_04268_ ) );
OAI211_X1 _12011_ ( .A(_04259_ ), .B(_04268_ ), .C1(_04097_ ), .C2(_02164_ ), .ZN(_04269_ ) );
NAND2_X1 _12012_ ( .A1(_04250_ ), .A2(_04269_ ), .ZN(_04270_ ) );
XNOR2_X1 _12013_ ( .A(_02271_ ), .B(_04270_ ), .ZN(_04271_ ) );
NAND3_X1 _12014_ ( .A1(_04226_ ), .A2(_04249_ ), .A3(_04271_ ), .ZN(_04272_ ) );
NOR2_X1 _12015_ ( .A1(_04177_ ), .A2(_04272_ ), .ZN(_04273_ ) );
CLKBUF_X2 _12016_ ( .A(_04051_ ), .Z(_04274_ ) );
BUF_X2 _12017_ ( .A(_04274_ ), .Z(_04275_ ) );
OR2_X1 _12018_ ( .A1(_04275_ ), .A2(\myreg.Reg[3][18] ), .ZN(_04276_ ) );
OAI211_X1 _12019_ ( .A(_04276_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[2][18] ), .ZN(_04277_ ) );
BUF_X4 _12020_ ( .A(_04058_ ), .Z(_04278_ ) );
BUF_X4 _12021_ ( .A(_04278_ ), .Z(_04279_ ) );
OR2_X1 _12022_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][18] ), .ZN(_04280_ ) );
BUF_X4 _12023_ ( .A(_04063_ ), .Z(_04281_ ) );
BUF_X4 _12024_ ( .A(_04281_ ), .Z(_04282_ ) );
BUF_X2 _12025_ ( .A(_04052_ ), .Z(_04283_ ) );
BUF_X2 _12026_ ( .A(_04283_ ), .Z(_04284_ ) );
OAI211_X1 _12027_ ( .A(_04280_ ), .B(_04282_ ), .C1(_04284_ ), .C2(\myreg.Reg[1][18] ), .ZN(_04285_ ) );
NAND3_X1 _12028_ ( .A1(_04277_ ), .A2(_04279_ ), .A3(_04285_ ), .ZN(_04286_ ) );
MUX2_X1 _12029_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_29 ), .Z(_04287_ ) );
MUX2_X1 _12030_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_29 ), .Z(_04288_ ) );
MUX2_X1 _12031_ ( .A(_04287_ ), .B(_04288_ ), .S(_04282_ ), .Z(_04289_ ) );
BUF_X4 _12032_ ( .A(_04278_ ), .Z(_04290_ ) );
OAI211_X1 _12033_ ( .A(_04049_ ), .B(_04286_ ), .C1(_04289_ ), .C2(_04290_ ), .ZN(_04291_ ) );
OR2_X1 _12034_ ( .A1(_04275_ ), .A2(\myreg.Reg[15][18] ), .ZN(_04292_ ) );
OAI211_X1 _12035_ ( .A(_04292_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[14][18] ), .ZN(_04293_ ) );
OR2_X1 _12036_ ( .A1(_04275_ ), .A2(\myreg.Reg[13][18] ), .ZN(_04294_ ) );
OAI211_X1 _12037_ ( .A(_04294_ ), .B(_04282_ ), .C1(fanout_net_29 ), .C2(\myreg.Reg[12][18] ), .ZN(_04295_ ) );
NAND3_X1 _12038_ ( .A1(_04293_ ), .A2(_04295_ ), .A3(fanout_net_38 ), .ZN(_04296_ ) );
MUX2_X1 _12039_ ( .A(\myreg.Reg[8][18] ), .B(\myreg.Reg[9][18] ), .S(fanout_net_29 ), .Z(_04297_ ) );
MUX2_X1 _12040_ ( .A(\myreg.Reg[10][18] ), .B(\myreg.Reg[11][18] ), .S(fanout_net_29 ), .Z(_04298_ ) );
MUX2_X1 _12041_ ( .A(_04297_ ), .B(_04298_ ), .S(fanout_net_36 ), .Z(_04299_ ) );
OAI211_X1 _12042_ ( .A(fanout_net_39 ), .B(_04296_ ), .C1(_04299_ ), .C2(fanout_net_38 ), .ZN(_04300_ ) );
CLKBUF_X2 _12043_ ( .A(_04094_ ), .Z(_04301_ ) );
BUF_X2 _12044_ ( .A(_04301_ ), .Z(_04302_ ) );
OAI211_X1 _12045_ ( .A(_04291_ ), .B(_04300_ ), .C1(_04302_ ), .C2(_02331_ ), .ZN(_04303_ ) );
OR3_X1 _12046_ ( .A1(_04095_ ), .A2(\EX_LS_result_reg [18] ), .A3(_02304_ ), .ZN(_04304_ ) );
NAND2_X1 _12047_ ( .A1(_04303_ ), .A2(_04304_ ), .ZN(_04305_ ) );
XOR2_X1 _12048_ ( .A(_02406_ ), .B(_04305_ ), .Z(_04306_ ) );
OR2_X1 _12049_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][19] ), .ZN(_04307_ ) );
OAI211_X1 _12050_ ( .A(_04307_ ), .B(_04282_ ), .C1(_04054_ ), .C2(\myreg.Reg[9][19] ), .ZN(_04308_ ) );
OR2_X1 _12051_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[10][19] ), .ZN(_04309_ ) );
OAI211_X1 _12052_ ( .A(_04309_ ), .B(fanout_net_36 ), .C1(_04054_ ), .C2(\myreg.Reg[11][19] ), .ZN(_04310_ ) );
NAND3_X1 _12053_ ( .A1(_04308_ ), .A2(_04310_ ), .A3(_04279_ ), .ZN(_04311_ ) );
MUX2_X1 _12054_ ( .A(\myreg.Reg[14][19] ), .B(\myreg.Reg[15][19] ), .S(fanout_net_29 ), .Z(_04312_ ) );
MUX2_X1 _12055_ ( .A(\myreg.Reg[12][19] ), .B(\myreg.Reg[13][19] ), .S(fanout_net_29 ), .Z(_04313_ ) );
BUF_X4 _12056_ ( .A(_04281_ ), .Z(_04314_ ) );
MUX2_X1 _12057_ ( .A(_04312_ ), .B(_04313_ ), .S(_04314_ ), .Z(_04315_ ) );
OAI211_X1 _12058_ ( .A(fanout_net_39 ), .B(_04311_ ), .C1(_04315_ ), .C2(_04290_ ), .ZN(_04316_ ) );
OR2_X1 _12059_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][19] ), .ZN(_04317_ ) );
OAI211_X1 _12060_ ( .A(_04317_ ), .B(_04314_ ), .C1(_04054_ ), .C2(\myreg.Reg[1][19] ), .ZN(_04318_ ) );
NOR2_X1 _12061_ ( .A1(_04284_ ), .A2(\myreg.Reg[3][19] ), .ZN(_04319_ ) );
OAI21_X1 _12062_ ( .A(fanout_net_36 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[2][19] ), .ZN(_04320_ ) );
OAI211_X1 _12063_ ( .A(_04318_ ), .B(_04060_ ), .C1(_04319_ ), .C2(_04320_ ), .ZN(_04321_ ) );
MUX2_X1 _12064_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_29 ), .Z(_04322_ ) );
MUX2_X1 _12065_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_29 ), .Z(_04323_ ) );
MUX2_X1 _12066_ ( .A(_04322_ ), .B(_04323_ ), .S(_04314_ ), .Z(_04324_ ) );
OAI211_X1 _12067_ ( .A(_04049_ ), .B(_04321_ ), .C1(_04324_ ), .C2(_04290_ ), .ZN(_04325_ ) );
OAI211_X1 _12068_ ( .A(_04316_ ), .B(_04325_ ), .C1(_04302_ ), .C2(_02331_ ), .ZN(_04326_ ) );
OR3_X1 _12069_ ( .A1(_04095_ ), .A2(\EX_LS_result_reg [19] ), .A3(_02162_ ), .ZN(_04327_ ) );
NAND2_X1 _12070_ ( .A1(_04326_ ), .A2(_04327_ ), .ZN(_04328_ ) );
INV_X1 _12071_ ( .A(_04328_ ), .ZN(_04329_ ) );
NAND2_X1 _12072_ ( .A1(_02429_ ), .A2(_02431_ ), .ZN(_04330_ ) );
XNOR2_X1 _12073_ ( .A(_04329_ ), .B(_04330_ ), .ZN(_04331_ ) );
AND2_X1 _12074_ ( .A1(_04306_ ), .A2(_04331_ ), .ZN(_04332_ ) );
OR2_X1 _12075_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][17] ), .ZN(_04333_ ) );
OAI211_X1 _12076_ ( .A(_04333_ ), .B(_04282_ ), .C1(_04054_ ), .C2(\myreg.Reg[9][17] ), .ZN(_04334_ ) );
OR2_X1 _12077_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[10][17] ), .ZN(_04335_ ) );
OAI211_X1 _12078_ ( .A(_04335_ ), .B(fanout_net_36 ), .C1(_04054_ ), .C2(\myreg.Reg[11][17] ), .ZN(_04336_ ) );
NAND3_X1 _12079_ ( .A1(_04334_ ), .A2(_04336_ ), .A3(_04060_ ), .ZN(_04337_ ) );
MUX2_X1 _12080_ ( .A(\myreg.Reg[14][17] ), .B(\myreg.Reg[15][17] ), .S(fanout_net_30 ), .Z(_04338_ ) );
MUX2_X1 _12081_ ( .A(\myreg.Reg[12][17] ), .B(\myreg.Reg[13][17] ), .S(fanout_net_30 ), .Z(_04339_ ) );
MUX2_X1 _12082_ ( .A(_04338_ ), .B(_04339_ ), .S(_04065_ ), .Z(_04340_ ) );
OAI211_X1 _12083_ ( .A(fanout_net_39 ), .B(_04337_ ), .C1(_04340_ ), .C2(_04290_ ), .ZN(_04341_ ) );
BUF_X4 _12084_ ( .A(_04059_ ), .Z(_04342_ ) );
BUF_X2 _12085_ ( .A(_04274_ ), .Z(_04343_ ) );
NOR2_X1 _12086_ ( .A1(_04343_ ), .A2(\myreg.Reg[3][17] ), .ZN(_04344_ ) );
OAI21_X1 _12087_ ( .A(fanout_net_36 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[2][17] ), .ZN(_04345_ ) );
NOR2_X1 _12088_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[0][17] ), .ZN(_04346_ ) );
OAI21_X1 _12089_ ( .A(_04065_ ), .B1(_04343_ ), .B2(\myreg.Reg[1][17] ), .ZN(_04347_ ) );
OAI221_X1 _12090_ ( .A(_04342_ ), .B1(_04344_ ), .B2(_04345_ ), .C1(_04346_ ), .C2(_04347_ ), .ZN(_04348_ ) );
MUX2_X1 _12091_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_30 ), .Z(_04349_ ) );
MUX2_X1 _12092_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_30 ), .Z(_04350_ ) );
MUX2_X1 _12093_ ( .A(_04349_ ), .B(_04350_ ), .S(_04065_ ), .Z(_04351_ ) );
OAI211_X1 _12094_ ( .A(_04049_ ), .B(_04348_ ), .C1(_04351_ ), .C2(_04290_ ), .ZN(_04352_ ) );
OAI211_X1 _12095_ ( .A(_04341_ ), .B(_04352_ ), .C1(_04302_ ), .C2(_02331_ ), .ZN(_04353_ ) );
OR3_X1 _12096_ ( .A1(_04095_ ), .A2(\EX_LS_result_reg [17] ), .A3(_02162_ ), .ZN(_04354_ ) );
NAND2_X1 _12097_ ( .A1(_04353_ ), .A2(_04354_ ), .ZN(_04355_ ) );
INV_X1 _12098_ ( .A(_04355_ ), .ZN(_04356_ ) );
XNOR2_X1 _12099_ ( .A(_04356_ ), .B(_02458_ ), .ZN(_04357_ ) );
OR2_X1 _12100_ ( .A1(_04054_ ), .A2(\myreg.Reg[1][16] ), .ZN(_04358_ ) );
OAI211_X1 _12101_ ( .A(_04358_ ), .B(_04066_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[0][16] ), .ZN(_04359_ ) );
OR2_X1 _12102_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[2][16] ), .ZN(_04360_ ) );
OAI211_X1 _12103_ ( .A(_04360_ ), .B(fanout_net_36 ), .C1(_04055_ ), .C2(\myreg.Reg[3][16] ), .ZN(_04361_ ) );
NAND3_X1 _12104_ ( .A1(_04359_ ), .A2(_04061_ ), .A3(_04361_ ), .ZN(_04362_ ) );
MUX2_X1 _12105_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_30 ), .Z(_04363_ ) );
MUX2_X1 _12106_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_30 ), .Z(_04364_ ) );
MUX2_X1 _12107_ ( .A(_04363_ ), .B(_04364_ ), .S(_04066_ ), .Z(_04365_ ) );
OAI211_X1 _12108_ ( .A(_04050_ ), .B(_04362_ ), .C1(_04365_ ), .C2(_04061_ ), .ZN(_04366_ ) );
OR2_X1 _12109_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[14][16] ), .ZN(_04367_ ) );
OAI211_X1 _12110_ ( .A(_04367_ ), .B(fanout_net_36 ), .C1(_04055_ ), .C2(\myreg.Reg[15][16] ), .ZN(_04368_ ) );
OR2_X1 _12111_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[12][16] ), .ZN(_04369_ ) );
OAI211_X1 _12112_ ( .A(_04369_ ), .B(_04066_ ), .C1(_04284_ ), .C2(\myreg.Reg[13][16] ), .ZN(_04370_ ) );
NAND3_X1 _12113_ ( .A1(_04368_ ), .A2(_04370_ ), .A3(fanout_net_38 ), .ZN(_04371_ ) );
MUX2_X1 _12114_ ( .A(\myreg.Reg[8][16] ), .B(\myreg.Reg[9][16] ), .S(fanout_net_30 ), .Z(_04372_ ) );
MUX2_X1 _12115_ ( .A(\myreg.Reg[10][16] ), .B(\myreg.Reg[11][16] ), .S(fanout_net_30 ), .Z(_04373_ ) );
MUX2_X1 _12116_ ( .A(_04372_ ), .B(_04373_ ), .S(fanout_net_36 ), .Z(_04374_ ) );
OAI211_X1 _12117_ ( .A(fanout_net_39 ), .B(_04371_ ), .C1(_04374_ ), .C2(fanout_net_38 ), .ZN(_04375_ ) );
OAI211_X1 _12118_ ( .A(_04366_ ), .B(_04375_ ), .C1(_04096_ ), .C2(_02163_ ), .ZN(_04376_ ) );
OR3_X1 _12119_ ( .A1(_04096_ ), .A2(\EX_LS_result_reg [16] ), .A3(_02163_ ), .ZN(_04377_ ) );
NAND2_X1 _12120_ ( .A1(_04376_ ), .A2(_04377_ ), .ZN(_04378_ ) );
INV_X1 _12121_ ( .A(_04378_ ), .ZN(_04379_ ) );
XNOR2_X1 _12122_ ( .A(_04379_ ), .B(_02480_ ), .ZN(_04380_ ) );
AND3_X1 _12123_ ( .A1(_04332_ ), .A2(_04357_ ), .A3(_04380_ ), .ZN(_04381_ ) );
OR2_X1 _12124_ ( .A1(_04053_ ), .A2(\myreg.Reg[9][23] ), .ZN(_04382_ ) );
OAI211_X1 _12125_ ( .A(_04382_ ), .B(_04065_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[8][23] ), .ZN(_04383_ ) );
OR2_X1 _12126_ ( .A1(_04053_ ), .A2(\myreg.Reg[11][23] ), .ZN(_04384_ ) );
OAI211_X1 _12127_ ( .A(_04384_ ), .B(fanout_net_37 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[10][23] ), .ZN(_04385_ ) );
NAND3_X1 _12128_ ( .A1(_04383_ ), .A2(_04385_ ), .A3(_04342_ ), .ZN(_04386_ ) );
MUX2_X1 _12129_ ( .A(\myreg.Reg[14][23] ), .B(\myreg.Reg[15][23] ), .S(fanout_net_30 ), .Z(_04387_ ) );
MUX2_X1 _12130_ ( .A(\myreg.Reg[12][23] ), .B(\myreg.Reg[13][23] ), .S(fanout_net_30 ), .Z(_04388_ ) );
BUF_X4 _12131_ ( .A(_04064_ ), .Z(_04389_ ) );
MUX2_X1 _12132_ ( .A(_04387_ ), .B(_04388_ ), .S(_04389_ ), .Z(_04390_ ) );
OAI211_X1 _12133_ ( .A(fanout_net_39 ), .B(_04386_ ), .C1(_04390_ ), .C2(_04279_ ), .ZN(_04391_ ) );
BUF_X4 _12134_ ( .A(_04064_ ), .Z(_04392_ ) );
BUF_X2 _12135_ ( .A(_04274_ ), .Z(_04393_ ) );
OAI21_X1 _12136_ ( .A(_04392_ ), .B1(_04393_ ), .B2(\myreg.Reg[1][23] ), .ZN(_04394_ ) );
NOR2_X1 _12137_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[0][23] ), .ZN(_04395_ ) );
NOR2_X1 _12138_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[2][23] ), .ZN(_04396_ ) );
OAI21_X1 _12139_ ( .A(fanout_net_37 ), .B1(_04393_ ), .B2(\myreg.Reg[3][23] ), .ZN(_04397_ ) );
OAI221_X1 _12140_ ( .A(_04342_ ), .B1(_04394_ ), .B2(_04395_ ), .C1(_04396_ ), .C2(_04397_ ), .ZN(_04398_ ) );
MUX2_X1 _12141_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_30 ), .Z(_04399_ ) );
MUX2_X1 _12142_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_30 ), .Z(_04400_ ) );
MUX2_X1 _12143_ ( .A(_04399_ ), .B(_04400_ ), .S(_04389_ ), .Z(_04401_ ) );
OAI211_X1 _12144_ ( .A(_04048_ ), .B(_04398_ ), .C1(_04401_ ), .C2(_04279_ ), .ZN(_04402_ ) );
OAI211_X1 _12145_ ( .A(_04391_ ), .B(_04402_ ), .C1(_04302_ ), .C2(_02304_ ), .ZN(_04403_ ) );
OR3_X1 _12146_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [23] ), .A3(_02456_ ), .ZN(_04404_ ) );
NAND2_X1 _12147_ ( .A1(_04403_ ), .A2(_04404_ ), .ZN(_04405_ ) );
INV_X1 _12148_ ( .A(_04405_ ), .ZN(_04406_ ) );
XNOR2_X1 _12149_ ( .A(_04406_ ), .B(_02307_ ), .ZN(_04407_ ) );
NOR2_X1 _12150_ ( .A1(_04393_ ), .A2(\myreg.Reg[11][22] ), .ZN(_04408_ ) );
OAI21_X1 _12151_ ( .A(fanout_net_37 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][22] ), .ZN(_04409_ ) );
NOR2_X1 _12152_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][22] ), .ZN(_04410_ ) );
OAI21_X1 _12153_ ( .A(_04389_ ), .B1(_04393_ ), .B2(\myreg.Reg[9][22] ), .ZN(_04411_ ) );
OAI221_X1 _12154_ ( .A(_04342_ ), .B1(_04408_ ), .B2(_04409_ ), .C1(_04410_ ), .C2(_04411_ ), .ZN(_04412_ ) );
MUX2_X1 _12155_ ( .A(\myreg.Reg[12][22] ), .B(\myreg.Reg[13][22] ), .S(fanout_net_30 ), .Z(_04413_ ) );
MUX2_X1 _12156_ ( .A(\myreg.Reg[14][22] ), .B(\myreg.Reg[15][22] ), .S(fanout_net_30 ), .Z(_04414_ ) );
MUX2_X1 _12157_ ( .A(_04413_ ), .B(_04414_ ), .S(fanout_net_37 ), .Z(_04415_ ) );
OAI211_X1 _12158_ ( .A(fanout_net_39 ), .B(_04412_ ), .C1(_04415_ ), .C2(_04279_ ), .ZN(_04416_ ) );
OR2_X1 _12159_ ( .A1(_04053_ ), .A2(\myreg.Reg[5][22] ), .ZN(_04417_ ) );
OAI211_X1 _12160_ ( .A(_04417_ ), .B(_04314_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[4][22] ), .ZN(_04418_ ) );
OR2_X1 _12161_ ( .A1(_04053_ ), .A2(\myreg.Reg[7][22] ), .ZN(_04419_ ) );
OAI211_X1 _12162_ ( .A(_04419_ ), .B(fanout_net_37 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[6][22] ), .ZN(_04420_ ) );
NAND3_X1 _12163_ ( .A1(_04418_ ), .A2(_04420_ ), .A3(fanout_net_38 ), .ZN(_04421_ ) );
MUX2_X1 _12164_ ( .A(\myreg.Reg[2][22] ), .B(\myreg.Reg[3][22] ), .S(fanout_net_30 ), .Z(_04422_ ) );
MUX2_X1 _12165_ ( .A(\myreg.Reg[0][22] ), .B(\myreg.Reg[1][22] ), .S(fanout_net_30 ), .Z(_04423_ ) );
MUX2_X1 _12166_ ( .A(_04422_ ), .B(_04423_ ), .S(_04389_ ), .Z(_04424_ ) );
OAI211_X1 _12167_ ( .A(_04048_ ), .B(_04421_ ), .C1(_04424_ ), .C2(fanout_net_38 ), .ZN(_04425_ ) );
OAI211_X1 _12168_ ( .A(_04416_ ), .B(_04425_ ), .C1(_02331_ ), .C2(_04302_ ), .ZN(_04426_ ) );
OR3_X1 _12169_ ( .A1(_04095_ ), .A2(\EX_LS_result_reg [22] ), .A3(_02456_ ), .ZN(_04427_ ) );
NAND2_X1 _12170_ ( .A1(_04426_ ), .A2(_04427_ ), .ZN(_04428_ ) );
INV_X1 _12171_ ( .A(_04428_ ), .ZN(_04429_ ) );
XNOR2_X1 _12172_ ( .A(_04429_ ), .B(_02333_ ), .ZN(_04430_ ) );
AND2_X1 _12173_ ( .A1(_04407_ ), .A2(_04430_ ), .ZN(_04431_ ) );
OR2_X1 _12174_ ( .A1(_04284_ ), .A2(\myreg.Reg[3][20] ), .ZN(_04432_ ) );
OAI211_X1 _12175_ ( .A(_04432_ ), .B(fanout_net_37 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[2][20] ), .ZN(_04433_ ) );
OR2_X1 _12176_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][20] ), .ZN(_04434_ ) );
OAI211_X1 _12177_ ( .A(_04434_ ), .B(_04066_ ), .C1(_04055_ ), .C2(\myreg.Reg[1][20] ), .ZN(_04435_ ) );
NAND3_X1 _12178_ ( .A1(_04433_ ), .A2(_04061_ ), .A3(_04435_ ), .ZN(_04436_ ) );
MUX2_X1 _12179_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_31 ), .Z(_04437_ ) );
MUX2_X1 _12180_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_31 ), .Z(_04438_ ) );
MUX2_X1 _12181_ ( .A(_04437_ ), .B(_04438_ ), .S(_04066_ ), .Z(_04439_ ) );
OAI211_X1 _12182_ ( .A(_04050_ ), .B(_04436_ ), .C1(_04439_ ), .C2(_04061_ ), .ZN(_04440_ ) );
OR2_X1 _12183_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][20] ), .ZN(_04441_ ) );
OAI211_X1 _12184_ ( .A(_04441_ ), .B(fanout_net_37 ), .C1(_04055_ ), .C2(\myreg.Reg[15][20] ), .ZN(_04442_ ) );
OR2_X1 _12185_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[12][20] ), .ZN(_04443_ ) );
OAI211_X1 _12186_ ( .A(_04443_ ), .B(_04066_ ), .C1(_04055_ ), .C2(\myreg.Reg[13][20] ), .ZN(_04444_ ) );
NAND3_X1 _12187_ ( .A1(_04442_ ), .A2(_04444_ ), .A3(fanout_net_38 ), .ZN(_04445_ ) );
MUX2_X1 _12188_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_31 ), .Z(_04446_ ) );
MUX2_X1 _12189_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_31 ), .Z(_04447_ ) );
MUX2_X1 _12190_ ( .A(_04446_ ), .B(_04447_ ), .S(fanout_net_37 ), .Z(_04448_ ) );
OAI211_X1 _12191_ ( .A(fanout_net_39 ), .B(_04445_ ), .C1(_04448_ ), .C2(fanout_net_38 ), .ZN(_04449_ ) );
OAI211_X1 _12192_ ( .A(_04440_ ), .B(_04449_ ), .C1(_04096_ ), .C2(_02163_ ), .ZN(_04450_ ) );
OR3_X1 _12193_ ( .A1(_04096_ ), .A2(\EX_LS_result_reg [20] ), .A3(_02163_ ), .ZN(_04451_ ) );
NAND2_X1 _12194_ ( .A1(_04450_ ), .A2(_04451_ ), .ZN(_04452_ ) );
INV_X1 _12195_ ( .A(_04452_ ), .ZN(_04453_ ) );
XNOR2_X1 _12196_ ( .A(_04453_ ), .B(_02382_ ), .ZN(_04454_ ) );
OR2_X1 _12197_ ( .A1(_04343_ ), .A2(\myreg.Reg[1][21] ), .ZN(_04455_ ) );
OAI211_X1 _12198_ ( .A(_04455_ ), .B(_04066_ ), .C1(\myreg.Reg[0][21] ), .C2(fanout_net_31 ), .ZN(_04456_ ) );
OR2_X1 _12199_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][21] ), .ZN(_04457_ ) );
OAI211_X1 _12200_ ( .A(_04457_ ), .B(fanout_net_37 ), .C1(_04284_ ), .C2(\myreg.Reg[3][21] ), .ZN(_04458_ ) );
NAND3_X1 _12201_ ( .A1(_04456_ ), .A2(_04290_ ), .A3(_04458_ ), .ZN(_04459_ ) );
MUX2_X1 _12202_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_31 ), .Z(_04460_ ) );
MUX2_X1 _12203_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_31 ), .Z(_04461_ ) );
MUX2_X1 _12204_ ( .A(_04460_ ), .B(_04461_ ), .S(_04282_ ), .Z(_04462_ ) );
OAI211_X1 _12205_ ( .A(_04049_ ), .B(_04459_ ), .C1(_04462_ ), .C2(_04061_ ), .ZN(_04463_ ) );
OR2_X1 _12206_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][21] ), .ZN(_04464_ ) );
OAI211_X1 _12207_ ( .A(_04464_ ), .B(fanout_net_37 ), .C1(_04284_ ), .C2(\myreg.Reg[15][21] ), .ZN(_04465_ ) );
OR2_X1 _12208_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[12][21] ), .ZN(_04466_ ) );
OAI211_X1 _12209_ ( .A(_04466_ ), .B(_04066_ ), .C1(_04284_ ), .C2(\myreg.Reg[13][21] ), .ZN(_04467_ ) );
NAND3_X1 _12210_ ( .A1(_04465_ ), .A2(_04467_ ), .A3(fanout_net_38 ), .ZN(_04468_ ) );
MUX2_X1 _12211_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_31 ), .Z(_04469_ ) );
MUX2_X1 _12212_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_31 ), .Z(_04470_ ) );
MUX2_X1 _12213_ ( .A(_04469_ ), .B(_04470_ ), .S(fanout_net_37 ), .Z(_04471_ ) );
OAI211_X1 _12214_ ( .A(fanout_net_39 ), .B(_04468_ ), .C1(_04471_ ), .C2(fanout_net_38 ), .ZN(_04472_ ) );
AOI21_X1 _12215_ ( .A(_04099_ ), .B1(_04463_ ), .B2(_04472_ ), .ZN(_04473_ ) );
INV_X1 _12216_ ( .A(\EX_LS_result_reg [21] ), .ZN(_04474_ ) );
NOR3_X1 _12217_ ( .A1(_04096_ ), .A2(_02163_ ), .A3(_04474_ ), .ZN(_04475_ ) );
NOR2_X1 _12218_ ( .A1(_04473_ ), .A2(_04475_ ), .ZN(_04476_ ) );
NAND2_X1 _12219_ ( .A1(_02356_ ), .A2(_02358_ ), .ZN(_04477_ ) );
AND2_X1 _12220_ ( .A1(_04476_ ), .A2(_04477_ ), .ZN(_04478_ ) );
NOR2_X1 _12221_ ( .A1(_04476_ ), .A2(_04477_ ), .ZN(_04479_ ) );
NOR2_X1 _12222_ ( .A1(_04478_ ), .A2(_04479_ ), .ZN(_04480_ ) );
AND3_X1 _12223_ ( .A1(_04431_ ), .A2(_04454_ ), .A3(_04480_ ), .ZN(_04481_ ) );
AND2_X1 _12224_ ( .A1(_04381_ ), .A2(_04481_ ), .ZN(_04482_ ) );
OR2_X1 _12225_ ( .A1(_04283_ ), .A2(\myreg.Reg[11][10] ), .ZN(_04483_ ) );
OAI211_X1 _12226_ ( .A(_04483_ ), .B(fanout_net_37 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[10][10] ), .ZN(_04484_ ) );
OR2_X1 _12227_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][10] ), .ZN(_04485_ ) );
OAI211_X1 _12228_ ( .A(_04485_ ), .B(_04314_ ), .C1(_04054_ ), .C2(\myreg.Reg[9][10] ), .ZN(_04486_ ) );
NAND3_X1 _12229_ ( .A1(_04484_ ), .A2(_04060_ ), .A3(_04486_ ), .ZN(_04487_ ) );
MUX2_X1 _12230_ ( .A(\myreg.Reg[14][10] ), .B(\myreg.Reg[15][10] ), .S(fanout_net_31 ), .Z(_04488_ ) );
MUX2_X1 _12231_ ( .A(\myreg.Reg[12][10] ), .B(\myreg.Reg[13][10] ), .S(fanout_net_31 ), .Z(_04489_ ) );
MUX2_X1 _12232_ ( .A(_04488_ ), .B(_04489_ ), .S(_04065_ ), .Z(_04490_ ) );
OAI211_X1 _12233_ ( .A(fanout_net_39 ), .B(_04487_ ), .C1(_04490_ ), .C2(_04290_ ), .ZN(_04491_ ) );
OR2_X1 _12234_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][10] ), .ZN(_04492_ ) );
OAI211_X1 _12235_ ( .A(_04492_ ), .B(_04282_ ), .C1(_04054_ ), .C2(\myreg.Reg[1][10] ), .ZN(_04493_ ) );
OR2_X1 _12236_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][10] ), .ZN(_04494_ ) );
OAI211_X1 _12237_ ( .A(_04494_ ), .B(fanout_net_37 ), .C1(_04054_ ), .C2(\myreg.Reg[3][10] ), .ZN(_04495_ ) );
NAND3_X1 _12238_ ( .A1(_04493_ ), .A2(_04495_ ), .A3(_04060_ ), .ZN(_04496_ ) );
MUX2_X1 _12239_ ( .A(\myreg.Reg[6][10] ), .B(\myreg.Reg[7][10] ), .S(fanout_net_31 ), .Z(_04497_ ) );
MUX2_X1 _12240_ ( .A(\myreg.Reg[4][10] ), .B(\myreg.Reg[5][10] ), .S(fanout_net_31 ), .Z(_04498_ ) );
MUX2_X1 _12241_ ( .A(_04497_ ), .B(_04498_ ), .S(_04065_ ), .Z(_04499_ ) );
OAI211_X1 _12242_ ( .A(_04049_ ), .B(_04496_ ), .C1(_04499_ ), .C2(_04290_ ), .ZN(_04500_ ) );
OAI211_X1 _12243_ ( .A(_04491_ ), .B(_04500_ ), .C1(_04302_ ), .C2(_02331_ ), .ZN(_04501_ ) );
OR3_X1 _12244_ ( .A1(_04095_ ), .A2(\EX_LS_result_reg [10] ), .A3(_02162_ ), .ZN(_04502_ ) );
NAND2_X1 _12245_ ( .A1(_04501_ ), .A2(_04502_ ), .ZN(_04503_ ) );
XOR2_X1 _12246_ ( .A(_02647_ ), .B(_04503_ ), .Z(_04504_ ) );
OR2_X1 _12247_ ( .A1(_04283_ ), .A2(\myreg.Reg[9][11] ), .ZN(_04505_ ) );
OAI211_X1 _12248_ ( .A(_04505_ ), .B(_04314_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[8][11] ), .ZN(_04506_ ) );
OR2_X1 _12249_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[10][11] ), .ZN(_04507_ ) );
OAI211_X1 _12250_ ( .A(_04507_ ), .B(fanout_net_37 ), .C1(_04343_ ), .C2(\myreg.Reg[11][11] ), .ZN(_04508_ ) );
NAND3_X1 _12251_ ( .A1(_04506_ ), .A2(_04060_ ), .A3(_04508_ ), .ZN(_04509_ ) );
MUX2_X1 _12252_ ( .A(\myreg.Reg[14][11] ), .B(\myreg.Reg[15][11] ), .S(fanout_net_31 ), .Z(_04510_ ) );
MUX2_X1 _12253_ ( .A(\myreg.Reg[12][11] ), .B(\myreg.Reg[13][11] ), .S(fanout_net_31 ), .Z(_04511_ ) );
MUX2_X1 _12254_ ( .A(_04510_ ), .B(_04511_ ), .S(_04065_ ), .Z(_04512_ ) );
OAI211_X1 _12255_ ( .A(fanout_net_39 ), .B(_04509_ ), .C1(_04512_ ), .C2(_04290_ ), .ZN(_04513_ ) );
NOR2_X1 _12256_ ( .A1(_04393_ ), .A2(\myreg.Reg[3][11] ), .ZN(_04514_ ) );
OAI21_X1 _12257_ ( .A(fanout_net_37 ), .B1(fanout_net_31 ), .B2(\myreg.Reg[2][11] ), .ZN(_04515_ ) );
NOR2_X1 _12258_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][11] ), .ZN(_04516_ ) );
OAI21_X1 _12259_ ( .A(_04065_ ), .B1(_04393_ ), .B2(\myreg.Reg[1][11] ), .ZN(_04517_ ) );
OAI221_X1 _12260_ ( .A(_04342_ ), .B1(_04514_ ), .B2(_04515_ ), .C1(_04516_ ), .C2(_04517_ ), .ZN(_04518_ ) );
MUX2_X1 _12261_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_32 ), .Z(_04519_ ) );
MUX2_X1 _12262_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_32 ), .Z(_04520_ ) );
MUX2_X1 _12263_ ( .A(_04519_ ), .B(_04520_ ), .S(_04065_ ), .Z(_04521_ ) );
OAI211_X1 _12264_ ( .A(_04049_ ), .B(_04518_ ), .C1(_04521_ ), .C2(_04279_ ), .ZN(_04522_ ) );
OAI211_X1 _12265_ ( .A(_04513_ ), .B(_04522_ ), .C1(_04302_ ), .C2(_02331_ ), .ZN(_04523_ ) );
OR3_X1 _12266_ ( .A1(_04095_ ), .A2(\EX_LS_result_reg [11] ), .A3(_02162_ ), .ZN(_04524_ ) );
NAND2_X1 _12267_ ( .A1(_04523_ ), .A2(_04524_ ), .ZN(_04525_ ) );
INV_X1 _12268_ ( .A(_04525_ ), .ZN(_04526_ ) );
XNOR2_X2 _12269_ ( .A(_04526_ ), .B(_02670_ ), .ZN(_04527_ ) );
AND2_X1 _12270_ ( .A1(_04504_ ), .A2(_04527_ ), .ZN(_04528_ ) );
OR2_X1 _12271_ ( .A1(_04393_ ), .A2(\myreg.Reg[3][8] ), .ZN(_04529_ ) );
OAI211_X1 _12272_ ( .A(_04529_ ), .B(fanout_net_37 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[2][8] ), .ZN(_04530_ ) );
OR2_X1 _12273_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][8] ), .ZN(_04531_ ) );
OAI211_X1 _12274_ ( .A(_04531_ ), .B(_04282_ ), .C1(_04284_ ), .C2(\myreg.Reg[1][8] ), .ZN(_04532_ ) );
NAND3_X1 _12275_ ( .A1(_04530_ ), .A2(_04290_ ), .A3(_04532_ ), .ZN(_04533_ ) );
MUX2_X1 _12276_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_32 ), .Z(_04534_ ) );
MUX2_X1 _12277_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_32 ), .Z(_04535_ ) );
MUX2_X1 _12278_ ( .A(_04534_ ), .B(_04535_ ), .S(_04282_ ), .Z(_04536_ ) );
OAI211_X1 _12279_ ( .A(_04049_ ), .B(_04533_ ), .C1(_04536_ ), .C2(_04061_ ), .ZN(_04537_ ) );
OR2_X1 _12280_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[14][8] ), .ZN(_04538_ ) );
OAI211_X1 _12281_ ( .A(_04538_ ), .B(fanout_net_37 ), .C1(_04284_ ), .C2(\myreg.Reg[15][8] ), .ZN(_04539_ ) );
OR2_X1 _12282_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][8] ), .ZN(_04540_ ) );
OAI211_X1 _12283_ ( .A(_04540_ ), .B(_04282_ ), .C1(_04284_ ), .C2(\myreg.Reg[13][8] ), .ZN(_04541_ ) );
NAND3_X1 _12284_ ( .A1(_04539_ ), .A2(_04541_ ), .A3(fanout_net_38 ), .ZN(_04542_ ) );
MUX2_X1 _12285_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_32 ), .Z(_04543_ ) );
MUX2_X1 _12286_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_32 ), .Z(_04544_ ) );
MUX2_X1 _12287_ ( .A(_04543_ ), .B(_04544_ ), .S(fanout_net_37 ), .Z(_04545_ ) );
OAI211_X1 _12288_ ( .A(fanout_net_39 ), .B(_04542_ ), .C1(_04545_ ), .C2(fanout_net_38 ), .ZN(_04546_ ) );
OAI211_X1 _12289_ ( .A(_04537_ ), .B(_04546_ ), .C1(_04096_ ), .C2(_02163_ ), .ZN(_04547_ ) );
OR3_X1 _12290_ ( .A1(_04302_ ), .A2(\EX_LS_result_reg [8] ), .A3(_02304_ ), .ZN(_04548_ ) );
NAND2_X1 _12291_ ( .A1(_04547_ ), .A2(_04548_ ), .ZN(_04549_ ) );
XOR2_X1 _12292_ ( .A(_02600_ ), .B(_04549_ ), .Z(_04550_ ) );
OR2_X1 _12293_ ( .A1(_04053_ ), .A2(\myreg.Reg[11][9] ), .ZN(_04551_ ) );
OAI211_X1 _12294_ ( .A(_04551_ ), .B(fanout_net_37 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[10][9] ), .ZN(_04552_ ) );
OR2_X1 _12295_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][9] ), .ZN(_04553_ ) );
OAI211_X1 _12296_ ( .A(_04553_ ), .B(_04389_ ), .C1(_04393_ ), .C2(\myreg.Reg[9][9] ), .ZN(_04554_ ) );
NAND3_X1 _12297_ ( .A1(_04552_ ), .A2(_04342_ ), .A3(_04554_ ), .ZN(_04555_ ) );
MUX2_X1 _12298_ ( .A(\myreg.Reg[14][9] ), .B(\myreg.Reg[15][9] ), .S(fanout_net_32 ), .Z(_04556_ ) );
MUX2_X1 _12299_ ( .A(\myreg.Reg[12][9] ), .B(\myreg.Reg[13][9] ), .S(fanout_net_32 ), .Z(_04557_ ) );
MUX2_X1 _12300_ ( .A(_04556_ ), .B(_04557_ ), .S(_04389_ ), .Z(_04558_ ) );
OAI211_X1 _12301_ ( .A(fanout_net_39 ), .B(_04555_ ), .C1(_04558_ ), .C2(_04279_ ), .ZN(_04559_ ) );
OR2_X1 _12302_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][9] ), .ZN(_04560_ ) );
OAI211_X1 _12303_ ( .A(_04560_ ), .B(_04389_ ), .C1(_04393_ ), .C2(\myreg.Reg[1][9] ), .ZN(_04561_ ) );
NOR2_X1 _12304_ ( .A1(_04343_ ), .A2(\myreg.Reg[3][9] ), .ZN(_04562_ ) );
OAI21_X1 _12305_ ( .A(fanout_net_37 ), .B1(fanout_net_32 ), .B2(\myreg.Reg[2][9] ), .ZN(_04563_ ) );
OAI211_X1 _12306_ ( .A(_04561_ ), .B(_04278_ ), .C1(_04562_ ), .C2(_04563_ ), .ZN(_04564_ ) );
MUX2_X1 _12307_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_32 ), .Z(_04565_ ) );
MUX2_X1 _12308_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_32 ), .Z(_04566_ ) );
MUX2_X1 _12309_ ( .A(_04565_ ), .B(_04566_ ), .S(_04389_ ), .Z(_04567_ ) );
OAI211_X1 _12310_ ( .A(_04048_ ), .B(_04564_ ), .C1(_04567_ ), .C2(_04279_ ), .ZN(_04568_ ) );
OAI211_X1 _12311_ ( .A(_04559_ ), .B(_04568_ ), .C1(_04095_ ), .C2(_02304_ ), .ZN(_04569_ ) );
OR3_X1 _12312_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [9] ), .A3(_02456_ ), .ZN(_04570_ ) );
NAND2_X1 _12313_ ( .A1(_04569_ ), .A2(_04570_ ), .ZN(_04571_ ) );
AND2_X1 _12314_ ( .A1(_02624_ ), .A2(_04571_ ), .ZN(_04572_ ) );
NOR2_X1 _12315_ ( .A1(_02624_ ), .A2(_04571_ ), .ZN(_04573_ ) );
NOR2_X1 _12316_ ( .A1(_04572_ ), .A2(_04573_ ), .ZN(_04574_ ) );
AND3_X1 _12317_ ( .A1(_04528_ ), .A2(_04550_ ), .A3(_04574_ ), .ZN(_04575_ ) );
INV_X1 _12318_ ( .A(_04575_ ), .ZN(_04576_ ) );
OR2_X1 _12319_ ( .A1(_04051_ ), .A2(\myreg.Reg[1][15] ), .ZN(_04577_ ) );
OAI211_X1 _12320_ ( .A(_04577_ ), .B(_04063_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[0][15] ), .ZN(_04578_ ) );
OR2_X1 _12321_ ( .A1(_04051_ ), .A2(\myreg.Reg[3][15] ), .ZN(_04579_ ) );
OAI211_X1 _12322_ ( .A(_04579_ ), .B(fanout_net_37 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[2][15] ), .ZN(_04580_ ) );
NAND3_X1 _12323_ ( .A1(_04578_ ), .A2(_04580_ ), .A3(_04058_ ), .ZN(_04581_ ) );
MUX2_X1 _12324_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_32 ), .Z(_04582_ ) );
MUX2_X1 _12325_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_32 ), .Z(_04583_ ) );
MUX2_X1 _12326_ ( .A(_04582_ ), .B(_04583_ ), .S(_04063_ ), .Z(_04584_ ) );
OAI211_X1 _12327_ ( .A(_04047_ ), .B(_04581_ ), .C1(_04584_ ), .C2(_04058_ ), .ZN(_04585_ ) );
OR2_X1 _12328_ ( .A1(_04051_ ), .A2(\myreg.Reg[15][15] ), .ZN(_04586_ ) );
OAI211_X1 _12329_ ( .A(_04586_ ), .B(fanout_net_37 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[14][15] ), .ZN(_04587_ ) );
OR2_X1 _12330_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][15] ), .ZN(_04588_ ) );
OAI211_X1 _12331_ ( .A(_04588_ ), .B(_04063_ ), .C1(_04051_ ), .C2(\myreg.Reg[13][15] ), .ZN(_04589_ ) );
NAND3_X1 _12332_ ( .A1(_04587_ ), .A2(fanout_net_38 ), .A3(_04589_ ), .ZN(_04590_ ) );
MUX2_X1 _12333_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_32 ), .Z(_04591_ ) );
MUX2_X1 _12334_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_32 ), .Z(_04592_ ) );
MUX2_X1 _12335_ ( .A(_04591_ ), .B(_04592_ ), .S(fanout_net_37 ), .Z(_04593_ ) );
OAI211_X1 _12336_ ( .A(fanout_net_39 ), .B(_04590_ ), .C1(_04593_ ), .C2(fanout_net_38 ), .ZN(_04594_ ) );
NAND2_X1 _12337_ ( .A1(_04585_ ), .A2(_04594_ ), .ZN(_04595_ ) );
OAI21_X1 _12338_ ( .A(_04595_ ), .B1(_02161_ ), .B2(_04094_ ), .ZN(_04596_ ) );
INV_X1 _12339_ ( .A(\EX_LS_result_reg [15] ), .ZN(_04597_ ) );
OR3_X1 _12340_ ( .A1(_04093_ ), .A2(_04597_ ), .A3(_02131_ ), .ZN(_04598_ ) );
AND2_X2 _12341_ ( .A1(_04596_ ), .A2(_04598_ ), .ZN(_04599_ ) );
XOR2_X1 _12342_ ( .A(_02503_ ), .B(_04599_ ), .Z(_04600_ ) );
OR2_X1 _12343_ ( .A1(_04052_ ), .A2(\myreg.Reg[1][14] ), .ZN(_04601_ ) );
OAI211_X1 _12344_ ( .A(_04601_ ), .B(_04064_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[0][14] ), .ZN(_04602_ ) );
OR2_X1 _12345_ ( .A1(_04052_ ), .A2(\myreg.Reg[3][14] ), .ZN(_04603_ ) );
OAI211_X1 _12346_ ( .A(_04603_ ), .B(fanout_net_37 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[2][14] ), .ZN(_04604_ ) );
NAND3_X1 _12347_ ( .A1(_04602_ ), .A2(_04604_ ), .A3(_04059_ ), .ZN(_04605_ ) );
MUX2_X1 _12348_ ( .A(\myreg.Reg[6][14] ), .B(\myreg.Reg[7][14] ), .S(fanout_net_32 ), .Z(_04606_ ) );
MUX2_X1 _12349_ ( .A(\myreg.Reg[4][14] ), .B(\myreg.Reg[5][14] ), .S(fanout_net_32 ), .Z(_04607_ ) );
MUX2_X1 _12350_ ( .A(_04606_ ), .B(_04607_ ), .S(_04064_ ), .Z(_04608_ ) );
OAI211_X1 _12351_ ( .A(_04047_ ), .B(_04605_ ), .C1(_04608_ ), .C2(_04278_ ), .ZN(_04609_ ) );
OR2_X1 _12352_ ( .A1(_04052_ ), .A2(\myreg.Reg[15][14] ), .ZN(_04610_ ) );
OAI211_X1 _12353_ ( .A(_04610_ ), .B(fanout_net_37 ), .C1(fanout_net_33 ), .C2(\myreg.Reg[14][14] ), .ZN(_04611_ ) );
OR2_X1 _12354_ ( .A1(_04052_ ), .A2(\myreg.Reg[13][14] ), .ZN(_04612_ ) );
OAI211_X1 _12355_ ( .A(_04612_ ), .B(_04064_ ), .C1(fanout_net_33 ), .C2(\myreg.Reg[12][14] ), .ZN(_04613_ ) );
NAND3_X1 _12356_ ( .A1(_04611_ ), .A2(_04613_ ), .A3(fanout_net_38 ), .ZN(_04614_ ) );
MUX2_X1 _12357_ ( .A(\myreg.Reg[8][14] ), .B(\myreg.Reg[9][14] ), .S(fanout_net_33 ), .Z(_04615_ ) );
MUX2_X1 _12358_ ( .A(\myreg.Reg[10][14] ), .B(\myreg.Reg[11][14] ), .S(fanout_net_33 ), .Z(_04616_ ) );
MUX2_X1 _12359_ ( .A(_04615_ ), .B(_04616_ ), .S(fanout_net_37 ), .Z(_04617_ ) );
OAI211_X1 _12360_ ( .A(fanout_net_39 ), .B(_04614_ ), .C1(_04617_ ), .C2(fanout_net_38 ), .ZN(_04618_ ) );
OAI211_X1 _12361_ ( .A(_04609_ ), .B(_04618_ ), .C1(_04094_ ), .C2(_02303_ ), .ZN(_04619_ ) );
OR3_X1 _12362_ ( .A1(_04094_ ), .A2(\EX_LS_result_reg [14] ), .A3(_02161_ ), .ZN(_04620_ ) );
NAND2_X1 _12363_ ( .A1(_04619_ ), .A2(_04620_ ), .ZN(_04621_ ) );
INV_X1 _12364_ ( .A(_04621_ ), .ZN(_04622_ ) );
XNOR2_X1 _12365_ ( .A(_04622_ ), .B(_02526_ ), .ZN(_04623_ ) );
AND2_X1 _12366_ ( .A1(_04600_ ), .A2(_04623_ ), .ZN(_04624_ ) );
NOR2_X1 _12367_ ( .A1(_04283_ ), .A2(\myreg.Reg[3][12] ), .ZN(_04625_ ) );
OAI21_X1 _12368_ ( .A(fanout_net_37 ), .B1(fanout_net_33 ), .B2(\myreg.Reg[2][12] ), .ZN(_04626_ ) );
NOR2_X1 _12369_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[0][12] ), .ZN(_04627_ ) );
OAI21_X1 _12370_ ( .A(_04281_ ), .B1(_04275_ ), .B2(\myreg.Reg[1][12] ), .ZN(_04628_ ) );
OAI221_X1 _12371_ ( .A(_04278_ ), .B1(_04625_ ), .B2(_04626_ ), .C1(_04627_ ), .C2(_04628_ ), .ZN(_04629_ ) );
MUX2_X1 _12372_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_33 ), .Z(_04630_ ) );
MUX2_X1 _12373_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_33 ), .Z(_04631_ ) );
MUX2_X1 _12374_ ( .A(_04630_ ), .B(_04631_ ), .S(_04392_ ), .Z(_04632_ ) );
OAI211_X1 _12375_ ( .A(_04048_ ), .B(_04629_ ), .C1(_04632_ ), .C2(_04060_ ), .ZN(_04633_ ) );
OR2_X1 _12376_ ( .A1(_04274_ ), .A2(\myreg.Reg[11][12] ), .ZN(_04634_ ) );
OAI211_X1 _12377_ ( .A(_04634_ ), .B(fanout_net_37 ), .C1(fanout_net_33 ), .C2(\myreg.Reg[10][12] ), .ZN(_04635_ ) );
OR2_X1 _12378_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[8][12] ), .ZN(_04636_ ) );
OAI211_X1 _12379_ ( .A(_04636_ ), .B(_04392_ ), .C1(_04275_ ), .C2(\myreg.Reg[9][12] ), .ZN(_04637_ ) );
NAND3_X1 _12380_ ( .A1(_04635_ ), .A2(_04278_ ), .A3(_04637_ ), .ZN(_04638_ ) );
MUX2_X1 _12381_ ( .A(\myreg.Reg[14][12] ), .B(\myreg.Reg[15][12] ), .S(fanout_net_33 ), .Z(_04639_ ) );
MUX2_X1 _12382_ ( .A(\myreg.Reg[12][12] ), .B(\myreg.Reg[13][12] ), .S(fanout_net_33 ), .Z(_04640_ ) );
MUX2_X1 _12383_ ( .A(_04639_ ), .B(_04640_ ), .S(_04281_ ), .Z(_04641_ ) );
OAI211_X1 _12384_ ( .A(fanout_net_39 ), .B(_04638_ ), .C1(_04641_ ), .C2(_04060_ ), .ZN(_04642_ ) );
OAI211_X1 _12385_ ( .A(_04633_ ), .B(_04642_ ), .C1(_02304_ ), .C2(_04301_ ), .ZN(_04643_ ) );
OR3_X1 _12386_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [12] ), .A3(_02303_ ), .ZN(_04644_ ) );
NAND2_X1 _12387_ ( .A1(_04643_ ), .A2(_04644_ ), .ZN(_04645_ ) );
INV_X1 _12388_ ( .A(_04645_ ), .ZN(_04646_ ) );
XNOR2_X1 _12389_ ( .A(_04646_ ), .B(_02574_ ), .ZN(_04647_ ) );
OR3_X1 _12390_ ( .A1(_04094_ ), .A2(\EX_LS_result_reg [13] ), .A3(_02161_ ), .ZN(_04648_ ) );
OR2_X1 _12391_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[0][13] ), .ZN(_04649_ ) );
OAI211_X1 _12392_ ( .A(_04649_ ), .B(_04281_ ), .C1(_04283_ ), .C2(\myreg.Reg[1][13] ), .ZN(_04650_ ) );
OR2_X1 _12393_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[2][13] ), .ZN(_04651_ ) );
OAI211_X1 _12394_ ( .A(_04651_ ), .B(fanout_net_37 ), .C1(_04283_ ), .C2(\myreg.Reg[3][13] ), .ZN(_04652_ ) );
NAND3_X1 _12395_ ( .A1(_04650_ ), .A2(_04652_ ), .A3(_04059_ ), .ZN(_04653_ ) );
MUX2_X1 _12396_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_33 ), .Z(_04654_ ) );
MUX2_X1 _12397_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_33 ), .Z(_04655_ ) );
MUX2_X1 _12398_ ( .A(_04654_ ), .B(_04655_ ), .S(_04064_ ), .Z(_04656_ ) );
OAI211_X1 _12399_ ( .A(_04048_ ), .B(_04653_ ), .C1(_04656_ ), .C2(_04278_ ), .ZN(_04657_ ) );
OR2_X1 _12400_ ( .A1(_04052_ ), .A2(\myreg.Reg[15][13] ), .ZN(_04658_ ) );
OAI211_X1 _12401_ ( .A(_04658_ ), .B(fanout_net_37 ), .C1(fanout_net_33 ), .C2(\myreg.Reg[14][13] ), .ZN(_04659_ ) );
OR2_X1 _12402_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[12][13] ), .ZN(_04660_ ) );
OAI211_X1 _12403_ ( .A(_04660_ ), .B(_04064_ ), .C1(_04053_ ), .C2(\myreg.Reg[13][13] ), .ZN(_04661_ ) );
NAND3_X1 _12404_ ( .A1(_04659_ ), .A2(fanout_net_38 ), .A3(_04661_ ), .ZN(_04662_ ) );
MUX2_X1 _12405_ ( .A(\myreg.Reg[8][13] ), .B(\myreg.Reg[9][13] ), .S(fanout_net_33 ), .Z(_04663_ ) );
MUX2_X1 _12406_ ( .A(\myreg.Reg[10][13] ), .B(\myreg.Reg[11][13] ), .S(fanout_net_33 ), .Z(_04664_ ) );
MUX2_X1 _12407_ ( .A(_04663_ ), .B(_04664_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04665_ ) );
OAI211_X1 _12408_ ( .A(fanout_net_39 ), .B(_04662_ ), .C1(_04665_ ), .C2(fanout_net_38 ), .ZN(_04666_ ) );
OAI211_X1 _12409_ ( .A(_04657_ ), .B(_04666_ ), .C1(_04301_ ), .C2(_02456_ ), .ZN(_04667_ ) );
NAND2_X1 _12410_ ( .A1(_04648_ ), .A2(_04667_ ), .ZN(_04668_ ) );
AND2_X1 _12411_ ( .A1(_02551_ ), .A2(_04668_ ), .ZN(_04669_ ) );
NOR2_X1 _12412_ ( .A1(_02552_ ), .A2(_04668_ ), .ZN(_04670_ ) );
NOR2_X1 _12413_ ( .A1(_04669_ ), .A2(_04670_ ), .ZN(_04671_ ) );
NAND3_X1 _12414_ ( .A1(_04624_ ), .A2(_04647_ ), .A3(_04671_ ), .ZN(_04672_ ) );
NOR2_X1 _12415_ ( .A1(_04576_ ), .A2(_04672_ ), .ZN(_04673_ ) );
NAND3_X1 _12416_ ( .A1(_04273_ ), .A2(_04482_ ), .A3(_04673_ ), .ZN(_04674_ ) );
OR2_X1 _12417_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04675_ ) );
OAI211_X1 _12418_ ( .A(_04675_ ), .B(_04392_ ), .C1(_04275_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04676_ ) );
OR2_X1 _12419_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04677_ ) );
OAI211_X1 _12420_ ( .A(_04677_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04275_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04678_ ) );
NAND3_X1 _12421_ ( .A1(_04676_ ), .A2(_04678_ ), .A3(_04278_ ), .ZN(_04679_ ) );
MUX2_X1 _12422_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04680_ ) );
MUX2_X1 _12423_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04681_ ) );
MUX2_X1 _12424_ ( .A(_04680_ ), .B(_04681_ ), .S(_04281_ ), .Z(_04682_ ) );
OAI211_X1 _12425_ ( .A(_04048_ ), .B(_04679_ ), .C1(_04682_ ), .C2(_04342_ ), .ZN(_04683_ ) );
OR2_X1 _12426_ ( .A1(_04274_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04684_ ) );
OAI211_X1 _12427_ ( .A(_04684_ ), .B(_04281_ ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04685_ ) );
OR2_X1 _12428_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04686_ ) );
OAI211_X1 _12429_ ( .A(_04686_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04283_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04687_ ) );
NAND3_X1 _12430_ ( .A1(_04685_ ), .A2(fanout_net_38 ), .A3(_04687_ ), .ZN(_04688_ ) );
MUX2_X1 _12431_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04689_ ) );
MUX2_X1 _12432_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04690_ ) );
MUX2_X1 _12433_ ( .A(_04689_ ), .B(_04690_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04691_ ) );
OAI211_X1 _12434_ ( .A(fanout_net_39 ), .B(_04688_ ), .C1(_04691_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04692_ ) );
AOI21_X1 _12435_ ( .A(_04099_ ), .B1(_04683_ ), .B2(_04692_ ), .ZN(_04693_ ) );
AND2_X1 _12436_ ( .A1(_04099_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04694_ ) );
NOR2_X1 _12437_ ( .A1(_04693_ ), .A2(_04694_ ), .ZN(_04695_ ) );
XNOR2_X1 _12438_ ( .A(_04695_ ), .B(_02766_ ), .ZN(_04696_ ) );
OR2_X1 _12439_ ( .A1(_04053_ ), .A2(\myreg.Reg[1][4] ), .ZN(_04697_ ) );
OAI211_X1 _12440_ ( .A(_04697_ ), .B(_04314_ ), .C1(fanout_net_33 ), .C2(\myreg.Reg[0][4] ), .ZN(_04698_ ) );
OR2_X1 _12441_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[2][4] ), .ZN(_04699_ ) );
OAI211_X1 _12442_ ( .A(_04699_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04343_ ), .C2(\myreg.Reg[3][4] ), .ZN(_04700_ ) );
NAND3_X1 _12443_ ( .A1(_04698_ ), .A2(_04342_ ), .A3(_04700_ ), .ZN(_04701_ ) );
MUX2_X1 _12444_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_34 ), .Z(_04702_ ) );
MUX2_X1 _12445_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_34 ), .Z(_04703_ ) );
MUX2_X1 _12446_ ( .A(_04702_ ), .B(_04703_ ), .S(_04389_ ), .Z(_04704_ ) );
OAI211_X1 _12447_ ( .A(_04049_ ), .B(_04701_ ), .C1(_04704_ ), .C2(_04279_ ), .ZN(_04705_ ) );
OR2_X1 _12448_ ( .A1(_04053_ ), .A2(\myreg.Reg[13][4] ), .ZN(_04706_ ) );
OAI211_X1 _12449_ ( .A(_04706_ ), .B(_04314_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[12][4] ), .ZN(_04707_ ) );
OR2_X1 _12450_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[14][4] ), .ZN(_04708_ ) );
OAI211_X1 _12451_ ( .A(_04708_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04343_ ), .C2(\myreg.Reg[15][4] ), .ZN(_04709_ ) );
NAND3_X1 _12452_ ( .A1(_04707_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04709_ ), .ZN(_04710_ ) );
MUX2_X1 _12453_ ( .A(\myreg.Reg[8][4] ), .B(\myreg.Reg[9][4] ), .S(fanout_net_34 ), .Z(_04711_ ) );
MUX2_X1 _12454_ ( .A(\myreg.Reg[10][4] ), .B(\myreg.Reg[11][4] ), .S(fanout_net_34 ), .Z(_04712_ ) );
MUX2_X1 _12455_ ( .A(_04711_ ), .B(_04712_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04713_ ) );
OAI211_X1 _12456_ ( .A(fanout_net_39 ), .B(_04710_ ), .C1(_04713_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04714_ ) );
OAI211_X1 _12457_ ( .A(_04705_ ), .B(_04714_ ), .C1(_04302_ ), .C2(_02331_ ), .ZN(_04715_ ) );
OR3_X1 _12458_ ( .A1(_04095_ ), .A2(\EX_LS_result_reg [4] ), .A3(_02456_ ), .ZN(_04716_ ) );
NAND2_X1 _12459_ ( .A1(_04715_ ), .A2(_04716_ ), .ZN(_04717_ ) );
INV_X1 _12460_ ( .A(_04717_ ), .ZN(_04718_ ) );
XNOR2_X1 _12461_ ( .A(_04718_ ), .B(_02864_ ), .ZN(_04719_ ) );
NOR2_X1 _12462_ ( .A1(_04283_ ), .A2(\myreg.Reg[11][2] ), .ZN(_04720_ ) );
OAI21_X1 _12463_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_34 ), .B2(\myreg.Reg[10][2] ), .ZN(_04721_ ) );
NOR2_X1 _12464_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[8][2] ), .ZN(_04722_ ) );
OAI21_X1 _12465_ ( .A(_04281_ ), .B1(_04283_ ), .B2(\myreg.Reg[9][2] ), .ZN(_04723_ ) );
OAI221_X1 _12466_ ( .A(_04059_ ), .B1(_04720_ ), .B2(_04721_ ), .C1(_04722_ ), .C2(_04723_ ), .ZN(_04724_ ) );
MUX2_X1 _12467_ ( .A(\myreg.Reg[12][2] ), .B(\myreg.Reg[13][2] ), .S(fanout_net_34 ), .Z(_04725_ ) );
MUX2_X1 _12468_ ( .A(\myreg.Reg[14][2] ), .B(\myreg.Reg[15][2] ), .S(fanout_net_34 ), .Z(_04726_ ) );
MUX2_X1 _12469_ ( .A(_04725_ ), .B(_04726_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04727_ ) );
OAI211_X1 _12470_ ( .A(fanout_net_39 ), .B(_04724_ ), .C1(_04727_ ), .C2(_04342_ ), .ZN(_04728_ ) );
OR2_X1 _12471_ ( .A1(_04274_ ), .A2(\myreg.Reg[7][2] ), .ZN(_04729_ ) );
OAI211_X1 _12472_ ( .A(_04729_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_34 ), .C2(\myreg.Reg[6][2] ), .ZN(_04730_ ) );
OR2_X1 _12473_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[4][2] ), .ZN(_04731_ ) );
OAI211_X1 _12474_ ( .A(_04731_ ), .B(_04281_ ), .C1(_04283_ ), .C2(\myreg.Reg[5][2] ), .ZN(_04732_ ) );
NAND3_X1 _12475_ ( .A1(_04730_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04732_ ), .ZN(_04733_ ) );
MUX2_X1 _12476_ ( .A(\myreg.Reg[2][2] ), .B(\myreg.Reg[3][2] ), .S(fanout_net_34 ), .Z(_04734_ ) );
MUX2_X1 _12477_ ( .A(\myreg.Reg[0][2] ), .B(\myreg.Reg[1][2] ), .S(fanout_net_34 ), .Z(_04735_ ) );
MUX2_X1 _12478_ ( .A(_04734_ ), .B(_04735_ ), .S(_04281_ ), .Z(_04736_ ) );
OAI211_X1 _12479_ ( .A(_04048_ ), .B(_04733_ ), .C1(_04736_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04737_ ) );
OAI211_X1 _12480_ ( .A(_04728_ ), .B(_04737_ ), .C1(_02162_ ), .C2(_04301_ ), .ZN(_04738_ ) );
OR3_X1 _12481_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [2] ), .A3(_02303_ ), .ZN(_04739_ ) );
NAND2_X1 _12482_ ( .A1(_04738_ ), .A2(_04739_ ), .ZN(_04740_ ) );
INV_X1 _12483_ ( .A(_04740_ ), .ZN(_04741_ ) );
XNOR2_X1 _12484_ ( .A(_04741_ ), .B(_02695_ ), .ZN(_04742_ ) );
NAND2_X2 _12485_ ( .A1(_02739_ ), .A2(_02740_ ), .ZN(_04743_ ) );
OR2_X1 _12486_ ( .A1(_04052_ ), .A2(\myreg.Reg[9][0] ), .ZN(_04744_ ) );
OAI211_X1 _12487_ ( .A(_04744_ ), .B(_04064_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[8][0] ), .ZN(_04745_ ) );
OR2_X1 _12488_ ( .A1(_04052_ ), .A2(\myreg.Reg[11][0] ), .ZN(_04746_ ) );
OAI211_X1 _12489_ ( .A(_04746_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_34 ), .C2(\myreg.Reg[10][0] ), .ZN(_04747_ ) );
NAND3_X1 _12490_ ( .A1(_04745_ ), .A2(_04747_ ), .A3(_04059_ ), .ZN(_04748_ ) );
MUX2_X1 _12491_ ( .A(\myreg.Reg[14][0] ), .B(\myreg.Reg[15][0] ), .S(fanout_net_34 ), .Z(_04749_ ) );
MUX2_X1 _12492_ ( .A(\myreg.Reg[12][0] ), .B(\myreg.Reg[13][0] ), .S(fanout_net_34 ), .Z(_04750_ ) );
MUX2_X1 _12493_ ( .A(_04749_ ), .B(_04750_ ), .S(_04064_ ), .Z(_04751_ ) );
OAI211_X1 _12494_ ( .A(fanout_net_39 ), .B(_04748_ ), .C1(_04751_ ), .C2(_04059_ ), .ZN(_04752_ ) );
NOR2_X1 _12495_ ( .A1(_04052_ ), .A2(\myreg.Reg[3][0] ), .ZN(_04753_ ) );
OAI21_X1 _12496_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_34 ), .B2(\myreg.Reg[2][0] ), .ZN(_04754_ ) );
NOR2_X1 _12497_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[0][0] ), .ZN(_04755_ ) );
OAI21_X1 _12498_ ( .A(_04063_ ), .B1(_04274_ ), .B2(\myreg.Reg[1][0] ), .ZN(_04756_ ) );
OAI221_X1 _12499_ ( .A(_04059_ ), .B1(_04753_ ), .B2(_04754_ ), .C1(_04755_ ), .C2(_04756_ ), .ZN(_04757_ ) );
MUX2_X1 _12500_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_34 ), .Z(_04758_ ) );
MUX2_X1 _12501_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_34 ), .Z(_04759_ ) );
MUX2_X1 _12502_ ( .A(_04758_ ), .B(_04759_ ), .S(_04063_ ), .Z(_04760_ ) );
OAI211_X1 _12503_ ( .A(_04047_ ), .B(_04757_ ), .C1(_04760_ ), .C2(_04059_ ), .ZN(_04761_ ) );
OAI211_X1 _12504_ ( .A(_04752_ ), .B(_04761_ ), .C1(_04094_ ), .C2(_02303_ ), .ZN(_04762_ ) );
OR3_X1 _12505_ ( .A1(_04094_ ), .A2(\EX_LS_result_reg [0] ), .A3(_02161_ ), .ZN(_04763_ ) );
NAND2_X1 _12506_ ( .A1(_04762_ ), .A2(_04763_ ), .ZN(_04764_ ) );
NAND2_X1 _12507_ ( .A1(_04743_ ), .A2(_04764_ ), .ZN(_04765_ ) );
AND4_X1 _12508_ ( .A1(_04696_ ), .A2(_04719_ ), .A3(_04742_ ), .A4(_04765_ ), .ZN(_04766_ ) );
OR2_X1 _12509_ ( .A1(_04051_ ), .A2(\myreg.Reg[1][1] ), .ZN(_04767_ ) );
OAI211_X1 _12510_ ( .A(_04767_ ), .B(_04063_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[0][1] ), .ZN(_04768_ ) );
OR2_X1 _12511_ ( .A1(_04051_ ), .A2(\myreg.Reg[3][1] ), .ZN(_04769_ ) );
OAI211_X1 _12512_ ( .A(_04769_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_34 ), .C2(\myreg.Reg[2][1] ), .ZN(_04770_ ) );
NAND3_X1 _12513_ ( .A1(_04768_ ), .A2(_04770_ ), .A3(_04058_ ), .ZN(_04771_ ) );
MUX2_X1 _12514_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(fanout_net_34 ), .Z(_04772_ ) );
MUX2_X1 _12515_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(fanout_net_34 ), .Z(_04773_ ) );
MUX2_X1 _12516_ ( .A(_04772_ ), .B(_04773_ ), .S(_04063_ ), .Z(_04774_ ) );
OAI211_X1 _12517_ ( .A(_04047_ ), .B(_04771_ ), .C1(_04774_ ), .C2(_04059_ ), .ZN(_04775_ ) );
OR2_X1 _12518_ ( .A1(_04051_ ), .A2(\myreg.Reg[15][1] ), .ZN(_04776_ ) );
OAI211_X1 _12519_ ( .A(_04776_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_34 ), .C2(\myreg.Reg[14][1] ), .ZN(_04777_ ) );
OR2_X1 _12520_ ( .A1(_04051_ ), .A2(\myreg.Reg[13][1] ), .ZN(_04778_ ) );
OAI211_X1 _12521_ ( .A(_04778_ ), .B(_04063_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[12][1] ), .ZN(_04779_ ) );
NAND3_X1 _12522_ ( .A1(_04777_ ), .A2(_04779_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04780_ ) );
MUX2_X1 _12523_ ( .A(\myreg.Reg[8][1] ), .B(\myreg.Reg[9][1] ), .S(fanout_net_34 ), .Z(_04781_ ) );
MUX2_X1 _12524_ ( .A(\myreg.Reg[10][1] ), .B(\myreg.Reg[11][1] ), .S(fanout_net_34 ), .Z(_04782_ ) );
MUX2_X1 _12525_ ( .A(_04781_ ), .B(_04782_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04783_ ) );
OAI211_X1 _12526_ ( .A(fanout_net_39 ), .B(_04780_ ), .C1(_04783_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04784_ ) );
OAI211_X1 _12527_ ( .A(_04775_ ), .B(_04784_ ), .C1(_04094_ ), .C2(_02161_ ), .ZN(_04785_ ) );
OR3_X1 _12528_ ( .A1(_04093_ ), .A2(\EX_LS_result_reg [1] ), .A3(_02131_ ), .ZN(_04786_ ) );
NAND2_X1 _12529_ ( .A1(_04785_ ), .A2(_04786_ ), .ZN(_04787_ ) );
XOR2_X1 _12530_ ( .A(_02717_ ), .B(_04787_ ), .Z(_04788_ ) );
NOR2_X1 _12531_ ( .A1(_04743_ ), .A2(_04764_ ), .ZN(_04789_ ) );
INV_X1 _12532_ ( .A(_04789_ ), .ZN(_04790_ ) );
AND2_X1 _12533_ ( .A1(_04788_ ), .A2(_04790_ ), .ZN(_04791_ ) );
AND2_X1 _12534_ ( .A1(_04766_ ), .A2(_04791_ ), .ZN(_04792_ ) );
OR2_X1 _12535_ ( .A1(_04274_ ), .A2(\myreg.Reg[5][7] ), .ZN(_04793_ ) );
OAI211_X1 _12536_ ( .A(_04793_ ), .B(_04392_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[4][7] ), .ZN(_04794_ ) );
OR2_X1 _12537_ ( .A1(_04274_ ), .A2(\myreg.Reg[7][7] ), .ZN(_04795_ ) );
OAI211_X1 _12538_ ( .A(_04795_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_35 ), .C2(\myreg.Reg[6][7] ), .ZN(_04796_ ) );
NAND3_X1 _12539_ ( .A1(_04794_ ), .A2(_04796_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04797_ ) );
MUX2_X1 _12540_ ( .A(\myreg.Reg[2][7] ), .B(\myreg.Reg[3][7] ), .S(fanout_net_35 ), .Z(_04798_ ) );
MUX2_X1 _12541_ ( .A(\myreg.Reg[0][7] ), .B(\myreg.Reg[1][7] ), .S(fanout_net_35 ), .Z(_04799_ ) );
MUX2_X1 _12542_ ( .A(_04798_ ), .B(_04799_ ), .S(_04392_ ), .Z(_04800_ ) );
OAI211_X1 _12543_ ( .A(_04048_ ), .B(_04797_ ), .C1(_04800_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04801_ ) );
NOR2_X1 _12544_ ( .A1(_04275_ ), .A2(\myreg.Reg[11][7] ), .ZN(_04802_ ) );
OAI21_X1 _12545_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_35 ), .B2(\myreg.Reg[10][7] ), .ZN(_04803_ ) );
NOR2_X1 _12546_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[8][7] ), .ZN(_04804_ ) );
OAI21_X1 _12547_ ( .A(_04392_ ), .B1(_04275_ ), .B2(\myreg.Reg[9][7] ), .ZN(_04805_ ) );
OAI221_X1 _12548_ ( .A(_04278_ ), .B1(_04802_ ), .B2(_04803_ ), .C1(_04804_ ), .C2(_04805_ ), .ZN(_04806_ ) );
MUX2_X1 _12549_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_35 ), .Z(_04807_ ) );
MUX2_X1 _12550_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_35 ), .Z(_04808_ ) );
MUX2_X1 _12551_ ( .A(_04807_ ), .B(_04808_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04809_ ) );
OAI211_X1 _12552_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04806_ ), .C1(_04809_ ), .C2(_04060_ ), .ZN(_04810_ ) );
OAI211_X1 _12553_ ( .A(_04801_ ), .B(_04810_ ), .C1(_04095_ ), .C2(_02162_ ), .ZN(_04811_ ) );
OR3_X1 _12554_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [7] ), .A3(_02303_ ), .ZN(_04812_ ) );
NAND2_X1 _12555_ ( .A1(_04811_ ), .A2(_04812_ ), .ZN(_04813_ ) );
INV_X1 _12556_ ( .A(_04813_ ), .ZN(_04814_ ) );
XNOR2_X1 _12557_ ( .A(_04814_ ), .B(_02816_ ), .ZN(_04815_ ) );
OR2_X1 _12558_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][6] ), .ZN(_04816_ ) );
OAI211_X1 _12559_ ( .A(_04816_ ), .B(_04314_ ), .C1(_04343_ ), .C2(\myreg.Reg[1][6] ), .ZN(_04817_ ) );
OR2_X1 _12560_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][6] ), .ZN(_04818_ ) );
OAI211_X1 _12561_ ( .A(_04818_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04343_ ), .C2(\myreg.Reg[3][6] ), .ZN(_04819_ ) );
NAND3_X1 _12562_ ( .A1(_04817_ ), .A2(_04819_ ), .A3(_04342_ ), .ZN(_04820_ ) );
MUX2_X1 _12563_ ( .A(\myreg.Reg[6][6] ), .B(\myreg.Reg[7][6] ), .S(fanout_net_35 ), .Z(_04821_ ) );
MUX2_X1 _12564_ ( .A(\myreg.Reg[4][6] ), .B(\myreg.Reg[5][6] ), .S(fanout_net_35 ), .Z(_04822_ ) );
MUX2_X1 _12565_ ( .A(_04821_ ), .B(_04822_ ), .S(_04389_ ), .Z(_04823_ ) );
OAI211_X1 _12566_ ( .A(_04049_ ), .B(_04820_ ), .C1(_04823_ ), .C2(_04279_ ), .ZN(_04824_ ) );
OR2_X1 _12567_ ( .A1(_04053_ ), .A2(\myreg.Reg[13][6] ), .ZN(_04825_ ) );
OAI211_X1 _12568_ ( .A(_04825_ ), .B(_04314_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[12][6] ), .ZN(_04826_ ) );
OR2_X1 _12569_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[14][6] ), .ZN(_04827_ ) );
OAI211_X1 _12570_ ( .A(_04827_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04343_ ), .C2(\myreg.Reg[15][6] ), .ZN(_04828_ ) );
NAND3_X1 _12571_ ( .A1(_04826_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04828_ ), .ZN(_04829_ ) );
MUX2_X1 _12572_ ( .A(\myreg.Reg[8][6] ), .B(\myreg.Reg[9][6] ), .S(fanout_net_35 ), .Z(_04830_ ) );
MUX2_X1 _12573_ ( .A(\myreg.Reg[10][6] ), .B(\myreg.Reg[11][6] ), .S(fanout_net_35 ), .Z(_04831_ ) );
MUX2_X1 _12574_ ( .A(_04830_ ), .B(_04831_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04832_ ) );
OAI211_X1 _12575_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04829_ ), .C1(_04832_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04833_ ) );
OAI211_X1 _12576_ ( .A(_04824_ ), .B(_04833_ ), .C1(_04302_ ), .C2(_02331_ ), .ZN(_04834_ ) );
OR3_X1 _12577_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [6] ), .A3(_02456_ ), .ZN(_04835_ ) );
NAND2_X1 _12578_ ( .A1(_04834_ ), .A2(_04835_ ), .ZN(_04836_ ) );
INV_X1 _12579_ ( .A(_04836_ ), .ZN(_04837_ ) );
XNOR2_X1 _12580_ ( .A(_04837_ ), .B(_02792_ ), .ZN(_04838_ ) );
AND2_X1 _12581_ ( .A1(_04815_ ), .A2(_04838_ ), .ZN(_04839_ ) );
OR2_X1 _12582_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04840_ ) );
OAI211_X1 _12583_ ( .A(_04840_ ), .B(_04392_ ), .C1(_04393_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04841_ ) );
NAND2_X1 _12584_ ( .A1(_02822_ ), .A2(fanout_net_35 ), .ZN(_04842_ ) );
OAI211_X1 _12585_ ( .A(_04842_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04843_ ) );
NAND3_X1 _12586_ ( .A1(_04841_ ), .A2(_04843_ ), .A3(_04278_ ), .ZN(_04844_ ) );
MUX2_X1 _12587_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04845_ ) );
MUX2_X1 _12588_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04846_ ) );
MUX2_X1 _12589_ ( .A(_04845_ ), .B(_04846_ ), .S(_04392_ ), .Z(_04847_ ) );
OAI211_X1 _12590_ ( .A(_04048_ ), .B(_04844_ ), .C1(_04847_ ), .C2(_04060_ ), .ZN(_04848_ ) );
OR2_X1 _12591_ ( .A1(_04274_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04849_ ) );
OAI211_X1 _12592_ ( .A(_04849_ ), .B(_04392_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04850_ ) );
OR2_X1 _12593_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04851_ ) );
OAI211_X1 _12594_ ( .A(_04851_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04275_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04852_ ) );
NAND3_X1 _12595_ ( .A1(_04850_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04852_ ), .ZN(_04853_ ) );
MUX2_X1 _12596_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04854_ ) );
MUX2_X1 _12597_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04855_ ) );
MUX2_X1 _12598_ ( .A(_04854_ ), .B(_04855_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04856_ ) );
OAI211_X1 _12599_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04853_ ), .C1(_04856_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04857_ ) );
AOI21_X1 _12600_ ( .A(_04099_ ), .B1(_04848_ ), .B2(_04857_ ), .ZN(_04858_ ) );
AND2_X1 _12601_ ( .A1(_04099_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04859_ ) );
NOR2_X2 _12602_ ( .A1(_04858_ ), .A2(_04859_ ), .ZN(_04860_ ) );
XNOR2_X1 _12603_ ( .A(_02841_ ), .B(_04860_ ), .ZN(_04861_ ) );
NAND3_X1 _12604_ ( .A1(_04792_ ), .A2(_04839_ ), .A3(_04861_ ), .ZN(_04862_ ) );
NOR2_X1 _12605_ ( .A1(_04674_ ), .A2(_04862_ ), .ZN(_04863_ ) );
INV_X1 _12606_ ( .A(_04863_ ), .ZN(_04864_ ) );
NOR2_X1 _12607_ ( .A1(_03886_ ), .A2(\ID_EX_typ [1] ), .ZN(_04865_ ) );
AND2_X2 _12608_ ( .A1(_04865_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04866_ ) );
INV_X1 _12609_ ( .A(\ID_EX_typ [1] ), .ZN(_04867_ ) );
NOR2_X1 _12610_ ( .A1(_04867_ ), .A2(fanout_net_4 ), .ZN(_04868_ ) );
INV_X1 _12611_ ( .A(\ID_EX_typ [2] ), .ZN(_04869_ ) );
AND2_X2 _12612_ ( .A1(_04868_ ), .A2(_04869_ ), .ZN(_04870_ ) );
INV_X2 _12613_ ( .A(_04870_ ), .ZN(_04871_ ) );
AND2_X1 _12614_ ( .A1(_04045_ ), .A2(\ID_EX_typ [2] ), .ZN(_04872_ ) );
INV_X1 _12615_ ( .A(_04872_ ), .ZN(_04873_ ) );
OR2_X1 _12616_ ( .A1(_04101_ ), .A2(fanout_net_5 ), .ZN(_04874_ ) );
NAND2_X1 _12617_ ( .A1(fanout_net_5 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04875_ ) );
AND2_X2 _12618_ ( .A1(_04874_ ), .A2(_04875_ ), .ZN(_04876_ ) );
XNOR2_X1 _12619_ ( .A(_04876_ ), .B(_02172_ ), .ZN(_04877_ ) );
INV_X1 _12620_ ( .A(_03004_ ), .ZN(_04878_ ) );
INV_X1 _12621_ ( .A(fanout_net_5 ), .ZN(_04879_ ) );
BUF_X2 _12622_ ( .A(_04879_ ), .Z(_04880_ ) );
BUF_X2 _12623_ ( .A(_04880_ ), .Z(_04881_ ) );
NAND3_X1 _12624_ ( .A1(_04125_ ), .A2(_04126_ ), .A3(_04881_ ), .ZN(_04882_ ) );
INV_X1 _12625_ ( .A(\ID_EX_imm [31] ), .ZN(_04883_ ) );
NAND2_X1 _12626_ ( .A1(_04883_ ), .A2(fanout_net_5 ), .ZN(_04884_ ) );
NAND2_X1 _12627_ ( .A1(_04882_ ), .A2(_04884_ ), .ZN(_04885_ ) );
NAND2_X1 _12628_ ( .A1(_04878_ ), .A2(_04885_ ), .ZN(_04886_ ) );
NAND3_X1 _12629_ ( .A1(_03004_ ), .A2(_04882_ ), .A3(_04884_ ), .ZN(_04887_ ) );
NAND2_X1 _12630_ ( .A1(_04886_ ), .A2(_04887_ ), .ZN(_04888_ ) );
INV_X1 _12631_ ( .A(_04888_ ), .ZN(_04889_ ) );
NOR2_X1 _12632_ ( .A1(_04877_ ), .A2(_04889_ ), .ZN(_04890_ ) );
NAND2_X1 _12633_ ( .A1(_04173_ ), .A2(_04881_ ), .ZN(_04891_ ) );
NAND2_X1 _12634_ ( .A1(_02978_ ), .A2(fanout_net_5 ), .ZN(_04892_ ) );
NAND2_X1 _12635_ ( .A1(_04891_ ), .A2(_04892_ ), .ZN(_04893_ ) );
INV_X1 _12636_ ( .A(_02199_ ), .ZN(_04894_ ) );
XNOR2_X1 _12637_ ( .A(_04893_ ), .B(_04894_ ), .ZN(_04895_ ) );
INV_X1 _12638_ ( .A(_04895_ ), .ZN(_04896_ ) );
OR2_X1 _12639_ ( .A1(_04151_ ), .A2(fanout_net_5 ), .ZN(_04897_ ) );
NAND2_X1 _12640_ ( .A1(fanout_net_5 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04898_ ) );
AND2_X1 _12641_ ( .A1(_04897_ ), .A2(_04898_ ), .ZN(_04899_ ) );
XNOR2_X1 _12642_ ( .A(_04899_ ), .B(_02976_ ), .ZN(_04900_ ) );
INV_X1 _12643_ ( .A(_04900_ ), .ZN(_04901_ ) );
AND3_X1 _12644_ ( .A1(_04890_ ), .A2(_04896_ ), .A3(_04901_ ), .ZN(_04902_ ) );
NAND3_X1 _12645_ ( .A1(_04403_ ), .A2(_04404_ ), .A3(_04880_ ), .ZN(_04903_ ) );
NAND2_X1 _12646_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [23] ), .ZN(_04904_ ) );
AND2_X1 _12647_ ( .A1(_04903_ ), .A2(_04904_ ), .ZN(_04905_ ) );
XNOR2_X1 _12648_ ( .A(_04905_ ), .B(_02307_ ), .ZN(_04906_ ) );
INV_X1 _12649_ ( .A(_04906_ ), .ZN(_04907_ ) );
BUF_X4 _12650_ ( .A(_04879_ ), .Z(_04908_ ) );
NAND2_X1 _12651_ ( .A1(_04428_ ), .A2(_04908_ ), .ZN(_04909_ ) );
NAND2_X1 _12652_ ( .A1(_02334_ ), .A2(fanout_net_5 ), .ZN(_04910_ ) );
NAND2_X1 _12653_ ( .A1(_04909_ ), .A2(_04910_ ), .ZN(_04911_ ) );
NAND3_X1 _12654_ ( .A1(_04907_ ), .A2(_02333_ ), .A3(_04911_ ), .ZN(_04912_ ) );
XNOR2_X1 _12655_ ( .A(_04911_ ), .B(_02333_ ), .ZN(_04913_ ) );
INV_X1 _12656_ ( .A(_04913_ ), .ZN(_04914_ ) );
NAND2_X1 _12657_ ( .A1(_04914_ ), .A2(_04907_ ), .ZN(_04915_ ) );
NAND3_X1 _12658_ ( .A1(_04450_ ), .A2(_04451_ ), .A3(_04881_ ), .ZN(_04916_ ) );
NAND2_X1 _12659_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [20] ), .ZN(_04917_ ) );
AND2_X2 _12660_ ( .A1(_04916_ ), .A2(_04917_ ), .ZN(_04918_ ) );
OAI21_X1 _12661_ ( .A(_04881_ ), .B1(_04473_ ), .B2(_04475_ ), .ZN(_04919_ ) );
NAND2_X1 _12662_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [21] ), .ZN(_04920_ ) );
AND2_X2 _12663_ ( .A1(_04919_ ), .A2(_04920_ ), .ZN(_04921_ ) );
INV_X1 _12664_ ( .A(_04477_ ), .ZN(_04922_ ) );
AND2_X1 _12665_ ( .A1(_04921_ ), .A2(_04922_ ), .ZN(_04923_ ) );
NOR2_X1 _12666_ ( .A1(_04921_ ), .A2(_04922_ ), .ZN(_04924_ ) );
OAI211_X1 _12667_ ( .A(_02382_ ), .B(_04918_ ), .C1(_04923_ ), .C2(_04924_ ), .ZN(_04925_ ) );
NAND3_X1 _12668_ ( .A1(_04919_ ), .A2(_04477_ ), .A3(_04920_ ), .ZN(_04926_ ) );
AOI21_X1 _12669_ ( .A(_04915_ ), .B1(_04925_ ), .B2(_04926_ ), .ZN(_04927_ ) );
NAND3_X1 _12670_ ( .A1(_04376_ ), .A2(_04377_ ), .A3(_04881_ ), .ZN(_04928_ ) );
NAND2_X1 _12671_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [16] ), .ZN(_04929_ ) );
AND2_X2 _12672_ ( .A1(_04928_ ), .A2(_04929_ ), .ZN(_04930_ ) );
NAND3_X1 _12673_ ( .A1(_04353_ ), .A2(_04354_ ), .A3(_04908_ ), .ZN(_04931_ ) );
NAND2_X1 _12674_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [17] ), .ZN(_04932_ ) );
AND2_X2 _12675_ ( .A1(_04931_ ), .A2(_04932_ ), .ZN(_04933_ ) );
INV_X1 _12676_ ( .A(_02458_ ), .ZN(_04934_ ) );
AND2_X1 _12677_ ( .A1(_04933_ ), .A2(_04934_ ), .ZN(_04935_ ) );
NOR2_X1 _12678_ ( .A1(_04933_ ), .A2(_04934_ ), .ZN(_04936_ ) );
OAI211_X1 _12679_ ( .A(_02480_ ), .B(_04930_ ), .C1(_04935_ ), .C2(_04936_ ), .ZN(_04937_ ) );
INV_X1 _12680_ ( .A(_04933_ ), .ZN(_04938_ ) );
OAI21_X1 _12681_ ( .A(_04937_ ), .B1(_04934_ ), .B2(_04938_ ), .ZN(_04939_ ) );
NAND3_X1 _12682_ ( .A1(_04326_ ), .A2(_04327_ ), .A3(_04908_ ), .ZN(_04940_ ) );
NAND2_X1 _12683_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [19] ), .ZN(_04941_ ) );
AND2_X2 _12684_ ( .A1(_04940_ ), .A2(_04941_ ), .ZN(_04942_ ) );
XNOR2_X1 _12685_ ( .A(_04942_ ), .B(_04330_ ), .ZN(_04943_ ) );
INV_X1 _12686_ ( .A(_04943_ ), .ZN(_04944_ ) );
NAND3_X1 _12687_ ( .A1(_04303_ ), .A2(_04304_ ), .A3(_04908_ ), .ZN(_04945_ ) );
NAND2_X1 _12688_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [18] ), .ZN(_04946_ ) );
AND2_X2 _12689_ ( .A1(_04945_ ), .A2(_04946_ ), .ZN(_04947_ ) );
XNOR2_X1 _12690_ ( .A(_04947_ ), .B(_02406_ ), .ZN(_04948_ ) );
INV_X1 _12691_ ( .A(_04948_ ), .ZN(_04949_ ) );
NAND3_X1 _12692_ ( .A1(_04939_ ), .A2(_04944_ ), .A3(_04949_ ), .ZN(_04950_ ) );
NAND3_X1 _12693_ ( .A1(_04944_ ), .A2(_02406_ ), .A3(_04947_ ), .ZN(_04951_ ) );
INV_X1 _12694_ ( .A(_04330_ ), .ZN(_04952_ ) );
INV_X1 _12695_ ( .A(_04942_ ), .ZN(_04953_ ) );
OAI211_X1 _12696_ ( .A(_04950_ ), .B(_04951_ ), .C1(_04952_ ), .C2(_04953_ ), .ZN(_04954_ ) );
XNOR2_X1 _12697_ ( .A(_04918_ ), .B(_02382_ ), .ZN(_04955_ ) );
XNOR2_X1 _12698_ ( .A(_04921_ ), .B(_04477_ ), .ZN(_04956_ ) );
NOR3_X1 _12699_ ( .A1(_04915_ ), .A2(_04955_ ), .A3(_04956_ ), .ZN(_04957_ ) );
AOI221_X4 _12700_ ( .A(_04927_ ), .B1(_02307_ ), .B2(_04905_ ), .C1(_04954_ ), .C2(_04957_ ), .ZN(_04958_ ) );
NAND3_X1 _12701_ ( .A1(_04619_ ), .A2(_04620_ ), .A3(_04879_ ), .ZN(_04959_ ) );
NAND2_X1 _12702_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [14] ), .ZN(_04960_ ) );
AND2_X2 _12703_ ( .A1(_04959_ ), .A2(_04960_ ), .ZN(_04961_ ) );
XNOR2_X2 _12704_ ( .A(_04961_ ), .B(_02525_ ), .ZN(_04962_ ) );
OR2_X1 _12705_ ( .A1(_04599_ ), .A2(fanout_net_5 ), .ZN(_04963_ ) );
NAND2_X1 _12706_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [15] ), .ZN(_04964_ ) );
AND2_X2 _12707_ ( .A1(_04963_ ), .A2(_04964_ ), .ZN(_04965_ ) );
INV_X2 _12708_ ( .A(_02503_ ), .ZN(_04966_ ) );
OR2_X1 _12709_ ( .A1(_04965_ ), .A2(_04966_ ), .ZN(_04967_ ) );
NAND3_X1 _12710_ ( .A1(_04963_ ), .A2(_04966_ ), .A3(_04964_ ), .ZN(_04968_ ) );
AOI21_X4 _12711_ ( .A(_04962_ ), .B1(_04967_ ), .B2(_04968_ ), .ZN(_04969_ ) );
NAND3_X1 _12712_ ( .A1(_04667_ ), .A2(_04648_ ), .A3(_04879_ ), .ZN(_04970_ ) );
NAND2_X1 _12713_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [13] ), .ZN(_04971_ ) );
AND2_X2 _12714_ ( .A1(_04970_ ), .A2(_04971_ ), .ZN(_04972_ ) );
XNOR2_X1 _12715_ ( .A(_04972_ ), .B(_02551_ ), .ZN(_04973_ ) );
INV_X1 _12716_ ( .A(_04973_ ), .ZN(_04974_ ) );
NAND3_X1 _12717_ ( .A1(_04643_ ), .A2(_04644_ ), .A3(_04880_ ), .ZN(_04975_ ) );
NAND2_X1 _12718_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [12] ), .ZN(_04976_ ) );
AND2_X2 _12719_ ( .A1(_04975_ ), .A2(_04976_ ), .ZN(_04977_ ) );
XNOR2_X1 _12720_ ( .A(_04977_ ), .B(_02574_ ), .ZN(_04978_ ) );
INV_X1 _12721_ ( .A(_04978_ ), .ZN(_04979_ ) );
AND3_X2 _12722_ ( .A1(_04969_ ), .A2(_04974_ ), .A3(_04979_ ), .ZN(_04980_ ) );
NAND3_X1 _12723_ ( .A1(_04523_ ), .A2(_04524_ ), .A3(_04908_ ), .ZN(_04981_ ) );
NAND2_X1 _12724_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [11] ), .ZN(_04982_ ) );
AND2_X1 _12725_ ( .A1(_04981_ ), .A2(_04982_ ), .ZN(_04983_ ) );
XNOR2_X2 _12726_ ( .A(_04983_ ), .B(_02670_ ), .ZN(_04984_ ) );
INV_X1 _12727_ ( .A(_04984_ ), .ZN(_04985_ ) );
NAND3_X1 _12728_ ( .A1(_04501_ ), .A2(_04502_ ), .A3(_04908_ ), .ZN(_04986_ ) );
NAND2_X1 _12729_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [10] ), .ZN(_04987_ ) );
AND2_X2 _12730_ ( .A1(_04986_ ), .A2(_04987_ ), .ZN(_04988_ ) );
XNOR2_X1 _12731_ ( .A(_04988_ ), .B(_02647_ ), .ZN(_04989_ ) );
INV_X1 _12732_ ( .A(_04989_ ), .ZN(_04990_ ) );
NAND3_X1 _12733_ ( .A1(_04980_ ), .A2(_04985_ ), .A3(_04990_ ), .ZN(_04991_ ) );
NAND3_X1 _12734_ ( .A1(_04569_ ), .A2(_04570_ ), .A3(_04908_ ), .ZN(_04992_ ) );
NAND2_X1 _12735_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [9] ), .ZN(_04993_ ) );
AND2_X2 _12736_ ( .A1(_04992_ ), .A2(_04993_ ), .ZN(_04994_ ) );
XNOR2_X1 _12737_ ( .A(_04994_ ), .B(_02624_ ), .ZN(_04995_ ) );
NAND3_X1 _12738_ ( .A1(_04547_ ), .A2(_04548_ ), .A3(_04908_ ), .ZN(_04996_ ) );
NAND2_X1 _12739_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [8] ), .ZN(_04997_ ) );
AND2_X2 _12740_ ( .A1(_04996_ ), .A2(_04997_ ), .ZN(_04998_ ) );
XNOR2_X1 _12741_ ( .A(_04998_ ), .B(_02600_ ), .ZN(_04999_ ) );
OR3_X4 _12742_ ( .A1(_04991_ ), .A2(_04995_ ), .A3(_04999_ ), .ZN(_05000_ ) );
NAND3_X1 _12743_ ( .A1(_04811_ ), .A2(_04812_ ), .A3(_04880_ ), .ZN(_05001_ ) );
NAND2_X1 _12744_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [7] ), .ZN(_05002_ ) );
AND2_X2 _12745_ ( .A1(_05001_ ), .A2(_05002_ ), .ZN(_05003_ ) );
XNOR2_X1 _12746_ ( .A(_05003_ ), .B(_02816_ ), .ZN(_05004_ ) );
INV_X1 _12747_ ( .A(_05004_ ), .ZN(_05005_ ) );
NAND3_X1 _12748_ ( .A1(_04834_ ), .A2(_04835_ ), .A3(_04880_ ), .ZN(_05006_ ) );
NAND2_X1 _12749_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [6] ), .ZN(_05007_ ) );
AND2_X2 _12750_ ( .A1(_05006_ ), .A2(_05007_ ), .ZN(_05008_ ) );
XNOR2_X1 _12751_ ( .A(_05008_ ), .B(_02792_ ), .ZN(_05009_ ) );
INV_X1 _12752_ ( .A(_05009_ ), .ZN(_05010_ ) );
NAND3_X1 _12753_ ( .A1(_04715_ ), .A2(_04716_ ), .A3(_04880_ ), .ZN(_05011_ ) );
NAND2_X1 _12754_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [4] ), .ZN(_05012_ ) );
AND2_X1 _12755_ ( .A1(_05011_ ), .A2(_05012_ ), .ZN(_05013_ ) );
INV_X1 _12756_ ( .A(_05013_ ), .ZN(_05014_ ) );
BUF_X4 _12757_ ( .A(_05014_ ), .Z(_05015_ ) );
NAND2_X1 _12758_ ( .A1(_04860_ ), .A2(_04908_ ), .ZN(_05016_ ) );
OR2_X1 _12759_ ( .A1(_04880_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05017_ ) );
NAND2_X2 _12760_ ( .A1(_05016_ ), .A2(_05017_ ), .ZN(_05018_ ) );
XNOR2_X1 _12761_ ( .A(_05018_ ), .B(_02875_ ), .ZN(_05019_ ) );
AOI211_X1 _12762_ ( .A(_05015_ ), .B(_05019_ ), .C1(_02862_ ), .C2(_02861_ ), .ZN(_05020_ ) );
AND3_X1 _12763_ ( .A1(_05016_ ), .A2(_02841_ ), .A3(_05017_ ), .ZN(_05021_ ) );
OAI211_X1 _12764_ ( .A(_05005_ ), .B(_05010_ ), .C1(_05020_ ), .C2(_05021_ ), .ZN(_05022_ ) );
NAND3_X1 _12765_ ( .A1(_02816_ ), .A2(_05002_ ), .A3(_05001_ ), .ZN(_05023_ ) );
NAND3_X1 _12766_ ( .A1(_05005_ ), .A2(_02792_ ), .A3(_05008_ ), .ZN(_05024_ ) );
AND3_X1 _12767_ ( .A1(_05022_ ), .A2(_05023_ ), .A3(_05024_ ), .ZN(_05025_ ) );
NAND3_X1 _12768_ ( .A1(_04738_ ), .A2(_04739_ ), .A3(_04908_ ), .ZN(_05026_ ) );
NAND2_X1 _12769_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [2] ), .ZN(_05027_ ) );
AND2_X2 _12770_ ( .A1(_05026_ ), .A2(_05027_ ), .ZN(_05028_ ) );
XNOR2_X1 _12771_ ( .A(_05028_ ), .B(_02695_ ), .ZN(_05029_ ) );
OAI21_X1 _12772_ ( .A(_04880_ ), .B1(_04693_ ), .B2(_04694_ ), .ZN(_05030_ ) );
NAND2_X1 _12773_ ( .A1(fanout_net_5 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_05031_ ) );
AND2_X1 _12774_ ( .A1(_05030_ ), .A2(_05031_ ), .ZN(_05032_ ) );
BUF_X4 _12775_ ( .A(_05032_ ), .Z(_05033_ ) );
XNOR2_X1 _12776_ ( .A(_05033_ ), .B(_02769_ ), .ZN(_05034_ ) );
NAND2_X1 _12777_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [1] ), .ZN(_05035_ ) );
NAND3_X1 _12778_ ( .A1(_04785_ ), .A2(_04786_ ), .A3(_04880_ ), .ZN(_05036_ ) );
NAND3_X1 _12779_ ( .A1(_02717_ ), .A2(_05035_ ), .A3(_05036_ ), .ZN(_05037_ ) );
INV_X1 _12780_ ( .A(_02717_ ), .ZN(_05038_ ) );
AND3_X1 _12781_ ( .A1(_05038_ ), .A2(_05035_ ), .A3(_05036_ ), .ZN(_05039_ ) );
AND2_X2 _12782_ ( .A1(_05036_ ), .A2(_05035_ ), .ZN(_05040_ ) );
NOR2_X1 _12783_ ( .A1(_05040_ ), .A2(_05038_ ), .ZN(_05041_ ) );
NAND2_X1 _12784_ ( .A1(_04764_ ), .A2(_04880_ ), .ZN(_05042_ ) );
NAND2_X1 _12785_ ( .A1(_02720_ ), .A2(\ID_EX_typ [4] ), .ZN(_05043_ ) );
NAND2_X2 _12786_ ( .A1(_05042_ ), .A2(_05043_ ), .ZN(_05044_ ) );
OAI22_X1 _12787_ ( .A1(_05039_ ), .A2(_05041_ ), .B1(_04743_ ), .B2(_05044_ ), .ZN(_05045_ ) );
AOI211_X1 _12788_ ( .A(_05029_ ), .B(_05034_ ), .C1(_05037_ ), .C2(_05045_ ), .ZN(_05046_ ) );
INV_X1 _12789_ ( .A(_02695_ ), .ZN(_05047_ ) );
INV_X1 _12790_ ( .A(_05028_ ), .ZN(_05048_ ) );
NOR3_X1 _12791_ ( .A1(_05034_ ), .A2(_05047_ ), .A3(_05048_ ), .ZN(_05049_ ) );
AOI21_X1 _12792_ ( .A(_02769_ ), .B1(_05030_ ), .B2(_05031_ ), .ZN(_05050_ ) );
OR3_X1 _12793_ ( .A1(_05046_ ), .A2(_05049_ ), .A3(_05050_ ), .ZN(_05051_ ) );
XNOR2_X1 _12794_ ( .A(_05013_ ), .B(_02864_ ), .ZN(_05052_ ) );
NOR4_X1 _12795_ ( .A1(_05019_ ), .A2(_05004_ ), .A3(_05009_ ), .A4(_05052_ ), .ZN(_05053_ ) );
NAND2_X1 _12796_ ( .A1(_05051_ ), .A2(_05053_ ), .ZN(_05054_ ) );
AOI21_X2 _12797_ ( .A(_05000_ ), .B1(_05025_ ), .B2(_05054_ ), .ZN(_05055_ ) );
XNOR2_X1 _12798_ ( .A(_04965_ ), .B(_02503_ ), .ZN(_05056_ ) );
INV_X1 _12799_ ( .A(_02526_ ), .ZN(_05057_ ) );
INV_X1 _12800_ ( .A(_04961_ ), .ZN(_05058_ ) );
NOR3_X1 _12801_ ( .A1(_05056_ ), .A2(_05057_ ), .A3(_05058_ ), .ZN(_05059_ ) );
NAND2_X1 _12802_ ( .A1(_04990_ ), .A2(_04985_ ), .ZN(_05060_ ) );
NAND3_X1 _12803_ ( .A1(_02624_ ), .A2(_04992_ ), .A3(_04993_ ), .ZN(_05061_ ) );
INV_X1 _12804_ ( .A(_02624_ ), .ZN(_05062_ ) );
AND2_X1 _12805_ ( .A1(_04994_ ), .A2(_05062_ ), .ZN(_05063_ ) );
NOR2_X1 _12806_ ( .A1(_04994_ ), .A2(_05062_ ), .ZN(_05064_ ) );
OAI211_X1 _12807_ ( .A(_02600_ ), .B(_04998_ ), .C1(_05063_ ), .C2(_05064_ ), .ZN(_05065_ ) );
AOI21_X1 _12808_ ( .A(_05060_ ), .B1(_05061_ ), .B2(_05065_ ), .ZN(_05066_ ) );
NAND3_X1 _12809_ ( .A1(_04985_ ), .A2(_02647_ ), .A3(_04988_ ), .ZN(_05067_ ) );
INV_X1 _12810_ ( .A(_02670_ ), .ZN(_05068_ ) );
INV_X1 _12811_ ( .A(_04983_ ), .ZN(_05069_ ) );
OAI21_X1 _12812_ ( .A(_05067_ ), .B1(_05068_ ), .B2(_05069_ ), .ZN(_05070_ ) );
OAI21_X1 _12813_ ( .A(_04980_ ), .B1(_05066_ ), .B2(_05070_ ), .ZN(_05071_ ) );
INV_X1 _12814_ ( .A(_02574_ ), .ZN(_05072_ ) );
INV_X1 _12815_ ( .A(_04977_ ), .ZN(_05073_ ) );
NOR3_X1 _12816_ ( .A1(_04973_ ), .A2(_05072_ ), .A3(_05073_ ), .ZN(_05074_ ) );
AND3_X1 _12817_ ( .A1(_02552_ ), .A2(_04971_ ), .A3(_04970_ ), .ZN(_05075_ ) );
OAI21_X1 _12818_ ( .A(_04969_ ), .B1(_05074_ ), .B2(_05075_ ), .ZN(_05076_ ) );
INV_X1 _12819_ ( .A(_04965_ ), .ZN(_05077_ ) );
OAI211_X1 _12820_ ( .A(_05071_ ), .B(_05076_ ), .C1(_04966_ ), .C2(_05077_ ), .ZN(_05078_ ) );
NOR3_X1 _12821_ ( .A1(_05055_ ), .A2(_05059_ ), .A3(_05078_ ), .ZN(_05079_ ) );
XNOR2_X1 _12822_ ( .A(_04933_ ), .B(_02458_ ), .ZN(_05080_ ) );
XNOR2_X1 _12823_ ( .A(_04930_ ), .B(_02480_ ), .ZN(_05081_ ) );
NOR4_X1 _12824_ ( .A1(_04943_ ), .A2(_04948_ ), .A3(_05080_ ), .A4(_05081_ ), .ZN(_05082_ ) );
NAND2_X1 _12825_ ( .A1(_04957_ ), .A2(_05082_ ), .ZN(_05083_ ) );
OAI211_X2 _12826_ ( .A(_04912_ ), .B(_04958_ ), .C1(_05079_ ), .C2(_05083_ ), .ZN(_05084_ ) );
NAND3_X1 _12827_ ( .A1(_04196_ ), .A2(_04198_ ), .A3(_04881_ ), .ZN(_05085_ ) );
NAND2_X1 _12828_ ( .A1(_02249_ ), .A2(\ID_EX_typ [4] ), .ZN(_05086_ ) );
NAND2_X1 _12829_ ( .A1(_05085_ ), .A2(_05086_ ), .ZN(_05087_ ) );
XNOR2_X1 _12830_ ( .A(_02248_ ), .B(_05087_ ), .ZN(_05088_ ) );
NAND3_X1 _12831_ ( .A1(_04221_ ), .A2(_04223_ ), .A3(_04881_ ), .ZN(_05089_ ) );
NAND2_X1 _12832_ ( .A1(_02966_ ), .A2(\ID_EX_typ [4] ), .ZN(_05090_ ) );
NAND2_X1 _12833_ ( .A1(_05089_ ), .A2(_05090_ ), .ZN(_05091_ ) );
XNOR2_X1 _12834_ ( .A(_05091_ ), .B(_02964_ ), .ZN(_05092_ ) );
NOR2_X1 _12835_ ( .A1(_05088_ ), .A2(_05092_ ), .ZN(_05093_ ) );
NAND3_X1 _12836_ ( .A1(_04269_ ), .A2(_04250_ ), .A3(_04881_ ), .ZN(_05094_ ) );
NAND2_X1 _12837_ ( .A1(_02272_ ), .A2(\ID_EX_typ [4] ), .ZN(_05095_ ) );
NAND2_X1 _12838_ ( .A1(_05094_ ), .A2(_05095_ ), .ZN(_05096_ ) );
XNOR2_X1 _12839_ ( .A(_05096_ ), .B(_02271_ ), .ZN(_05097_ ) );
INV_X1 _12840_ ( .A(_05097_ ), .ZN(_05098_ ) );
NAND3_X1 _12841_ ( .A1(_04245_ ), .A2(_04247_ ), .A3(_04881_ ), .ZN(_05099_ ) );
NAND2_X1 _12842_ ( .A1(_02968_ ), .A2(\ID_EX_typ [4] ), .ZN(_05100_ ) );
NAND2_X1 _12843_ ( .A1(_05099_ ), .A2(_05100_ ), .ZN(_05101_ ) );
XNOR2_X1 _12844_ ( .A(_05101_ ), .B(_02940_ ), .ZN(_05102_ ) );
INV_X1 _12845_ ( .A(_05102_ ), .ZN(_05103_ ) );
AND4_X2 _12846_ ( .A1(_05084_ ), .A2(_05093_ ), .A3(_05098_ ), .A4(_05103_ ), .ZN(_05104_ ) );
AND3_X1 _12847_ ( .A1(_05103_ ), .A2(_02271_ ), .A3(_05096_ ), .ZN(_05105_ ) );
AOI22_X1 _12848_ ( .A1(_05099_ ), .A2(_05100_ ), .B1(_02939_ ), .B2(_02938_ ), .ZN(_05106_ ) );
OAI21_X1 _12849_ ( .A(_05093_ ), .B1(_05105_ ), .B2(_05106_ ), .ZN(_05107_ ) );
INV_X1 _12850_ ( .A(_05088_ ), .ZN(_05108_ ) );
NAND3_X1 _12851_ ( .A1(_05108_ ), .A2(_02965_ ), .A3(_05091_ ), .ZN(_05109_ ) );
NAND2_X1 _12852_ ( .A1(_02248_ ), .A2(_05087_ ), .ZN(_05110_ ) );
NAND3_X1 _12853_ ( .A1(_05107_ ), .A2(_05109_ ), .A3(_05110_ ), .ZN(_05111_ ) );
OAI21_X2 _12854_ ( .A(_04902_ ), .B1(_05104_ ), .B2(_05111_ ), .ZN(_05112_ ) );
NOR2_X1 _12855_ ( .A1(_04885_ ), .A2(_03005_ ), .ZN(_05113_ ) );
NOR2_X1 _12856_ ( .A1(_04876_ ), .A2(_02172_ ), .ZN(_05114_ ) );
AND2_X1 _12857_ ( .A1(_05114_ ), .A2(_04888_ ), .ZN(_05115_ ) );
INV_X1 _12858_ ( .A(_04899_ ), .ZN(_05116_ ) );
NAND3_X1 _12859_ ( .A1(_05116_ ), .A2(_04896_ ), .A3(_02226_ ), .ZN(_05117_ ) );
OAI21_X1 _12860_ ( .A(_05117_ ), .B1(_04894_ ), .B2(_04893_ ), .ZN(_05118_ ) );
AOI211_X1 _12861_ ( .A(_05113_ ), .B(_05115_ ), .C1(_04890_ ), .C2(_05118_ ), .ZN(_05119_ ) );
AND2_X2 _12862_ ( .A1(_05112_ ), .A2(_05119_ ), .ZN(_05120_ ) );
MUX2_X1 _12863_ ( .A(_04871_ ), .B(_04873_ ), .S(_05120_ ), .Z(_05121_ ) );
AND2_X1 _12864_ ( .A1(_02717_ ), .A2(_04787_ ), .ZN(_05122_ ) );
OAI21_X1 _12865_ ( .A(_04742_ ), .B1(_04791_ ), .B2(_05122_ ), .ZN(_05123_ ) );
AND2_X1 _12866_ ( .A1(_02695_ ), .A2(_04740_ ), .ZN(_05124_ ) );
INV_X1 _12867_ ( .A(_05124_ ), .ZN(_05125_ ) );
OAI211_X1 _12868_ ( .A(_05123_ ), .B(_05125_ ), .C1(_02769_ ), .C2(_04695_ ), .ZN(_05126_ ) );
NAND3_X1 _12869_ ( .A1(_04695_ ), .A2(_02765_ ), .A3(_02764_ ), .ZN(_05127_ ) );
AND2_X1 _12870_ ( .A1(_05126_ ), .A2(_05127_ ), .ZN(_05128_ ) );
AND3_X1 _12871_ ( .A1(_05128_ ), .A2(_04861_ ), .A3(_04719_ ), .ZN(_05129_ ) );
NAND2_X1 _12872_ ( .A1(_05129_ ), .A2(_04839_ ), .ZN(_05130_ ) );
AND3_X1 _12873_ ( .A1(_04815_ ), .A2(_02792_ ), .A3(_04836_ ), .ZN(_05131_ ) );
NAND3_X1 _12874_ ( .A1(_04861_ ), .A2(_02864_ ), .A3(_04717_ ), .ZN(_05132_ ) );
OAI21_X1 _12875_ ( .A(_05132_ ), .B1(_02875_ ), .B2(_04860_ ), .ZN(_05133_ ) );
AOI221_X1 _12876_ ( .A(_05131_ ), .B1(_02816_ ), .B2(_04813_ ), .C1(_05133_ ), .C2(_04839_ ), .ZN(_05134_ ) );
NAND2_X1 _12877_ ( .A1(_05130_ ), .A2(_05134_ ), .ZN(_05135_ ) );
NAND2_X1 _12878_ ( .A1(_05135_ ), .A2(_04673_ ), .ZN(_05136_ ) );
NAND3_X1 _12879_ ( .A1(_04600_ ), .A2(_02526_ ), .A3(_04621_ ), .ZN(_05137_ ) );
INV_X1 _12880_ ( .A(_04599_ ), .ZN(_05138_ ) );
NAND3_X1 _12881_ ( .A1(_04527_ ), .A2(_02647_ ), .A3(_04503_ ), .ZN(_05139_ ) );
OAI21_X1 _12882_ ( .A(_05139_ ), .B1(_05068_ ), .B2(_04526_ ), .ZN(_05140_ ) );
AND3_X1 _12883_ ( .A1(_04574_ ), .A2(_02600_ ), .A3(_04549_ ), .ZN(_05141_ ) );
OR2_X1 _12884_ ( .A1(_05141_ ), .A2(_04572_ ), .ZN(_05142_ ) );
AOI21_X2 _12885_ ( .A(_05140_ ), .B1(_05142_ ), .B2(_04528_ ), .ZN(_05143_ ) );
OAI221_X1 _12886_ ( .A(_05137_ ), .B1(_04966_ ), .B2(_05138_ ), .C1(_05143_ ), .C2(_04672_ ), .ZN(_05144_ ) );
NAND2_X1 _12887_ ( .A1(_02574_ ), .A2(_04645_ ), .ZN(_05145_ ) );
NOR3_X1 _12888_ ( .A1(_04669_ ), .A2(_04670_ ), .A3(_05145_ ), .ZN(_05146_ ) );
OR2_X1 _12889_ ( .A1(_05146_ ), .A2(_04669_ ), .ZN(_05147_ ) );
AOI21_X1 _12890_ ( .A(_05144_ ), .B1(_04624_ ), .B2(_05147_ ), .ZN(_05148_ ) );
AND2_X1 _12891_ ( .A1(_05136_ ), .A2(_05148_ ), .ZN(_05149_ ) );
INV_X1 _12892_ ( .A(_05149_ ), .ZN(_05150_ ) );
NAND2_X1 _12893_ ( .A1(_05150_ ), .A2(_04482_ ), .ZN(_05151_ ) );
AND2_X1 _12894_ ( .A1(_02406_ ), .A2(_04305_ ), .ZN(_05152_ ) );
NAND2_X1 _12895_ ( .A1(_04331_ ), .A2(_05152_ ), .ZN(_05153_ ) );
OAI21_X1 _12896_ ( .A(_05153_ ), .B1(_04952_ ), .B2(_04329_ ), .ZN(_05154_ ) );
AND2_X1 _12897_ ( .A1(_02480_ ), .A2(_04378_ ), .ZN(_05155_ ) );
AND2_X1 _12898_ ( .A1(_04357_ ), .A2(_05155_ ), .ZN(_05156_ ) );
AOI21_X1 _12899_ ( .A(_05156_ ), .B1(_02458_ ), .B2(_04355_ ), .ZN(_05157_ ) );
INV_X1 _12900_ ( .A(_05157_ ), .ZN(_05158_ ) );
AOI21_X1 _12901_ ( .A(_05154_ ), .B1(_05158_ ), .B2(_04332_ ), .ZN(_05159_ ) );
INV_X1 _12902_ ( .A(_04481_ ), .ZN(_05160_ ) );
NOR2_X1 _12903_ ( .A1(_05159_ ), .A2(_05160_ ), .ZN(_05161_ ) );
AND2_X1 _12904_ ( .A1(_02333_ ), .A2(_04428_ ), .ZN(_05162_ ) );
NAND2_X1 _12905_ ( .A1(_04407_ ), .A2(_05162_ ), .ZN(_05163_ ) );
OAI21_X1 _12906_ ( .A(_05163_ ), .B1(_02900_ ), .B2(_04406_ ), .ZN(_05164_ ) );
INV_X1 _12907_ ( .A(_04431_ ), .ZN(_05165_ ) );
INV_X1 _12908_ ( .A(_04478_ ), .ZN(_05166_ ) );
AND2_X1 _12909_ ( .A1(_02382_ ), .A2(_04452_ ), .ZN(_05167_ ) );
NAND2_X1 _12910_ ( .A1(_04480_ ), .A2(_05167_ ), .ZN(_05168_ ) );
AOI21_X1 _12911_ ( .A(_05165_ ), .B1(_05166_ ), .B2(_05168_ ), .ZN(_05169_ ) );
NOR3_X1 _12912_ ( .A1(_05161_ ), .A2(_05164_ ), .A3(_05169_ ), .ZN(_05170_ ) );
NAND2_X2 _12913_ ( .A1(_05151_ ), .A2(_05170_ ), .ZN(_05171_ ) );
NAND2_X1 _12914_ ( .A1(_05171_ ), .A2(_04273_ ), .ZN(_05172_ ) );
INV_X1 _12915_ ( .A(_02271_ ), .ZN(_05173_ ) );
NOR2_X1 _12916_ ( .A1(_05173_ ), .A2(_04270_ ), .ZN(_05174_ ) );
AND2_X1 _12917_ ( .A1(_04249_ ), .A2(_05174_ ), .ZN(_05175_ ) );
INV_X1 _12918_ ( .A(_04248_ ), .ZN(_05176_ ) );
AND2_X1 _12919_ ( .A1(_05176_ ), .A2(_02940_ ), .ZN(_05177_ ) );
OAI211_X1 _12920_ ( .A(_04203_ ), .B(_04225_ ), .C1(_05175_ ), .C2(_05177_ ), .ZN(_05178_ ) );
INV_X1 _12921_ ( .A(_04224_ ), .ZN(_05179_ ) );
NAND4_X1 _12922_ ( .A1(_04201_ ), .A2(_02965_ ), .A3(_04202_ ), .A4(_05179_ ), .ZN(_05180_ ) );
AND3_X1 _12923_ ( .A1(_05178_ ), .A2(_04201_ ), .A3(_05180_ ), .ZN(_05181_ ) );
NOR2_X1 _12924_ ( .A1(_04177_ ), .A2(_05181_ ), .ZN(_05182_ ) );
INV_X1 _12925_ ( .A(_04129_ ), .ZN(_05183_ ) );
INV_X1 _12926_ ( .A(_04151_ ), .ZN(_05184_ ) );
AOI21_X1 _12927_ ( .A(_04175_ ), .B1(_05184_ ), .B2(_02226_ ), .ZN(_05185_ ) );
NOR3_X1 _12928_ ( .A1(_05183_ ), .A2(_04174_ ), .A3(_05185_ ), .ZN(_05186_ ) );
INV_X1 _12929_ ( .A(_02172_ ), .ZN(_05187_ ) );
NAND3_X1 _12930_ ( .A1(_05187_ ), .A2(_04128_ ), .A3(_04102_ ), .ZN(_05188_ ) );
OAI21_X1 _12931_ ( .A(_05188_ ), .B1(_04878_ ), .B2(_04127_ ), .ZN(_05189_ ) );
NOR3_X1 _12932_ ( .A1(_05182_ ), .A2(_05186_ ), .A3(_05189_ ), .ZN(_05190_ ) );
AND2_X1 _12933_ ( .A1(_04865_ ), .A2(\ID_EX_typ [2] ), .ZN(_05191_ ) );
AND3_X1 _12934_ ( .A1(_05172_ ), .A2(_05190_ ), .A3(_05191_ ), .ZN(_05192_ ) );
AND2_X1 _12935_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_4 ), .ZN(_05193_ ) );
AND2_X2 _12936_ ( .A1(_05193_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05194_ ) );
INV_X1 _12937_ ( .A(_05194_ ), .ZN(_05195_ ) );
AOI21_X1 _12938_ ( .A(_05195_ ), .B1(_05172_ ), .B2(_05190_ ), .ZN(_05196_ ) );
NOR3_X1 _12939_ ( .A1(_05192_ ), .A2(_05196_ ), .A3(_04866_ ), .ZN(_05197_ ) );
AOI221_X4 _12940_ ( .A(_04046_ ), .B1(_04864_ ), .B2(_04866_ ), .C1(_05121_ ), .C2(_05197_ ), .ZN(_05198_ ) );
NOR3_X1 _12941_ ( .A1(_04862_ ), .A2(_04672_ ), .A3(_04576_ ), .ZN(_05199_ ) );
NAND3_X1 _12942_ ( .A1(_04273_ ), .A2(_04482_ ), .A3(_05199_ ), .ZN(_05200_ ) );
AND2_X2 _12943_ ( .A1(_05200_ ), .A2(_04046_ ), .ZN(_05201_ ) );
NOR2_X4 _12944_ ( .A1(_05198_ ), .A2(_05201_ ), .ZN(_05202_ ) );
BUF_X8 _12945_ ( .A(_05202_ ), .Z(_05203_ ) );
MUX2_X1 _12946_ ( .A(_03926_ ), .B(_04044_ ), .S(_05203_ ), .Z(_05204_ ) );
OR2_X2 _12947_ ( .A1(_05204_ ), .A2(\ID_EX_typ [3] ), .ZN(_05205_ ) );
INV_X2 _12948_ ( .A(_03885_ ), .ZN(_05206_ ) );
BUF_X4 _12949_ ( .A(_05206_ ), .Z(_05207_ ) );
BUF_X4 _12950_ ( .A(_05207_ ), .Z(_05208_ ) );
INV_X1 _12951_ ( .A(\ID_EX_typ [3] ), .ZN(_05209_ ) );
BUF_X2 _12952_ ( .A(_05209_ ), .Z(_05210_ ) );
BUF_X4 _12953_ ( .A(_05210_ ), .Z(_05211_ ) );
XNOR2_X1 _12954_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_05212_ ) );
XNOR2_X1 _12955_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_05213_ ) );
AND2_X1 _12956_ ( .A1(_05212_ ), .A2(_05213_ ), .ZN(_05214_ ) );
XNOR2_X1 _12957_ ( .A(fanout_net_3 ), .B(\ID_EX_csr [0] ), .ZN(_05215_ ) );
XNOR2_X1 _12958_ ( .A(\EX_LS_dest_csreg_mem [1] ), .B(\ID_EX_csr [1] ), .ZN(_05216_ ) );
AND2_X1 _12959_ ( .A1(_05215_ ), .A2(_05216_ ), .ZN(_05217_ ) );
XNOR2_X1 _12960_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_05218_ ) );
XNOR2_X1 _12961_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_05219_ ) );
AND2_X1 _12962_ ( .A1(_05218_ ), .A2(_05219_ ), .ZN(_05220_ ) );
XNOR2_X1 _12963_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_05221_ ) );
XNOR2_X1 _12964_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_05222_ ) );
AND2_X1 _12965_ ( .A1(_05221_ ), .A2(_05222_ ), .ZN(_05223_ ) );
AND4_X2 _12966_ ( .A1(_05214_ ), .A2(_05217_ ), .A3(_05220_ ), .A4(_05223_ ), .ZN(_05224_ ) );
XNOR2_X1 _12967_ ( .A(\EX_LS_dest_csreg_mem [8] ), .B(\ID_EX_csr [8] ), .ZN(_05225_ ) );
XNOR2_X1 _12968_ ( .A(\EX_LS_dest_csreg_mem [9] ), .B(\ID_EX_csr [9] ), .ZN(_05226_ ) );
XNOR2_X1 _12969_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .ZN(_05227_ ) );
XNOR2_X1 _12970_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_05228_ ) );
AND4_X2 _12971_ ( .A1(_05225_ ), .A2(_05226_ ), .A3(_05227_ ), .A4(_05228_ ), .ZN(_05229_ ) );
NAND2_X1 _12972_ ( .A1(_05224_ ), .A2(_05229_ ), .ZN(_05230_ ) );
BUF_X4 _12973_ ( .A(_05230_ ), .Z(_05231_ ) );
INV_X2 _12974_ ( .A(_02128_ ), .ZN(_05232_ ) );
NOR2_X1 _12975_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_05233_ ) );
INV_X1 _12976_ ( .A(\ID_EX_csr [7] ), .ZN(_05234_ ) );
AND3_X2 _12977_ ( .A1(_05233_ ), .A2(_05234_ ), .A3(\ID_EX_csr [6] ), .ZN(_05235_ ) );
AND2_X1 _12978_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_05236_ ) );
NOR2_X1 _12979_ ( .A1(\ID_EX_csr [10] ), .A2(\ID_EX_csr [11] ), .ZN(_05237_ ) );
AND2_X1 _12980_ ( .A1(_05236_ ), .A2(_05237_ ), .ZN(_05238_ ) );
AND2_X1 _12981_ ( .A1(_05235_ ), .A2(_05238_ ), .ZN(_05239_ ) );
BUF_X4 _12982_ ( .A(_05239_ ), .Z(_05240_ ) );
BUF_X4 _12983_ ( .A(_05240_ ), .Z(_05241_ ) );
INV_X1 _12984_ ( .A(\ID_EX_csr [3] ), .ZN(_05242_ ) );
INV_X1 _12985_ ( .A(\ID_EX_csr [2] ), .ZN(_05243_ ) );
NAND3_X1 _12986_ ( .A1(_05242_ ), .A2(_05243_ ), .A3(\ID_EX_csr [1] ), .ZN(_05244_ ) );
NOR2_X1 _12987_ ( .A1(_05244_ ), .A2(\ID_EX_csr [0] ), .ZN(_05245_ ) );
BUF_X2 _12988_ ( .A(_05245_ ), .Z(_05246_ ) );
NAND3_X1 _12989_ ( .A1(_05241_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_05246_ ), .ZN(_05247_ ) );
INV_X1 _12990_ ( .A(\ID_EX_csr [1] ), .ZN(_05248_ ) );
NAND3_X1 _12991_ ( .A1(_05248_ ), .A2(_05242_ ), .A3(\ID_EX_csr [0] ), .ZN(_05249_ ) );
NOR2_X1 _12992_ ( .A1(_05249_ ), .A2(\ID_EX_csr [2] ), .ZN(_05250_ ) );
NOR2_X1 _12993_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_05251_ ) );
INV_X1 _12994_ ( .A(\ID_EX_csr [5] ), .ZN(_05252_ ) );
AND3_X1 _12995_ ( .A1(_05251_ ), .A2(_05252_ ), .A3(\ID_EX_csr [4] ), .ZN(_05253_ ) );
AND2_X1 _12996_ ( .A1(_05250_ ), .A2(_05253_ ), .ZN(_05254_ ) );
AND3_X1 _12997_ ( .A1(_05236_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_05255_ ) );
NAND2_X1 _12998_ ( .A1(_05254_ ), .A2(_05255_ ), .ZN(_05256_ ) );
BUF_X4 _12999_ ( .A(_05250_ ), .Z(_05257_ ) );
BUF_X4 _13000_ ( .A(_05257_ ), .Z(_05258_ ) );
BUF_X4 _13001_ ( .A(_05235_ ), .Z(_05259_ ) );
BUF_X4 _13002_ ( .A(_05238_ ), .Z(_05260_ ) );
BUF_X2 _13003_ ( .A(_05260_ ), .Z(_05261_ ) );
NAND4_X1 _13004_ ( .A1(_05258_ ), .A2(_05259_ ), .A3(_05261_ ), .A4(\mepc [30] ), .ZN(_05262_ ) );
NOR2_X1 _13005_ ( .A1(_05249_ ), .A2(_05243_ ), .ZN(_05263_ ) );
BUF_X2 _13006_ ( .A(_05263_ ), .Z(_05264_ ) );
BUF_X2 _13007_ ( .A(_05260_ ), .Z(_05265_ ) );
AND2_X1 _13008_ ( .A1(_05251_ ), .A2(_05233_ ), .ZN(_05266_ ) );
BUF_X4 _13009_ ( .A(_05266_ ), .Z(_05267_ ) );
BUF_X2 _13010_ ( .A(_05267_ ), .Z(_05268_ ) );
NAND4_X1 _13011_ ( .A1(_05264_ ), .A2(_05265_ ), .A3(_05268_ ), .A4(\mtvec [30] ), .ZN(_05269_ ) );
NAND4_X1 _13012_ ( .A1(_05247_ ), .A2(_05256_ ), .A3(_05262_ ), .A4(_05269_ ), .ZN(_05270_ ) );
NOR2_X1 _13013_ ( .A1(\ID_EX_csr [1] ), .A2(\ID_EX_csr [0] ), .ZN(_05271_ ) );
AND3_X1 _13014_ ( .A1(_05271_ ), .A2(_05242_ ), .A3(_05243_ ), .ZN(_05272_ ) );
AND2_X2 _13015_ ( .A1(_05272_ ), .A2(_05267_ ), .ZN(_05273_ ) );
AND3_X1 _13016_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_05265_ ), .ZN(_05274_ ) );
OAI22_X1 _13017_ ( .A1(_05231_ ), .A2(_05232_ ), .B1(_05270_ ), .B2(_05274_ ), .ZN(_05275_ ) );
NAND4_X1 _13018_ ( .A1(_05224_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_02128_ ), .A4(_05229_ ), .ZN(_05276_ ) );
NAND2_X1 _13019_ ( .A1(_05275_ ), .A2(_05276_ ), .ZN(_05277_ ) );
OAI211_X1 _13020_ ( .A(_05205_ ), .B(_05208_ ), .C1(_05211_ ), .C2(_05277_ ), .ZN(_05278_ ) );
BUF_X2 _13021_ ( .A(_03885_ ), .Z(_05279_ ) );
BUF_X4 _13022_ ( .A(_05279_ ), .Z(_05280_ ) );
OAI21_X1 _13023_ ( .A(fanout_net_4 ), .B1(_03010_ ), .B2(_02980_ ), .ZN(_05281_ ) );
OAI211_X1 _13024_ ( .A(_05280_ ), .B(_05281_ ), .C1(_04044_ ), .C2(fanout_net_4 ), .ZN(_05282_ ) );
AOI21_X1 _13025_ ( .A(_03907_ ), .B1(_05278_ ), .B2(_05282_ ), .ZN(_00122_ ) );
BUF_X4 _13026_ ( .A(_05209_ ), .Z(_05283_ ) );
AND4_X1 _13027_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_05284_ ) );
AND4_X1 _13028_ ( .A1(\ID_EX_pc [13] ), .A2(_05284_ ), .A3(\ID_EX_pc [12] ), .A4(_03915_ ), .ZN(_05285_ ) );
AND2_X1 _13029_ ( .A1(_03914_ ), .A2(_05285_ ), .ZN(_05286_ ) );
AND4_X1 _13030_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_05287_ ) );
AND2_X1 _13031_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_05288_ ) );
AND4_X1 _13032_ ( .A1(\ID_EX_pc [21] ), .A2(_05287_ ), .A3(\ID_EX_pc [20] ), .A4(_05288_ ), .ZN(_05289_ ) );
NAND2_X1 _13033_ ( .A1(_05286_ ), .A2(_05289_ ), .ZN(_05290_ ) );
INV_X1 _13034_ ( .A(\ID_EX_pc [27] ), .ZN(_05291_ ) );
INV_X1 _13035_ ( .A(\ID_EX_pc [26] ), .ZN(_05292_ ) );
NOR3_X1 _13036_ ( .A1(_05290_ ), .A2(_05291_ ), .A3(_05292_ ), .ZN(_05293_ ) );
NAND2_X1 _13037_ ( .A1(_05293_ ), .A2(\ID_EX_pc [28] ), .ZN(_05294_ ) );
XNOR2_X1 _13038_ ( .A(_05294_ ), .B(\ID_EX_pc [29] ), .ZN(_05295_ ) );
OAI21_X1 _13039_ ( .A(_05295_ ), .B1(_05198_ ), .B2(_05201_ ), .ZN(_05296_ ) );
INV_X1 _13040_ ( .A(_05202_ ), .ZN(_05297_ ) );
NAND2_X1 _13041_ ( .A1(_04037_ ), .A2(_04038_ ), .ZN(_05298_ ) );
XOR2_X1 _13042_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .Z(_05299_ ) );
XNOR2_X1 _13043_ ( .A(_05298_ ), .B(_05299_ ), .ZN(_05300_ ) );
OAI211_X1 _13044_ ( .A(_05283_ ), .B(_05296_ ), .C1(_05297_ ), .C2(_05300_ ), .ZN(_05301_ ) );
INV_X1 _13045_ ( .A(\ID_EX_csr [6] ), .ZN(_05302_ ) );
OAI221_X1 _13046_ ( .A(_05225_ ), .B1(\EX_LS_dest_csreg_mem [3] ), .B2(_05242_ ), .C1(\EX_LS_dest_csreg_mem [6] ), .C2(_05302_ ), .ZN(_05303_ ) );
INV_X1 _13047_ ( .A(\EX_LS_dest_csreg_mem [3] ), .ZN(_05304_ ) );
OAI221_X1 _13048_ ( .A(_05212_ ), .B1(_05304_ ), .B2(\ID_EX_csr [3] ), .C1(_03876_ ), .C2(\ID_EX_csr [6] ), .ZN(_05305_ ) );
INV_X2 _13049_ ( .A(\EX_LS_dest_csreg_mem [1] ), .ZN(_05306_ ) );
INV_X1 _13050_ ( .A(\EX_LS_dest_csreg_mem [5] ), .ZN(_05307_ ) );
OAI22_X1 _13051_ ( .A1(_05306_ ), .A2(\ID_EX_csr [1] ), .B1(_05307_ ), .B2(\ID_EX_csr [5] ), .ZN(_05308_ ) );
OAI22_X1 _13052_ ( .A1(\EX_LS_dest_csreg_mem [1] ), .A2(_05248_ ), .B1(_05252_ ), .B2(\EX_LS_dest_csreg_mem [5] ), .ZN(_05309_ ) );
NOR4_X1 _13053_ ( .A1(_05303_ ), .A2(_05305_ ), .A3(_05308_ ), .A4(_05309_ ), .ZN(_05310_ ) );
AND4_X1 _13054_ ( .A1(_05227_ ), .A2(_05218_ ), .A3(_05228_ ), .A4(_05215_ ), .ZN(_05311_ ) );
AND4_X1 _13055_ ( .A1(_02128_ ), .A2(_05311_ ), .A3(_05226_ ), .A4(_05221_ ), .ZN(_05312_ ) );
AND2_X1 _13056_ ( .A1(_05310_ ), .A2(_05312_ ), .ZN(_05313_ ) );
INV_X1 _13057_ ( .A(_05313_ ), .ZN(_05314_ ) );
BUF_X4 _13058_ ( .A(_05314_ ), .Z(_05315_ ) );
AND4_X1 _13059_ ( .A1(\ID_EX_csr [10] ), .A2(_05252_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_05316_ ) );
AND3_X1 _13060_ ( .A1(_05316_ ), .A2(_05236_ ), .A3(_05251_ ), .ZN(_05317_ ) );
AND2_X1 _13061_ ( .A1(_05317_ ), .A2(_05250_ ), .ZN(_05318_ ) );
INV_X1 _13062_ ( .A(_05318_ ), .ZN(_05319_ ) );
BUF_X4 _13063_ ( .A(_05240_ ), .Z(_05320_ ) );
BUF_X4 _13064_ ( .A(_05320_ ), .Z(_05321_ ) );
BUF_X2 _13065_ ( .A(_05245_ ), .Z(_05322_ ) );
BUF_X2 _13066_ ( .A(_05322_ ), .Z(_05323_ ) );
NAND3_X1 _13067_ ( .A1(_05321_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_05323_ ), .ZN(_05324_ ) );
NAND3_X1 _13068_ ( .A1(_05241_ ), .A2(\mepc [29] ), .A3(_05258_ ), .ZN(_05325_ ) );
BUF_X4 _13069_ ( .A(_05263_ ), .Z(_05326_ ) );
BUF_X4 _13070_ ( .A(_05260_ ), .Z(_05327_ ) );
BUF_X4 _13071_ ( .A(_05327_ ), .Z(_05328_ ) );
NAND4_X1 _13072_ ( .A1(_05326_ ), .A2(_05328_ ), .A3(_05268_ ), .A4(\mtvec [29] ), .ZN(_05329_ ) );
BUF_X2 _13073_ ( .A(_05272_ ), .Z(_05330_ ) );
BUF_X2 _13074_ ( .A(_05330_ ), .Z(_05331_ ) );
NAND4_X1 _13075_ ( .A1(_05331_ ), .A2(_05328_ ), .A3(_05268_ ), .A4(\mycsreg.CSReg[0][29] ), .ZN(_05332_ ) );
AND4_X1 _13076_ ( .A1(_05324_ ), .A2(_05325_ ), .A3(_05329_ ), .A4(_05332_ ), .ZN(_05333_ ) );
NAND3_X1 _13077_ ( .A1(_05315_ ), .A2(_05319_ ), .A3(_05333_ ), .ZN(_05334_ ) );
BUF_X4 _13078_ ( .A(_05310_ ), .Z(_05335_ ) );
INV_X1 _13079_ ( .A(\EX_LS_result_csreg_mem [29] ), .ZN(_05336_ ) );
BUF_X4 _13080_ ( .A(_05312_ ), .Z(_05337_ ) );
AND3_X1 _13081_ ( .A1(_05335_ ), .A2(_05336_ ), .A3(_05337_ ), .ZN(_05338_ ) );
INV_X1 _13082_ ( .A(_05338_ ), .ZN(_05339_ ) );
AND2_X1 _13083_ ( .A1(_05334_ ), .A2(_05339_ ), .ZN(_05340_ ) );
OAI211_X1 _13084_ ( .A(_05301_ ), .B(_05208_ ), .C1(_05211_ ), .C2(_05340_ ), .ZN(_05341_ ) );
MUX2_X1 _13085_ ( .A(_05300_ ), .B(_03047_ ), .S(fanout_net_4 ), .Z(_05342_ ) );
BUF_X2 _13086_ ( .A(_05206_ ), .Z(_05343_ ) );
OR2_X1 _13087_ ( .A1(_05342_ ), .A2(_05343_ ), .ZN(_05344_ ) );
AOI21_X1 _13088_ ( .A(_03907_ ), .B1(_05341_ ), .B2(_05344_ ), .ZN(_00123_ ) );
BUF_X4 _13089_ ( .A(_05207_ ), .Z(_05345_ ) );
OAI21_X1 _13090_ ( .A(_03941_ ), .B1(_03986_ ), .B2(_04005_ ), .ZN(_05346_ ) );
NAND2_X1 _13091_ ( .A1(_05346_ ), .A2(_04016_ ), .ZN(_05347_ ) );
XOR2_X1 _13092_ ( .A(_05347_ ), .B(_03932_ ), .Z(_05348_ ) );
OR3_X1 _13093_ ( .A1(_05198_ ), .A2(_05201_ ), .A3(_05348_ ), .ZN(_05349_ ) );
NAND3_X1 _13094_ ( .A1(_03914_ ), .A2(_05285_ ), .A3(_05288_ ), .ZN(_05350_ ) );
XNOR2_X1 _13095_ ( .A(_05350_ ), .B(\ID_EX_pc [20] ), .ZN(_05351_ ) );
OR2_X1 _13096_ ( .A1(_05203_ ), .A2(_05351_ ), .ZN(_05352_ ) );
AND3_X1 _13097_ ( .A1(_05349_ ), .A2(_05210_ ), .A3(_05352_ ), .ZN(_05353_ ) );
BUF_X2 _13098_ ( .A(_05239_ ), .Z(_05354_ ) );
NAND3_X1 _13099_ ( .A1(_05354_ ), .A2(\mepc [20] ), .A3(_05257_ ), .ZN(_05355_ ) );
BUF_X2 _13100_ ( .A(_05238_ ), .Z(_05356_ ) );
BUF_X4 _13101_ ( .A(_05267_ ), .Z(_05357_ ) );
NAND4_X1 _13102_ ( .A1(_05264_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mtvec [20] ), .ZN(_05358_ ) );
NAND4_X1 _13103_ ( .A1(_05330_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mycsreg.CSReg[0][20] ), .ZN(_05359_ ) );
AND3_X1 _13104_ ( .A1(_05355_ ), .A2(_05358_ ), .A3(_05359_ ), .ZN(_05360_ ) );
NAND3_X1 _13105_ ( .A1(_05241_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_05323_ ), .ZN(_05361_ ) );
AND2_X1 _13106_ ( .A1(_05245_ ), .A2(_05253_ ), .ZN(_05362_ ) );
NAND2_X1 _13107_ ( .A1(_05362_ ), .A2(_05255_ ), .ZN(_05363_ ) );
AND2_X1 _13108_ ( .A1(_05256_ ), .A2(_05363_ ), .ZN(_05364_ ) );
NAND3_X1 _13109_ ( .A1(_05360_ ), .A2(_05361_ ), .A3(_05364_ ), .ZN(_05365_ ) );
OAI21_X1 _13110_ ( .A(_05365_ ), .B1(_05232_ ), .B2(_05231_ ), .ZN(_05366_ ) );
NAND4_X1 _13111_ ( .A1(_05224_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_03840_ ), .A4(_05229_ ), .ZN(_05367_ ) );
AOI21_X1 _13112_ ( .A(_05283_ ), .B1(_05366_ ), .B2(_05367_ ), .ZN(_05368_ ) );
OAI21_X1 _13113_ ( .A(_05345_ ), .B1(_05353_ ), .B2(_05368_ ), .ZN(_05369_ ) );
BUF_X4 _13114_ ( .A(_03887_ ), .Z(_05370_ ) );
AND2_X2 _13115_ ( .A1(_03885_ ), .A2(fanout_net_4 ), .ZN(_05371_ ) );
AOI22_X1 _13116_ ( .A1(_05348_ ), .A2(_05370_ ), .B1(_03017_ ), .B2(_05371_ ), .ZN(_05372_ ) );
AOI21_X1 _13117_ ( .A(_03907_ ), .B1(_05369_ ), .B2(_05372_ ), .ZN(_00124_ ) );
BUF_X2 _13118_ ( .A(_05202_ ), .Z(_05373_ ) );
NAND3_X1 _13119_ ( .A1(_03914_ ), .A2(\ID_EX_pc [18] ), .A3(_05285_ ), .ZN(_05374_ ) );
XNOR2_X1 _13120_ ( .A(_05374_ ), .B(\ID_EX_pc [19] ), .ZN(_05375_ ) );
NOR2_X1 _13121_ ( .A1(_05373_ ), .A2(_05375_ ), .ZN(_05376_ ) );
BUF_X4 _13122_ ( .A(_05203_ ), .Z(_05377_ ) );
NOR2_X1 _13123_ ( .A1(_03986_ ), .A2(_04005_ ), .ZN(_05378_ ) );
NOR2_X1 _13124_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_05379_ ) );
NOR3_X1 _13125_ ( .A1(_05378_ ), .A2(_04012_ ), .A3(_05379_ ), .ZN(_05380_ ) );
AND2_X1 _13126_ ( .A1(_05380_ ), .A2(_03939_ ), .ZN(_05381_ ) );
OAI21_X1 _13127_ ( .A(_03937_ ), .B1(_05381_ ), .B2(_04015_ ), .ZN(_05382_ ) );
NAND2_X1 _13128_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_05383_ ) );
NAND2_X1 _13129_ ( .A1(_05382_ ), .A2(_05383_ ), .ZN(_05384_ ) );
XNOR2_X1 _13130_ ( .A(_05384_ ), .B(_03936_ ), .ZN(_05385_ ) );
AOI211_X1 _13131_ ( .A(\ID_EX_typ [3] ), .B(_05376_ ), .C1(_05377_ ), .C2(_05385_ ), .ZN(_05386_ ) );
BUF_X4 _13132_ ( .A(_05232_ ), .Z(_05387_ ) );
NAND3_X1 _13133_ ( .A1(_05321_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_05323_ ), .ZN(_05388_ ) );
BUF_X4 _13134_ ( .A(_05258_ ), .Z(_05389_ ) );
BUF_X4 _13135_ ( .A(_05328_ ), .Z(_05390_ ) );
NAND4_X1 _13136_ ( .A1(_05389_ ), .A2(_05259_ ), .A3(_05390_ ), .A4(\mepc [19] ), .ZN(_05391_ ) );
BUF_X2 _13137_ ( .A(_05264_ ), .Z(_05392_ ) );
BUF_X4 _13138_ ( .A(_05267_ ), .Z(_05393_ ) );
BUF_X2 _13139_ ( .A(_05393_ ), .Z(_05394_ ) );
NAND4_X1 _13140_ ( .A1(_05392_ ), .A2(_05390_ ), .A3(_05394_ ), .A4(\mtvec [19] ), .ZN(_05395_ ) );
NAND4_X1 _13141_ ( .A1(_05388_ ), .A2(_05363_ ), .A3(_05391_ ), .A4(_05395_ ), .ZN(_05396_ ) );
CLKBUF_X2 _13142_ ( .A(_05273_ ), .Z(_05397_ ) );
AND3_X1 _13143_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_05328_ ), .ZN(_05398_ ) );
OAI22_X1 _13144_ ( .A1(_05231_ ), .A2(_05387_ ), .B1(_05396_ ), .B2(_05398_ ), .ZN(_05399_ ) );
BUF_X4 _13145_ ( .A(_05224_ ), .Z(_05400_ ) );
BUF_X4 _13146_ ( .A(_05229_ ), .Z(_05401_ ) );
NAND4_X1 _13147_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_03841_ ), .A4(_05401_ ), .ZN(_05402_ ) );
AOI21_X1 _13148_ ( .A(_05283_ ), .B1(_05399_ ), .B2(_05402_ ), .ZN(_05403_ ) );
OAI21_X1 _13149_ ( .A(_05345_ ), .B1(_05386_ ), .B2(_05403_ ), .ZN(_05404_ ) );
BUF_X4 _13150_ ( .A(_03886_ ), .Z(_05405_ ) );
BUF_X4 _13151_ ( .A(_05405_ ), .Z(_05406_ ) );
NOR3_X1 _13152_ ( .A1(_03025_ ), .A2(_05406_ ), .A3(_05207_ ), .ZN(_05407_ ) );
INV_X1 _13153_ ( .A(_05385_ ), .ZN(_05408_ ) );
AOI21_X1 _13154_ ( .A(_05407_ ), .B1(_05408_ ), .B2(_05370_ ), .ZN(_05409_ ) );
AOI21_X1 _13155_ ( .A(_03907_ ), .B1(_05404_ ), .B2(_05409_ ), .ZN(_00125_ ) );
INV_X1 _13156_ ( .A(\ID_EX_pc [18] ), .ZN(_05410_ ) );
XNOR2_X1 _13157_ ( .A(_05286_ ), .B(_05410_ ), .ZN(_05411_ ) );
OR3_X1 _13158_ ( .A1(_05381_ ), .A2(_03937_ ), .A3(_04015_ ), .ZN(_05412_ ) );
AND2_X1 _13159_ ( .A1(_05412_ ), .A2(_05382_ ), .ZN(_05413_ ) );
MUX2_X1 _13160_ ( .A(_05411_ ), .B(_05413_ ), .S(_05202_ ), .Z(_05414_ ) );
OR2_X1 _13161_ ( .A1(_05414_ ), .A2(\ID_EX_typ [3] ), .ZN(_05415_ ) );
BUF_X4 _13162_ ( .A(_05207_ ), .Z(_05416_ ) );
BUF_X2 _13163_ ( .A(_05250_ ), .Z(_05417_ ) );
NAND3_X1 _13164_ ( .A1(_05320_ ), .A2(\mepc [18] ), .A3(_05417_ ), .ZN(_05418_ ) );
NAND4_X1 _13165_ ( .A1(_05331_ ), .A2(_05261_ ), .A3(_05393_ ), .A4(\mycsreg.CSReg[0][18] ), .ZN(_05419_ ) );
AND2_X1 _13166_ ( .A1(_05418_ ), .A2(_05419_ ), .ZN(_05420_ ) );
NAND2_X1 _13167_ ( .A1(_05317_ ), .A2(_05245_ ), .ZN(_05421_ ) );
NAND4_X1 _13168_ ( .A1(_05264_ ), .A2(_05327_ ), .A3(_05393_ ), .A4(\mtvec [18] ), .ZN(_05422_ ) );
AND2_X1 _13169_ ( .A1(_05421_ ), .A2(_05422_ ), .ZN(_05423_ ) );
NAND3_X1 _13170_ ( .A1(_05241_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_05323_ ), .ZN(_05424_ ) );
NAND3_X1 _13171_ ( .A1(_05420_ ), .A2(_05423_ ), .A3(_05424_ ), .ZN(_05425_ ) );
OAI21_X1 _13172_ ( .A(_05425_ ), .B1(_05232_ ), .B2(_05231_ ), .ZN(_05426_ ) );
BUF_X4 _13173_ ( .A(_05335_ ), .Z(_05427_ ) );
BUF_X4 _13174_ ( .A(_05337_ ), .Z(_05428_ ) );
NAND3_X1 _13175_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_05428_ ), .ZN(_05429_ ) );
AND2_X1 _13176_ ( .A1(_05426_ ), .A2(_05429_ ), .ZN(_05430_ ) );
INV_X1 _13177_ ( .A(_05430_ ), .ZN(_05431_ ) );
OAI211_X1 _13178_ ( .A(_05415_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05431_ ), .ZN(_05432_ ) );
BUF_X4 _13179_ ( .A(_03886_ ), .Z(_05433_ ) );
NOR4_X1 _13180_ ( .A1(_03026_ ), .A2(_03023_ ), .A3(_05433_ ), .A4(_05206_ ), .ZN(_05434_ ) );
AOI21_X1 _13181_ ( .A(_05434_ ), .B1(_05413_ ), .B2(_05370_ ), .ZN(_05435_ ) );
AOI21_X1 _13182_ ( .A(_03907_ ), .B1(_05432_ ), .B2(_05435_ ), .ZN(_00126_ ) );
BUF_X4 _13183_ ( .A(_05209_ ), .Z(_05436_ ) );
NOR2_X1 _13184_ ( .A1(_05230_ ), .A2(_05232_ ), .ZN(_05437_ ) );
INV_X1 _13185_ ( .A(_05437_ ), .ZN(_05438_ ) );
NAND3_X1 _13186_ ( .A1(_05241_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_05323_ ), .ZN(_05439_ ) );
NAND4_X1 _13187_ ( .A1(_05258_ ), .A2(_05259_ ), .A3(_05328_ ), .A4(\mepc [17] ), .ZN(_05440_ ) );
BUF_X4 _13188_ ( .A(_05393_ ), .Z(_05441_ ) );
NAND4_X1 _13189_ ( .A1(_05326_ ), .A2(_05328_ ), .A3(_05441_ ), .A4(\mtvec [17] ), .ZN(_05442_ ) );
NAND4_X1 _13190_ ( .A1(_05364_ ), .A2(_05439_ ), .A3(_05440_ ), .A4(_05442_ ), .ZN(_05443_ ) );
BUF_X2 _13191_ ( .A(_05261_ ), .Z(_05444_ ) );
AND3_X1 _13192_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_05444_ ), .ZN(_05445_ ) );
OAI21_X1 _13193_ ( .A(_05438_ ), .B1(_05443_ ), .B2(_05445_ ), .ZN(_05446_ ) );
NAND3_X1 _13194_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_05428_ ), .ZN(_05447_ ) );
AND2_X1 _13195_ ( .A1(_05446_ ), .A2(_05447_ ), .ZN(_05448_ ) );
INV_X1 _13196_ ( .A(_05448_ ), .ZN(_05449_ ) );
BUF_X2 _13197_ ( .A(_05203_ ), .Z(_05450_ ) );
NOR2_X1 _13198_ ( .A1(_05380_ ), .A2(_04012_ ), .ZN(_05451_ ) );
XNOR2_X1 _13199_ ( .A(_05451_ ), .B(_03939_ ), .ZN(_05452_ ) );
AND2_X1 _13200_ ( .A1(_05450_ ), .A2(_05452_ ), .ZN(_05453_ ) );
BUF_X4 _13201_ ( .A(_05209_ ), .Z(_05454_ ) );
AND3_X1 _13202_ ( .A1(_03915_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_05455_ ) );
AND2_X1 _13203_ ( .A1(_03914_ ), .A2(_05455_ ), .ZN(_05456_ ) );
NAND3_X1 _13204_ ( .A1(_05456_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05457_ ) );
INV_X1 _13205_ ( .A(\ID_EX_pc [16] ), .ZN(_05458_ ) );
NOR2_X1 _13206_ ( .A1(_05457_ ), .A2(_05458_ ), .ZN(_05459_ ) );
XNOR2_X1 _13207_ ( .A(_05459_ ), .B(\ID_EX_pc [17] ), .ZN(_05460_ ) );
OAI21_X1 _13208_ ( .A(_05454_ ), .B1(_05377_ ), .B2(_05460_ ), .ZN(_05461_ ) );
OAI221_X1 _13209_ ( .A(_05416_ ), .B1(_05436_ ), .B2(_05449_ ), .C1(_05453_ ), .C2(_05461_ ), .ZN(_05462_ ) );
NOR3_X1 _13210_ ( .A1(_03030_ ), .A2(_05406_ ), .A3(_05207_ ), .ZN(_05463_ ) );
AOI21_X1 _13211_ ( .A(_05463_ ), .B1(_05370_ ), .B2(_05452_ ), .ZN(_05464_ ) );
AOI21_X1 _13212_ ( .A(_03907_ ), .B1(_05462_ ), .B2(_05464_ ), .ZN(_00127_ ) );
XNOR2_X1 _13213_ ( .A(_05457_ ), .B(\ID_EX_pc [16] ), .ZN(_05465_ ) );
NOR2_X1 _13214_ ( .A1(_05373_ ), .A2(_05465_ ), .ZN(_05466_ ) );
XNOR2_X1 _13215_ ( .A(_05378_ ), .B(_03940_ ), .ZN(_05467_ ) );
INV_X1 _13216_ ( .A(_05467_ ), .ZN(_05468_ ) );
AOI211_X1 _13217_ ( .A(\ID_EX_typ [3] ), .B(_05466_ ), .C1(_05377_ ), .C2(_05468_ ), .ZN(_05469_ ) );
NAND3_X1 _13218_ ( .A1(_05320_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_05322_ ), .ZN(_05470_ ) );
NAND4_X1 _13219_ ( .A1(_05389_ ), .A2(_05259_ ), .A3(_05390_ ), .A4(\mepc [16] ), .ZN(_05471_ ) );
NAND4_X1 _13220_ ( .A1(_05392_ ), .A2(_05390_ ), .A3(_05394_ ), .A4(\mtvec [16] ), .ZN(_05472_ ) );
NAND4_X1 _13221_ ( .A1(_05364_ ), .A2(_05470_ ), .A3(_05471_ ), .A4(_05472_ ), .ZN(_05473_ ) );
BUF_X4 _13222_ ( .A(_05327_ ), .Z(_05474_ ) );
BUF_X2 _13223_ ( .A(_05474_ ), .Z(_05475_ ) );
AND3_X1 _13224_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_05475_ ), .ZN(_05476_ ) );
OAI22_X1 _13225_ ( .A1(_05473_ ), .A2(_05476_ ), .B1(_05387_ ), .B2(_05231_ ), .ZN(_05477_ ) );
NAND4_X1 _13226_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [16] ), .A3(_03841_ ), .A4(_05401_ ), .ZN(_05478_ ) );
AOI21_X1 _13227_ ( .A(_05283_ ), .B1(_05477_ ), .B2(_05478_ ), .ZN(_05479_ ) );
OAI21_X1 _13228_ ( .A(_05345_ ), .B1(_05469_ ), .B2(_05479_ ), .ZN(_05480_ ) );
AOI22_X1 _13229_ ( .A1(_05467_ ), .A2(_05370_ ), .B1(_03031_ ), .B2(_05371_ ), .ZN(_05481_ ) );
AOI21_X1 _13230_ ( .A(_03907_ ), .B1(_05480_ ), .B2(_05481_ ), .ZN(_00128_ ) );
NAND3_X1 _13231_ ( .A1(_03914_ ), .A2(\ID_EX_pc [14] ), .A3(_05455_ ), .ZN(_05482_ ) );
XNOR2_X1 _13232_ ( .A(_05482_ ), .B(\ID_EX_pc [15] ), .ZN(_05483_ ) );
INV_X1 _13233_ ( .A(_03973_ ), .ZN(_05484_ ) );
OAI21_X1 _13234_ ( .A(_03985_ ), .B1(_03968_ ), .B2(_03969_ ), .ZN(_05485_ ) );
INV_X1 _13235_ ( .A(_03994_ ), .ZN(_05486_ ) );
NAND2_X1 _13236_ ( .A1(_05485_ ), .A2(_05486_ ), .ZN(_05487_ ) );
NAND2_X1 _13237_ ( .A1(_05487_ ), .A2(_03977_ ), .ZN(_05488_ ) );
AOI21_X1 _13238_ ( .A(_05484_ ), .B1(_05488_ ), .B2(_03998_ ), .ZN(_05489_ ) );
NOR2_X1 _13239_ ( .A1(_05489_ ), .A2(_04001_ ), .ZN(_05490_ ) );
XNOR2_X1 _13240_ ( .A(_05490_ ), .B(_03972_ ), .ZN(_05491_ ) );
MUX2_X1 _13241_ ( .A(_05483_ ), .B(_05491_ ), .S(_05202_ ), .Z(_05492_ ) );
OR2_X1 _13242_ ( .A1(_05492_ ), .A2(\ID_EX_typ [3] ), .ZN(_05493_ ) );
AND3_X1 _13243_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_05444_ ), .ZN(_05494_ ) );
NAND3_X1 _13244_ ( .A1(_05321_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_05323_ ), .ZN(_05495_ ) );
NAND4_X1 _13245_ ( .A1(_05258_ ), .A2(_05259_ ), .A3(_05328_ ), .A4(\mepc [15] ), .ZN(_05496_ ) );
NAND4_X1 _13246_ ( .A1(_05326_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mtvec [15] ), .ZN(_05497_ ) );
NAND4_X1 _13247_ ( .A1(_05495_ ), .A2(_05421_ ), .A3(_05496_ ), .A4(_05497_ ), .ZN(_05498_ ) );
OAI21_X1 _13248_ ( .A(_05438_ ), .B1(_05494_ ), .B2(_05498_ ), .ZN(_05499_ ) );
NAND3_X1 _13249_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_05428_ ), .ZN(_05500_ ) );
AND2_X1 _13250_ ( .A1(_05499_ ), .A2(_05500_ ), .ZN(_05501_ ) );
INV_X1 _13251_ ( .A(_05501_ ), .ZN(_05502_ ) );
OAI211_X1 _13252_ ( .A(_05493_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05502_ ), .ZN(_05503_ ) );
NOR3_X1 _13253_ ( .A1(_03038_ ), .A2(_05406_ ), .A3(_05206_ ), .ZN(_05504_ ) );
AOI21_X1 _13254_ ( .A(_05504_ ), .B1(_05370_ ), .B2(_05491_ ), .ZN(_05505_ ) );
AOI21_X1 _13255_ ( .A(_03907_ ), .B1(_05503_ ), .B2(_05505_ ), .ZN(_00129_ ) );
BUF_X4 _13256_ ( .A(_05207_ ), .Z(_05506_ ) );
BUF_X2 _13257_ ( .A(_05240_ ), .Z(_05507_ ) );
NAND3_X1 _13258_ ( .A1(_05507_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_05246_ ), .ZN(_05508_ ) );
NAND3_X1 _13259_ ( .A1(_05320_ ), .A2(\mepc [14] ), .A3(_05417_ ), .ZN(_05509_ ) );
NAND4_X1 _13260_ ( .A1(_05331_ ), .A2(_05261_ ), .A3(_05393_ ), .A4(\mycsreg.CSReg[0][14] ), .ZN(_05510_ ) );
AND3_X1 _13261_ ( .A1(_05508_ ), .A2(_05509_ ), .A3(_05510_ ), .ZN(_05511_ ) );
AND2_X1 _13262_ ( .A1(_05317_ ), .A2(_05245_ ), .ZN(_05512_ ) );
NOR2_X1 _13263_ ( .A1(_05318_ ), .A2(_05512_ ), .ZN(_05513_ ) );
NAND4_X1 _13264_ ( .A1(_05392_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mtvec [14] ), .ZN(_05514_ ) );
NAND3_X1 _13265_ ( .A1(_05511_ ), .A2(_05513_ ), .A3(_05514_ ), .ZN(_05515_ ) );
NAND2_X1 _13266_ ( .A1(_05315_ ), .A2(_05515_ ), .ZN(_05516_ ) );
NAND3_X1 _13267_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [14] ), .A3(_05428_ ), .ZN(_05517_ ) );
AND2_X1 _13268_ ( .A1(_05516_ ), .A2(_05517_ ), .ZN(_05518_ ) );
INV_X1 _13269_ ( .A(_05518_ ), .ZN(_05519_ ) );
AOI211_X1 _13270_ ( .A(_03973_ ), .B(_03999_ ), .C1(_05487_ ), .C2(_03977_ ), .ZN(_05520_ ) );
NOR2_X1 _13271_ ( .A1(_05489_ ), .A2(_05520_ ), .ZN(_05521_ ) );
AND2_X1 _13272_ ( .A1(_05450_ ), .A2(_05521_ ), .ZN(_05522_ ) );
XNOR2_X1 _13273_ ( .A(_05456_ ), .B(\ID_EX_pc [14] ), .ZN(_05523_ ) );
OAI21_X1 _13274_ ( .A(_05454_ ), .B1(_05377_ ), .B2(_05523_ ), .ZN(_05524_ ) );
OAI221_X1 _13275_ ( .A(_05506_ ), .B1(_05436_ ), .B2(_05519_ ), .C1(_05522_ ), .C2(_05524_ ), .ZN(_05525_ ) );
AND3_X1 _13276_ ( .A1(_03039_ ), .A2(_03036_ ), .A3(_05371_ ), .ZN(_05526_ ) );
AOI21_X1 _13277_ ( .A(_05526_ ), .B1(_05370_ ), .B2(_05521_ ), .ZN(_05527_ ) );
AOI21_X1 _13278_ ( .A(_03907_ ), .B1(_05525_ ), .B2(_05527_ ), .ZN(_00130_ ) );
BUF_X4 _13279_ ( .A(_03906_ ), .Z(_05528_ ) );
AND3_X1 _13280_ ( .A1(_05507_ ), .A2(\mepc [13] ), .A3(_05417_ ), .ZN(_05529_ ) );
INV_X1 _13281_ ( .A(_05529_ ), .ZN(_05530_ ) );
AND3_X1 _13282_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_05261_ ), .ZN(_05531_ ) );
INV_X1 _13283_ ( .A(_05531_ ), .ZN(_05532_ ) );
AND4_X1 _13284_ ( .A1(_02128_ ), .A2(_05225_ ), .A3(_05226_ ), .A4(_05227_ ), .ZN(_05533_ ) );
NAND3_X1 _13285_ ( .A1(_05533_ ), .A2(_05214_ ), .A3(_05217_ ), .ZN(_05534_ ) );
NAND3_X1 _13286_ ( .A1(_05220_ ), .A2(_05223_ ), .A3(_05228_ ), .ZN(_05535_ ) );
BUF_X2 _13287_ ( .A(_05535_ ), .Z(_05536_ ) );
OAI211_X1 _13288_ ( .A(_05530_ ), .B(_05532_ ), .C1(_05534_ ), .C2(_05536_ ), .ZN(_05537_ ) );
AND3_X1 _13289_ ( .A1(_05507_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_05246_ ), .ZN(_05538_ ) );
INV_X1 _13290_ ( .A(_05538_ ), .ZN(_05539_ ) );
AND2_X1 _13291_ ( .A1(_05255_ ), .A2(_05253_ ), .ZN(_05540_ ) );
AND2_X1 _13292_ ( .A1(_05540_ ), .A2(_05257_ ), .ZN(_05541_ ) );
INV_X1 _13293_ ( .A(_05541_ ), .ZN(_05542_ ) );
AND4_X2 _13294_ ( .A1(_05248_ ), .A2(_05267_ ), .A3(\ID_EX_csr [0] ), .A4(_05242_ ), .ZN(_05543_ ) );
NAND4_X1 _13295_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [13] ), .A4(_05444_ ), .ZN(_05544_ ) );
NAND3_X1 _13296_ ( .A1(_05539_ ), .A2(_05542_ ), .A3(_05544_ ), .ZN(_05545_ ) );
NOR2_X1 _13297_ ( .A1(_05537_ ), .A2(_05545_ ), .ZN(_05546_ ) );
BUF_X2 _13298_ ( .A(_05534_ ), .Z(_05547_ ) );
NOR3_X1 _13299_ ( .A1(_05547_ ), .A2(\EX_LS_result_csreg_mem [13] ), .A3(_05536_ ), .ZN(_05548_ ) );
NOR2_X1 _13300_ ( .A1(_05546_ ), .A2(_05548_ ), .ZN(_05549_ ) );
INV_X1 _13301_ ( .A(_03975_ ), .ZN(_05550_ ) );
AOI21_X1 _13302_ ( .A(_05550_ ), .B1(_05485_ ), .B2(_05486_ ), .ZN(_05551_ ) );
NOR2_X1 _13303_ ( .A1(_05551_ ), .A2(_03997_ ), .ZN(_05552_ ) );
XNOR2_X1 _13304_ ( .A(_05552_ ), .B(_03976_ ), .ZN(_05553_ ) );
AND2_X1 _13305_ ( .A1(_05450_ ), .A2(_05553_ ), .ZN(_05554_ ) );
AND2_X1 _13306_ ( .A1(_03916_ ), .A2(\ID_EX_pc [12] ), .ZN(_05555_ ) );
XNOR2_X1 _13307_ ( .A(_05555_ ), .B(\ID_EX_pc [13] ), .ZN(_05556_ ) );
OAI21_X1 _13308_ ( .A(_05454_ ), .B1(_05377_ ), .B2(_05556_ ), .ZN(_05557_ ) );
OAI221_X1 _13309_ ( .A(_05506_ ), .B1(_05436_ ), .B2(_05549_ ), .C1(_05554_ ), .C2(_05557_ ), .ZN(_05558_ ) );
NOR3_X1 _13310_ ( .A1(_03042_ ), .A2(_05406_ ), .A3(_05206_ ), .ZN(_05559_ ) );
AOI21_X1 _13311_ ( .A(_05559_ ), .B1(_05370_ ), .B2(_05553_ ), .ZN(_05560_ ) );
AOI21_X1 _13312_ ( .A(_05528_ ), .B1(_05558_ ), .B2(_05560_ ), .ZN(_00131_ ) );
INV_X1 _13313_ ( .A(\ID_EX_pc [12] ), .ZN(_05561_ ) );
XNOR2_X1 _13314_ ( .A(_03916_ ), .B(_05561_ ), .ZN(_05562_ ) );
XNOR2_X1 _13315_ ( .A(_05487_ ), .B(_05550_ ), .ZN(_05563_ ) );
MUX2_X1 _13316_ ( .A(_05562_ ), .B(_05563_ ), .S(_05202_ ), .Z(_05564_ ) );
OR2_X1 _13317_ ( .A1(_05564_ ), .A2(\ID_EX_typ [3] ), .ZN(_05565_ ) );
NAND3_X1 _13318_ ( .A1(_05320_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_05322_ ), .ZN(_05566_ ) );
NAND3_X1 _13319_ ( .A1(_05354_ ), .A2(\mepc [12] ), .A3(_05417_ ), .ZN(_05567_ ) );
NAND4_X1 _13320_ ( .A1(_05330_ ), .A2(_05327_ ), .A3(_05393_ ), .A4(\mycsreg.CSReg[0][12] ), .ZN(_05568_ ) );
AND3_X1 _13321_ ( .A1(_05566_ ), .A2(_05567_ ), .A3(_05568_ ), .ZN(_05569_ ) );
NAND4_X1 _13322_ ( .A1(_05326_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mtvec [12] ), .ZN(_05570_ ) );
NAND3_X1 _13323_ ( .A1(_05569_ ), .A2(_05513_ ), .A3(_05570_ ), .ZN(_05571_ ) );
NAND2_X1 _13324_ ( .A1(_05314_ ), .A2(_05571_ ), .ZN(_05572_ ) );
NAND3_X1 _13325_ ( .A1(_05335_ ), .A2(\EX_LS_result_csreg_mem [12] ), .A3(_05337_ ), .ZN(_05573_ ) );
AND2_X1 _13326_ ( .A1(_05572_ ), .A2(_05573_ ), .ZN(_05574_ ) );
INV_X1 _13327_ ( .A(_05574_ ), .ZN(_05575_ ) );
OAI211_X1 _13328_ ( .A(_05565_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05575_ ), .ZN(_05576_ ) );
BUF_X4 _13329_ ( .A(_05371_ ), .Z(_05577_ ) );
BUF_X4 _13330_ ( .A(_03887_ ), .Z(_05578_ ) );
AOI22_X1 _13331_ ( .A1(_03043_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05563_ ), .ZN(_05579_ ) );
AOI21_X1 _13332_ ( .A(_05528_ ), .B1(_05576_ ), .B2(_05579_ ), .ZN(_00132_ ) );
NAND3_X1 _13333_ ( .A1(_05507_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_05246_ ), .ZN(_05580_ ) );
NAND3_X1 _13334_ ( .A1(_05320_ ), .A2(\mepc [11] ), .A3(_05417_ ), .ZN(_05581_ ) );
NAND4_X1 _13335_ ( .A1(_05331_ ), .A2(_05327_ ), .A3(_05393_ ), .A4(\mycsreg.CSReg[0][11] ), .ZN(_05582_ ) );
AND3_X1 _13336_ ( .A1(_05580_ ), .A2(_05581_ ), .A3(_05582_ ), .ZN(_05583_ ) );
NAND4_X1 _13337_ ( .A1(_05392_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mtvec [11] ), .ZN(_05584_ ) );
NAND3_X1 _13338_ ( .A1(_05583_ ), .A2(_05513_ ), .A3(_05584_ ), .ZN(_05585_ ) );
NAND2_X1 _13339_ ( .A1(_05315_ ), .A2(_05585_ ), .ZN(_05586_ ) );
NAND3_X1 _13340_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [11] ), .A3(_05428_ ), .ZN(_05587_ ) );
AND2_X1 _13341_ ( .A1(_05586_ ), .A2(_05587_ ), .ZN(_05588_ ) );
INV_X1 _13342_ ( .A(_05588_ ), .ZN(_05589_ ) );
INV_X1 _13343_ ( .A(_03980_ ), .ZN(_05590_ ) );
OAI21_X1 _13344_ ( .A(_03984_ ), .B1(_03968_ ), .B2(_03969_ ), .ZN(_05591_ ) );
AOI21_X1 _13345_ ( .A(_05590_ ), .B1(_05591_ ), .B2(_03992_ ), .ZN(_05592_ ) );
NOR2_X1 _13346_ ( .A1(_05592_ ), .A2(_03987_ ), .ZN(_05593_ ) );
XNOR2_X1 _13347_ ( .A(_05593_ ), .B(_03979_ ), .ZN(_05594_ ) );
AND2_X1 _13348_ ( .A1(_05450_ ), .A2(_05594_ ), .ZN(_05595_ ) );
AND2_X1 _13349_ ( .A1(_03914_ ), .A2(\ID_EX_pc [10] ), .ZN(_05596_ ) );
XNOR2_X1 _13350_ ( .A(_05596_ ), .B(\ID_EX_pc [11] ), .ZN(_05597_ ) );
OAI21_X1 _13351_ ( .A(_05454_ ), .B1(_05450_ ), .B2(_05597_ ), .ZN(_05598_ ) );
OAI221_X1 _13352_ ( .A(_05506_ ), .B1(_05436_ ), .B2(_05589_ ), .C1(_05595_ ), .C2(_05598_ ), .ZN(_05599_ ) );
NAND2_X1 _13353_ ( .A1(_02869_ ), .A2(_02877_ ), .ZN(_05600_ ) );
AOI21_X1 _13354_ ( .A(_02884_ ), .B1(_05600_ ), .B2(_02626_ ), .ZN(_05601_ ) );
AND3_X1 _13355_ ( .A1(_02645_ ), .A2(_02648_ ), .A3(_02646_ ), .ZN(_05602_ ) );
NOR3_X1 _13356_ ( .A1(_05601_ ), .A2(_02879_ ), .A3(_05602_ ), .ZN(_05603_ ) );
NOR2_X1 _13357_ ( .A1(_05603_ ), .A2(_02879_ ), .ZN(_05604_ ) );
XNOR2_X1 _13358_ ( .A(_05604_ ), .B(_02672_ ), .ZN(_05605_ ) );
AOI22_X1 _13359_ ( .A1(_05605_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05594_ ), .ZN(_05606_ ) );
AOI21_X1 _13360_ ( .A(_05528_ ), .B1(_05599_ ), .B2(_05606_ ), .ZN(_00133_ ) );
INV_X1 _13361_ ( .A(\ID_EX_pc [28] ), .ZN(_05607_ ) );
XNOR2_X1 _13362_ ( .A(_05293_ ), .B(_05607_ ), .ZN(_05608_ ) );
OAI21_X1 _13363_ ( .A(_05608_ ), .B1(_05198_ ), .B2(_05201_ ), .ZN(_05609_ ) );
XNOR2_X1 _13364_ ( .A(_04035_ ), .B(_04036_ ), .ZN(_05610_ ) );
OAI211_X1 _13365_ ( .A(_05283_ ), .B(_05609_ ), .C1(_05297_ ), .C2(_05610_ ), .ZN(_05611_ ) );
NAND3_X1 _13366_ ( .A1(_05321_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_05323_ ), .ZN(_05612_ ) );
NAND3_X1 _13367_ ( .A1(_05241_ ), .A2(\mepc [28] ), .A3(_05258_ ), .ZN(_05613_ ) );
NAND4_X1 _13368_ ( .A1(_05331_ ), .A2(_05328_ ), .A3(_05268_ ), .A4(\mycsreg.CSReg[0][28] ), .ZN(_05614_ ) );
NAND4_X1 _13369_ ( .A1(_05326_ ), .A2(_05265_ ), .A3(_05268_ ), .A4(\mtvec [28] ), .ZN(_05615_ ) );
AND4_X1 _13370_ ( .A1(_05612_ ), .A2(_05613_ ), .A3(_05614_ ), .A4(_05615_ ), .ZN(_05616_ ) );
NAND3_X1 _13371_ ( .A1(_05315_ ), .A2(_05319_ ), .A3(_05616_ ), .ZN(_05617_ ) );
INV_X1 _13372_ ( .A(\EX_LS_result_csreg_mem [28] ), .ZN(_05618_ ) );
AND3_X1 _13373_ ( .A1(_05335_ ), .A2(_05618_ ), .A3(_05337_ ), .ZN(_05619_ ) );
INV_X1 _13374_ ( .A(_05619_ ), .ZN(_05620_ ) );
AND2_X1 _13375_ ( .A1(_05617_ ), .A2(_05620_ ), .ZN(_05621_ ) );
OAI211_X1 _13376_ ( .A(_05611_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05621_ ), .ZN(_05622_ ) );
BUF_X4 _13377_ ( .A(_05405_ ), .Z(_05623_ ) );
AOI21_X1 _13378_ ( .A(_05207_ ), .B1(_05610_ ), .B2(_05623_ ), .ZN(_05624_ ) );
OAI21_X1 _13379_ ( .A(_05624_ ), .B1(_03048_ ), .B2(_05623_ ), .ZN(_05625_ ) );
AOI21_X1 _13380_ ( .A(_05528_ ), .B1(_05622_ ), .B2(_05625_ ), .ZN(_00134_ ) );
INV_X1 _13381_ ( .A(\ID_EX_pc [10] ), .ZN(_05626_ ) );
XNOR2_X1 _13382_ ( .A(_03914_ ), .B(_05626_ ), .ZN(_05627_ ) );
AND3_X1 _13383_ ( .A1(_05591_ ), .A2(_05590_ ), .A3(_03992_ ), .ZN(_05628_ ) );
NOR2_X1 _13384_ ( .A1(_05628_ ), .A2(_05592_ ), .ZN(_05629_ ) );
MUX2_X1 _13385_ ( .A(_05627_ ), .B(_05629_ ), .S(_05203_ ), .Z(_05630_ ) );
AND2_X1 _13386_ ( .A1(_05630_ ), .A2(_05210_ ), .ZN(_05631_ ) );
NAND3_X1 _13387_ ( .A1(_05354_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_05322_ ), .ZN(_05632_ ) );
NAND4_X1 _13388_ ( .A1(_05257_ ), .A2(_05235_ ), .A3(_05260_ ), .A4(\mepc [10] ), .ZN(_05633_ ) );
AND3_X1 _13389_ ( .A1(_05632_ ), .A2(_05363_ ), .A3(_05633_ ), .ZN(_05634_ ) );
NAND4_X1 _13390_ ( .A1(_05326_ ), .A2(_05328_ ), .A3(_05441_ ), .A4(\mtvec [10] ), .ZN(_05635_ ) );
NAND2_X1 _13391_ ( .A1(_05634_ ), .A2(_05635_ ), .ZN(_05636_ ) );
AND3_X1 _13392_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][10] ), .A3(_05328_ ), .ZN(_05637_ ) );
OAI21_X1 _13393_ ( .A(_05438_ ), .B1(_05636_ ), .B2(_05637_ ), .ZN(_05638_ ) );
NAND4_X1 _13394_ ( .A1(_05224_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_03840_ ), .A4(_05229_ ), .ZN(_05639_ ) );
AOI21_X1 _13395_ ( .A(_05283_ ), .B1(_05638_ ), .B2(_05639_ ), .ZN(_05640_ ) );
OAI21_X1 _13396_ ( .A(_05345_ ), .B1(_05631_ ), .B2(_05640_ ), .ZN(_05641_ ) );
XNOR2_X1 _13397_ ( .A(_05601_ ), .B(_02649_ ), .ZN(_05642_ ) );
AOI22_X1 _13398_ ( .A1(_05642_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05629_ ), .ZN(_05643_ ) );
AOI21_X1 _13399_ ( .A(_05528_ ), .B1(_05641_ ), .B2(_05643_ ), .ZN(_00135_ ) );
NAND3_X1 _13400_ ( .A1(_05240_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_05245_ ), .ZN(_05644_ ) );
NAND3_X1 _13401_ ( .A1(_05240_ ), .A2(\mepc [9] ), .A3(_05257_ ), .ZN(_05645_ ) );
NAND4_X1 _13402_ ( .A1(_05330_ ), .A2(_05260_ ), .A3(_05267_ ), .A4(\mycsreg.CSReg[0][9] ), .ZN(_05646_ ) );
NAND3_X1 _13403_ ( .A1(_05644_ ), .A2(_05645_ ), .A3(_05646_ ), .ZN(_05647_ ) );
NAND4_X1 _13404_ ( .A1(_05263_ ), .A2(_05260_ ), .A3(_05267_ ), .A4(\mtvec [9] ), .ZN(_05648_ ) );
NAND2_X1 _13405_ ( .A1(_05421_ ), .A2(_05648_ ), .ZN(_05649_ ) );
OAI21_X1 _13406_ ( .A(_05314_ ), .B1(_05647_ ), .B2(_05649_ ), .ZN(_05650_ ) );
NAND3_X1 _13407_ ( .A1(_05310_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_05312_ ), .ZN(_05651_ ) );
AND2_X1 _13408_ ( .A1(_05650_ ), .A2(_05651_ ), .ZN(_05652_ ) );
INV_X1 _13409_ ( .A(_05652_ ), .ZN(_05653_ ) );
AND2_X1 _13410_ ( .A1(_03971_ ), .A2(_03982_ ), .ZN(_05654_ ) );
NOR2_X1 _13411_ ( .A1(_05654_ ), .A2(_03990_ ), .ZN(_05655_ ) );
XNOR2_X1 _13412_ ( .A(_05655_ ), .B(_03983_ ), .ZN(_05656_ ) );
AND2_X1 _13413_ ( .A1(_05373_ ), .A2(_05656_ ), .ZN(_05657_ ) );
XNOR2_X1 _13414_ ( .A(_03913_ ), .B(\ID_EX_pc [9] ), .ZN(_05658_ ) );
OAI21_X1 _13415_ ( .A(_05454_ ), .B1(_05450_ ), .B2(_05658_ ), .ZN(_05659_ ) );
OAI221_X1 _13416_ ( .A(_05506_ ), .B1(_05436_ ), .B2(_05653_ ), .C1(_05657_ ), .C2(_05659_ ), .ZN(_05660_ ) );
NAND2_X1 _13417_ ( .A1(_05600_ ), .A2(_02602_ ), .ZN(_05661_ ) );
AND2_X1 _13418_ ( .A1(_05661_ ), .A2(_02883_ ), .ZN(_05662_ ) );
XNOR2_X1 _13419_ ( .A(_05662_ ), .B(_02625_ ), .ZN(_05663_ ) );
NOR3_X1 _13420_ ( .A1(_05663_ ), .A2(_05406_ ), .A3(_05206_ ), .ZN(_05664_ ) );
AOI21_X1 _13421_ ( .A(_05664_ ), .B1(_05370_ ), .B2(_05656_ ), .ZN(_05665_ ) );
AOI21_X1 _13422_ ( .A(_05528_ ), .B1(_05660_ ), .B2(_05665_ ), .ZN(_00136_ ) );
NAND3_X1 _13423_ ( .A1(_05240_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_05245_ ), .ZN(_05666_ ) );
NAND3_X1 _13424_ ( .A1(_05240_ ), .A2(\mepc [8] ), .A3(_05257_ ), .ZN(_05667_ ) );
NAND4_X1 _13425_ ( .A1(_05330_ ), .A2(_05260_ ), .A3(_05267_ ), .A4(\mycsreg.CSReg[0][8] ), .ZN(_05668_ ) );
AND3_X1 _13426_ ( .A1(_05666_ ), .A2(_05667_ ), .A3(_05668_ ), .ZN(_05669_ ) );
NAND4_X1 _13427_ ( .A1(_05326_ ), .A2(_05265_ ), .A3(_05268_ ), .A4(\mtvec [8] ), .ZN(_05670_ ) );
NAND3_X1 _13428_ ( .A1(_05669_ ), .A2(_05513_ ), .A3(_05670_ ), .ZN(_05671_ ) );
OAI21_X1 _13429_ ( .A(_05671_ ), .B1(_05232_ ), .B2(_05230_ ), .ZN(_05672_ ) );
NAND3_X1 _13430_ ( .A1(_05335_ ), .A2(\EX_LS_result_csreg_mem [8] ), .A3(_05337_ ), .ZN(_05673_ ) );
AND2_X1 _13431_ ( .A1(_05672_ ), .A2(_05673_ ), .ZN(_05674_ ) );
INV_X1 _13432_ ( .A(_05674_ ), .ZN(_05675_ ) );
XNOR2_X1 _13433_ ( .A(_03970_ ), .B(_03982_ ), .ZN(_05676_ ) );
AND2_X1 _13434_ ( .A1(_05373_ ), .A2(_05676_ ), .ZN(_05677_ ) );
XNOR2_X1 _13435_ ( .A(_03912_ ), .B(\ID_EX_pc [8] ), .ZN(_05678_ ) );
OAI21_X1 _13436_ ( .A(_05454_ ), .B1(_05450_ ), .B2(_05678_ ), .ZN(_05679_ ) );
OAI221_X1 _13437_ ( .A(_05506_ ), .B1(_05436_ ), .B2(_05675_ ), .C1(_05677_ ), .C2(_05679_ ), .ZN(_05680_ ) );
XNOR2_X1 _13438_ ( .A(_05600_ ), .B(_02603_ ), .ZN(_05681_ ) );
AOI22_X1 _13439_ ( .A1(_05681_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05676_ ), .ZN(_05682_ ) );
AOI21_X1 _13440_ ( .A(_05528_ ), .B1(_05680_ ), .B2(_05682_ ), .ZN(_00137_ ) );
AND3_X1 _13441_ ( .A1(_05320_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_05246_ ), .ZN(_05683_ ) );
AND4_X1 _13442_ ( .A1(\mycsreg.CSReg[0][7] ), .A2(_05330_ ), .A3(_05356_ ), .A4(_05393_ ), .ZN(_05684_ ) );
NOR2_X1 _13443_ ( .A1(_05683_ ), .A2(_05684_ ), .ZN(_05685_ ) );
NAND3_X1 _13444_ ( .A1(_05507_ ), .A2(\mepc [7] ), .A3(_05417_ ), .ZN(_05686_ ) );
NAND4_X1 _13445_ ( .A1(_05264_ ), .A2(_05261_ ), .A3(_05393_ ), .A4(\mtvec [7] ), .ZN(_05687_ ) );
AND2_X1 _13446_ ( .A1(_05686_ ), .A2(_05687_ ), .ZN(_05688_ ) );
OAI211_X1 _13447_ ( .A(_05685_ ), .B(_05688_ ), .C1(_05534_ ), .C2(_05535_ ), .ZN(_05689_ ) );
OR3_X1 _13448_ ( .A1(_05534_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_05535_ ), .ZN(_05690_ ) );
NAND2_X1 _13449_ ( .A1(_05689_ ), .A2(_05690_ ), .ZN(_05691_ ) );
INV_X1 _13450_ ( .A(_05691_ ), .ZN(_05692_ ) );
NOR2_X1 _13451_ ( .A1(_03969_ ), .A2(_03967_ ), .ZN(_05693_ ) );
XNOR2_X1 _13452_ ( .A(_03966_ ), .B(_05693_ ), .ZN(_05694_ ) );
AND2_X1 _13453_ ( .A1(_05373_ ), .A2(_05694_ ), .ZN(_05695_ ) );
XNOR2_X1 _13454_ ( .A(_03911_ ), .B(\ID_EX_pc [7] ), .ZN(_05696_ ) );
OAI21_X1 _13455_ ( .A(_05210_ ), .B1(_05450_ ), .B2(_05696_ ), .ZN(_05697_ ) );
OAI221_X1 _13456_ ( .A(_05506_ ), .B1(_05436_ ), .B2(_05692_ ), .C1(_05695_ ), .C2(_05697_ ), .ZN(_05698_ ) );
AND2_X1 _13457_ ( .A1(_02771_ ), .A2(_02868_ ), .ZN(_05699_ ) );
NOR2_X1 _13458_ ( .A1(_05699_ ), .A2(_02876_ ), .ZN(_05700_ ) );
NOR2_X1 _13459_ ( .A1(_05700_ ), .A2(_02795_ ), .ZN(_05701_ ) );
AND2_X1 _13460_ ( .A1(_02792_ ), .A2(\ID_EX_imm [6] ), .ZN(_05702_ ) );
OR2_X1 _13461_ ( .A1(_05701_ ), .A2(_05702_ ), .ZN(_05703_ ) );
XNOR2_X1 _13462_ ( .A(_05703_ ), .B(_02817_ ), .ZN(_05704_ ) );
AOI22_X1 _13463_ ( .A1(_05704_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05694_ ), .ZN(_05705_ ) );
AOI21_X1 _13464_ ( .A(_05528_ ), .B1(_05698_ ), .B2(_05705_ ), .ZN(_00138_ ) );
XOR2_X1 _13465_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_05706_ ) );
XNOR2_X1 _13466_ ( .A(_03962_ ), .B(_05706_ ), .ZN(_05707_ ) );
NAND2_X1 _13467_ ( .A1(_05373_ ), .A2(_05707_ ), .ZN(_05708_ ) );
INV_X1 _13468_ ( .A(\ID_EX_pc [6] ), .ZN(_05709_ ) );
XNOR2_X1 _13469_ ( .A(_03910_ ), .B(_05709_ ), .ZN(_05710_ ) );
OAI21_X1 _13470_ ( .A(_05710_ ), .B1(_05198_ ), .B2(_05201_ ), .ZN(_05711_ ) );
NAND3_X1 _13471_ ( .A1(_05708_ ), .A2(_05436_ ), .A3(_05711_ ), .ZN(_05712_ ) );
NAND3_X1 _13472_ ( .A1(_05320_ ), .A2(\mepc [6] ), .A3(_05417_ ), .ZN(_05713_ ) );
NAND3_X1 _13473_ ( .A1(_05354_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_05322_ ), .ZN(_05714_ ) );
NAND4_X1 _13474_ ( .A1(_05330_ ), .A2(_05327_ ), .A3(_05357_ ), .A4(\mycsreg.CSReg[0][6] ), .ZN(_05715_ ) );
NAND4_X1 _13475_ ( .A1(_05264_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mtvec [6] ), .ZN(_05716_ ) );
NAND4_X1 _13476_ ( .A1(_05713_ ), .A2(_05714_ ), .A3(_05715_ ), .A4(_05716_ ), .ZN(_05717_ ) );
AOI211_X1 _13477_ ( .A(_05318_ ), .B(_05717_ ), .C1(_05335_ ), .C2(_05337_ ), .ZN(_05718_ ) );
INV_X1 _13478_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_05719_ ) );
AND3_X1 _13479_ ( .A1(_05335_ ), .A2(_05719_ ), .A3(_05337_ ), .ZN(_05720_ ) );
NOR2_X1 _13480_ ( .A1(_05718_ ), .A2(_05720_ ), .ZN(_05721_ ) );
OAI211_X1 _13481_ ( .A(_05712_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05721_ ), .ZN(_05722_ ) );
XNOR2_X1 _13482_ ( .A(_05700_ ), .B(_02794_ ), .ZN(_05723_ ) );
AOI22_X1 _13483_ ( .A1(_05723_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05707_ ), .ZN(_05724_ ) );
AOI21_X1 _13484_ ( .A(_05528_ ), .B1(_05722_ ), .B2(_05724_ ), .ZN(_00139_ ) );
XOR2_X1 _13485_ ( .A(_03909_ ), .B(\ID_EX_pc [5] ), .Z(_05725_ ) );
NOR2_X1 _13486_ ( .A1(_03961_ ), .A2(_03959_ ), .ZN(_05726_ ) );
XNOR2_X1 _13487_ ( .A(_03958_ ), .B(_05726_ ), .ZN(_05727_ ) );
MUX2_X1 _13488_ ( .A(_05725_ ), .B(_05727_ ), .S(_05203_ ), .Z(_05728_ ) );
AND2_X1 _13489_ ( .A1(_05728_ ), .A2(_05210_ ), .ZN(_05729_ ) );
NAND3_X1 _13490_ ( .A1(_05241_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_05246_ ), .ZN(_05730_ ) );
NAND4_X1 _13491_ ( .A1(_05389_ ), .A2(_05259_ ), .A3(_05390_ ), .A4(\mepc [5] ), .ZN(_05731_ ) );
NAND4_X1 _13492_ ( .A1(_05392_ ), .A2(_05390_ ), .A3(_05394_ ), .A4(\mtvec [5] ), .ZN(_05732_ ) );
NAND4_X1 _13493_ ( .A1(_05730_ ), .A2(_05256_ ), .A3(_05731_ ), .A4(_05732_ ), .ZN(_05733_ ) );
AND3_X1 _13494_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_05265_ ), .ZN(_05734_ ) );
OAI22_X1 _13495_ ( .A1(_05231_ ), .A2(_05387_ ), .B1(_05733_ ), .B2(_05734_ ), .ZN(_05735_ ) );
BUF_X4 _13496_ ( .A(_03840_ ), .Z(_05736_ ) );
NAND4_X1 _13497_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [5] ), .A3(_05736_ ), .A4(_05401_ ), .ZN(_05737_ ) );
AOI21_X1 _13498_ ( .A(_05283_ ), .B1(_05735_ ), .B2(_05737_ ), .ZN(_05738_ ) );
OAI21_X1 _13499_ ( .A(_05345_ ), .B1(_05729_ ), .B2(_05738_ ), .ZN(_05739_ ) );
AOI21_X1 _13500_ ( .A(_02872_ ), .B1(_02771_ ), .B2(_02866_ ), .ZN(_05740_ ) );
XOR2_X1 _13501_ ( .A(_05740_ ), .B(_02842_ ), .Z(_05741_ ) );
AOI22_X1 _13502_ ( .A1(_05741_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05727_ ), .ZN(_05742_ ) );
AOI21_X1 _13503_ ( .A(_05528_ ), .B1(_05739_ ), .B2(_05742_ ), .ZN(_00140_ ) );
BUF_X4 _13504_ ( .A(_03906_ ), .Z(_05743_ ) );
NOR2_X1 _13505_ ( .A1(_05534_ ), .A2(_05535_ ), .ZN(_05744_ ) );
INV_X1 _13506_ ( .A(_05744_ ), .ZN(_05745_ ) );
NAND4_X1 _13507_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [4] ), .A4(_05474_ ), .ZN(_05746_ ) );
AND3_X1 _13508_ ( .A1(_05354_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_05322_ ), .ZN(_05747_ ) );
NOR2_X1 _13509_ ( .A1(_05747_ ), .A2(_05541_ ), .ZN(_05748_ ) );
AND3_X1 _13510_ ( .A1(_05354_ ), .A2(\mepc [4] ), .A3(_05257_ ), .ZN(_05749_ ) );
AND3_X1 _13511_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_05327_ ), .ZN(_05750_ ) );
NOR2_X1 _13512_ ( .A1(_05749_ ), .A2(_05750_ ), .ZN(_05751_ ) );
NAND4_X1 _13513_ ( .A1(_05745_ ), .A2(_05746_ ), .A3(_05748_ ), .A4(_05751_ ), .ZN(_05752_ ) );
OR3_X1 _13514_ ( .A1(_05534_ ), .A2(\EX_LS_result_csreg_mem [4] ), .A3(_05535_ ), .ZN(_05753_ ) );
AND2_X1 _13515_ ( .A1(_05752_ ), .A2(_05753_ ), .ZN(_05754_ ) );
XOR2_X1 _13516_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_05755_ ) );
XNOR2_X1 _13517_ ( .A(_03954_ ), .B(_05755_ ), .ZN(_05756_ ) );
AND2_X1 _13518_ ( .A1(_05373_ ), .A2(_05756_ ), .ZN(_05757_ ) );
XNOR2_X1 _13519_ ( .A(_03908_ ), .B(\ID_EX_pc [4] ), .ZN(_05758_ ) );
OAI21_X1 _13520_ ( .A(_05210_ ), .B1(_05450_ ), .B2(_05758_ ), .ZN(_05759_ ) );
OAI221_X1 _13521_ ( .A(_05506_ ), .B1(_05436_ ), .B2(_05754_ ), .C1(_05757_ ), .C2(_05759_ ), .ZN(_05760_ ) );
XNOR2_X1 _13522_ ( .A(_02771_ ), .B(_02867_ ), .ZN(_05761_ ) );
AOI22_X1 _13523_ ( .A1(_05761_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05756_ ), .ZN(_05762_ ) );
AOI21_X1 _13524_ ( .A(_05743_ ), .B1(_05760_ ), .B2(_05762_ ), .ZN(_00141_ ) );
NAND3_X1 _13525_ ( .A1(_05507_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_05246_ ), .ZN(_05763_ ) );
NAND4_X1 _13526_ ( .A1(_05417_ ), .A2(_05235_ ), .A3(_05261_ ), .A4(\mepc [3] ), .ZN(_05764_ ) );
NAND3_X1 _13527_ ( .A1(_05763_ ), .A2(_05256_ ), .A3(_05764_ ), .ZN(_05765_ ) );
AND4_X1 _13528_ ( .A1(\mtvec [3] ), .A2(_05264_ ), .A3(_05261_ ), .A4(_05268_ ), .ZN(_05766_ ) );
NOR2_X1 _13529_ ( .A1(_05765_ ), .A2(_05766_ ), .ZN(_05767_ ) );
NAND3_X1 _13530_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_05444_ ), .ZN(_05768_ ) );
NAND3_X1 _13531_ ( .A1(_05745_ ), .A2(_05767_ ), .A3(_05768_ ), .ZN(_05769_ ) );
OR3_X1 _13532_ ( .A1(_05534_ ), .A2(\EX_LS_result_csreg_mem [3] ), .A3(_05535_ ), .ZN(_05770_ ) );
AND2_X1 _13533_ ( .A1(_05769_ ), .A2(_05770_ ), .ZN(_05771_ ) );
XOR2_X1 _13534_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .Z(_05772_ ) );
NOR2_X1 _13535_ ( .A1(_03953_ ), .A2(_03951_ ), .ZN(_05773_ ) );
XNOR2_X1 _13536_ ( .A(_03950_ ), .B(_05773_ ), .ZN(_05774_ ) );
MUX2_X1 _13537_ ( .A(_05772_ ), .B(_05774_ ), .S(_05202_ ), .Z(_05775_ ) );
MUX2_X1 _13538_ ( .A(_05771_ ), .B(_05775_ ), .S(_05210_ ), .Z(_05776_ ) );
NAND2_X1 _13539_ ( .A1(_05776_ ), .A2(_05345_ ), .ZN(_05777_ ) );
XOR2_X1 _13540_ ( .A(_02745_ ), .B(_02767_ ), .Z(_05778_ ) );
AOI22_X1 _13541_ ( .A1(_05778_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05774_ ), .ZN(_05779_ ) );
AOI21_X1 _13542_ ( .A(_05743_ ), .B1(_05777_ ), .B2(_05779_ ), .ZN(_00142_ ) );
AOI211_X1 _13543_ ( .A(_03946_ ), .B(_03942_ ), .C1(_03944_ ), .C2(_03943_ ), .ZN(_05780_ ) );
NOR2_X1 _13544_ ( .A1(_03948_ ), .A2(_05780_ ), .ZN(_05781_ ) );
MUX2_X1 _13545_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B(_05781_ ), .S(_05203_ ), .Z(_05782_ ) );
AND2_X1 _13546_ ( .A1(_05782_ ), .A2(_05210_ ), .ZN(_05783_ ) );
NAND3_X1 _13547_ ( .A1(_05239_ ), .A2(\mycsreg.CSReg[3][2] ), .A3(_05245_ ), .ZN(_05784_ ) );
NAND4_X1 _13548_ ( .A1(_05250_ ), .A2(_05235_ ), .A3(_05238_ ), .A4(\mepc [2] ), .ZN(_05785_ ) );
AND3_X1 _13549_ ( .A1(_05784_ ), .A2(_05363_ ), .A3(_05785_ ), .ZN(_05786_ ) );
NAND4_X1 _13550_ ( .A1(_05263_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mtvec [2] ), .ZN(_05787_ ) );
NAND3_X1 _13551_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_05327_ ), .ZN(_05788_ ) );
NAND3_X1 _13552_ ( .A1(_05786_ ), .A2(_05787_ ), .A3(_05788_ ), .ZN(_05789_ ) );
OAI21_X1 _13553_ ( .A(_05789_ ), .B1(_05232_ ), .B2(_05230_ ), .ZN(_05790_ ) );
NAND4_X1 _13554_ ( .A1(_05224_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_02128_ ), .A4(_05229_ ), .ZN(_05791_ ) );
AOI21_X1 _13555_ ( .A(_05283_ ), .B1(_05790_ ), .B2(_05791_ ), .ZN(_05792_ ) );
OAI21_X1 _13556_ ( .A(_05345_ ), .B1(_05783_ ), .B2(_05792_ ), .ZN(_05793_ ) );
XOR2_X1 _13557_ ( .A(_02743_ ), .B(_02744_ ), .Z(_05794_ ) );
AOI22_X1 _13558_ ( .A1(_05794_ ), .A2(_05577_ ), .B1(_05578_ ), .B2(_05781_ ), .ZN(_05795_ ) );
AOI21_X1 _13559_ ( .A(_05743_ ), .B1(_05793_ ), .B2(_05795_ ), .ZN(_00143_ ) );
NOR2_X1 _13560_ ( .A1(_05373_ ), .A2(\ID_EX_pc [1] ), .ZN(_05796_ ) );
XOR2_X1 _13561_ ( .A(_03943_ ), .B(_03944_ ), .Z(_05797_ ) );
INV_X1 _13562_ ( .A(_05797_ ), .ZN(_05798_ ) );
AOI211_X1 _13563_ ( .A(\ID_EX_typ [3] ), .B(_05796_ ), .C1(_05377_ ), .C2(_05798_ ), .ZN(_05799_ ) );
NAND3_X1 _13564_ ( .A1(_05240_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_05322_ ), .ZN(_05800_ ) );
NAND3_X1 _13565_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_05475_ ), .ZN(_05801_ ) );
NAND4_X1 _13566_ ( .A1(_05389_ ), .A2(_05259_ ), .A3(_05475_ ), .A4(\mepc [1] ), .ZN(_05802_ ) );
NAND4_X1 _13567_ ( .A1(_05392_ ), .A2(_05475_ ), .A3(_05394_ ), .A4(\mtvec [1] ), .ZN(_05803_ ) );
NAND4_X1 _13568_ ( .A1(_05800_ ), .A2(_05801_ ), .A3(_05802_ ), .A4(_05803_ ), .ZN(_05804_ ) );
OAI21_X1 _13569_ ( .A(_05804_ ), .B1(_05231_ ), .B2(_05387_ ), .ZN(_05805_ ) );
NAND4_X1 _13570_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_03841_ ), .A4(_05401_ ), .ZN(_05806_ ) );
AOI21_X1 _13571_ ( .A(_05454_ ), .B1(_05805_ ), .B2(_05806_ ), .ZN(_05807_ ) );
OAI21_X1 _13572_ ( .A(_05345_ ), .B1(_05799_ ), .B2(_05807_ ), .ZN(_05808_ ) );
XOR2_X1 _13573_ ( .A(_02719_ ), .B(_02741_ ), .Z(_05809_ ) );
AOI22_X1 _13574_ ( .A1(_05809_ ), .A2(_05371_ ), .B1(_03887_ ), .B2(_05797_ ), .ZN(_05810_ ) );
AOI21_X1 _13575_ ( .A(_05743_ ), .B1(_05808_ ), .B2(_05810_ ), .ZN(_00144_ ) );
NAND3_X1 _13576_ ( .A1(_05286_ ), .A2(\ID_EX_pc [26] ), .A3(_05289_ ), .ZN(_05811_ ) );
XNOR2_X1 _13577_ ( .A(_05811_ ), .B(\ID_EX_pc [27] ), .ZN(_05812_ ) );
OAI21_X1 _13578_ ( .A(_05812_ ), .B1(_05198_ ), .B2(_05201_ ), .ZN(_05813_ ) );
OR2_X1 _13579_ ( .A1(_04029_ ), .A2(_04030_ ), .ZN(_05814_ ) );
AND2_X1 _13580_ ( .A1(_05814_ ), .A2(_03928_ ), .ZN(_05815_ ) );
OR2_X1 _13581_ ( .A1(_05815_ ), .A2(_04032_ ), .ZN(_05816_ ) );
XNOR2_X1 _13582_ ( .A(_05816_ ), .B(_03927_ ), .ZN(_05817_ ) );
OAI211_X1 _13583_ ( .A(_05283_ ), .B(_05813_ ), .C1(_05297_ ), .C2(_05817_ ), .ZN(_05818_ ) );
NAND3_X1 _13584_ ( .A1(_05241_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_05246_ ), .ZN(_05819_ ) );
NAND3_X1 _13585_ ( .A1(_05507_ ), .A2(\mepc [27] ), .A3(_05258_ ), .ZN(_05820_ ) );
NAND4_X1 _13586_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [27] ), .A4(_05444_ ), .ZN(_05821_ ) );
NAND4_X1 _13587_ ( .A1(_05542_ ), .A2(_05819_ ), .A3(_05820_ ), .A4(_05821_ ), .ZN(_05822_ ) );
AND3_X1 _13588_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_05444_ ), .ZN(_05823_ ) );
NOR3_X1 _13589_ ( .A1(_05822_ ), .A2(_05744_ ), .A3(_05823_ ), .ZN(_05824_ ) );
NOR3_X1 _13590_ ( .A1(_05547_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_05536_ ), .ZN(_05825_ ) );
NOR2_X1 _13591_ ( .A1(_05824_ ), .A2(_05825_ ), .ZN(_05826_ ) );
OAI211_X1 _13592_ ( .A(_05818_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05826_ ), .ZN(_05827_ ) );
MUX2_X1 _13593_ ( .A(_03051_ ), .B(_05817_ ), .S(_05405_ ), .Z(_05828_ ) );
OR2_X1 _13594_ ( .A1(_05828_ ), .A2(_05343_ ), .ZN(_05829_ ) );
AOI21_X1 _13595_ ( .A(_05743_ ), .B1(_05827_ ), .B2(_05829_ ), .ZN(_00145_ ) );
XOR2_X1 _13596_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05830_ ) );
MUX2_X1 _13597_ ( .A(\ID_EX_pc [0] ), .B(_05830_ ), .S(_05203_ ), .Z(_05831_ ) );
AND2_X1 _13598_ ( .A1(_05831_ ), .A2(_05210_ ), .ZN(_05832_ ) );
OR3_X1 _13599_ ( .A1(_05547_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_05536_ ), .ZN(_05833_ ) );
AND2_X1 _13600_ ( .A1(_05540_ ), .A2(_05323_ ), .ZN(_05834_ ) );
INV_X1 _13601_ ( .A(_05834_ ), .ZN(_05835_ ) );
NAND3_X1 _13602_ ( .A1(_05321_ ), .A2(\mepc [0] ), .A3(_05389_ ), .ZN(_05836_ ) );
NAND3_X1 _13603_ ( .A1(_05321_ ), .A2(\mycsreg.CSReg[3][0] ), .A3(_05323_ ), .ZN(_05837_ ) );
NAND3_X1 _13604_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_05390_ ), .ZN(_05838_ ) );
NAND4_X1 _13605_ ( .A1(_05835_ ), .A2(_05836_ ), .A3(_05837_ ), .A4(_05838_ ), .ZN(_05839_ ) );
NAND4_X1 _13606_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [0] ), .A4(_05390_ ), .ZN(_05840_ ) );
OAI21_X1 _13607_ ( .A(_05840_ ), .B1(_05547_ ), .B2(_05536_ ), .ZN(_05841_ ) );
OAI211_X1 _13608_ ( .A(_05833_ ), .B(\ID_EX_typ [3] ), .C1(_05839_ ), .C2(_05841_ ), .ZN(_05842_ ) );
INV_X1 _13609_ ( .A(_05842_ ), .ZN(_05843_ ) );
OAI21_X1 _13610_ ( .A(_05345_ ), .B1(_05832_ ), .B2(_05843_ ), .ZN(_05844_ ) );
NAND4_X1 _13611_ ( .A1(_05830_ ), .A2(\ID_EX_typ [5] ), .A3(_05623_ ), .A4(_03884_ ), .ZN(_05845_ ) );
AOI21_X1 _13612_ ( .A(_05743_ ), .B1(_05844_ ), .B2(_05845_ ), .ZN(_00146_ ) );
XNOR2_X1 _13613_ ( .A(_05290_ ), .B(_05292_ ), .ZN(_05846_ ) );
AND2_X1 _13614_ ( .A1(_05297_ ), .A2(_05846_ ), .ZN(_05847_ ) );
XOR2_X1 _13615_ ( .A(_05814_ ), .B(_03928_ ), .Z(_05848_ ) );
INV_X1 _13616_ ( .A(_05848_ ), .ZN(_05849_ ) );
AOI211_X1 _13617_ ( .A(\ID_EX_typ [3] ), .B(_05847_ ), .C1(_05377_ ), .C2(_05849_ ), .ZN(_05850_ ) );
NAND3_X1 _13618_ ( .A1(_05240_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_05322_ ), .ZN(_05851_ ) );
NAND3_X1 _13619_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_05475_ ), .ZN(_05852_ ) );
NAND4_X1 _13620_ ( .A1(_05389_ ), .A2(_05259_ ), .A3(_05475_ ), .A4(\mepc [26] ), .ZN(_05853_ ) );
NAND4_X1 _13621_ ( .A1(_05392_ ), .A2(_05475_ ), .A3(_05394_ ), .A4(\mtvec [26] ), .ZN(_05854_ ) );
NAND4_X1 _13622_ ( .A1(_05851_ ), .A2(_05852_ ), .A3(_05853_ ), .A4(_05854_ ), .ZN(_05855_ ) );
OAI21_X1 _13623_ ( .A(_05855_ ), .B1(_05231_ ), .B2(_05387_ ), .ZN(_05856_ ) );
NAND4_X1 _13624_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_03841_ ), .A4(_05401_ ), .ZN(_05857_ ) );
AOI21_X1 _13625_ ( .A(_05454_ ), .B1(_05856_ ), .B2(_05857_ ), .ZN(_05858_ ) );
OAI21_X1 _13626_ ( .A(_05208_ ), .B1(_05850_ ), .B2(_05858_ ), .ZN(_05859_ ) );
OAI21_X1 _13627_ ( .A(fanout_net_4 ), .B1(_03049_ ), .B2(_03052_ ), .ZN(_05860_ ) );
OAI211_X1 _13628_ ( .A(_05280_ ), .B(_05860_ ), .C1(_05848_ ), .C2(fanout_net_4 ), .ZN(_05861_ ) );
AOI21_X1 _13629_ ( .A(_05743_ ), .B1(_05859_ ), .B2(_05861_ ), .ZN(_00147_ ) );
AND3_X1 _13630_ ( .A1(_05288_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05862_ ) );
AND2_X1 _13631_ ( .A1(_05286_ ), .A2(_05862_ ), .ZN(_05863_ ) );
NAND3_X1 _13632_ ( .A1(_05863_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05864_ ) );
INV_X1 _13633_ ( .A(\ID_EX_pc [24] ), .ZN(_05865_ ) );
NOR2_X1 _13634_ ( .A1(_05864_ ), .A2(_05865_ ), .ZN(_05866_ ) );
XNOR2_X1 _13635_ ( .A(_05866_ ), .B(_04028_ ), .ZN(_05867_ ) );
NOR2_X1 _13636_ ( .A1(_05373_ ), .A2(_05867_ ), .ZN(_05868_ ) );
NAND2_X1 _13637_ ( .A1(_04026_ ), .A2(_04027_ ), .ZN(_05869_ ) );
XOR2_X1 _13638_ ( .A(\ID_EX_pc [25] ), .B(\ID_EX_imm [25] ), .Z(_05870_ ) );
XNOR2_X1 _13639_ ( .A(_05869_ ), .B(_05870_ ), .ZN(_05871_ ) );
AOI211_X1 _13640_ ( .A(\ID_EX_typ [3] ), .B(_05868_ ), .C1(_05377_ ), .C2(_05871_ ), .ZN(_05872_ ) );
NAND3_X1 _13641_ ( .A1(_05507_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_05246_ ), .ZN(_05873_ ) );
NAND3_X1 _13642_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_05265_ ), .ZN(_05874_ ) );
NAND4_X1 _13643_ ( .A1(_05389_ ), .A2(_05259_ ), .A3(_05475_ ), .A4(\mepc [25] ), .ZN(_05875_ ) );
NAND4_X1 _13644_ ( .A1(_05392_ ), .A2(_05475_ ), .A3(_05394_ ), .A4(\mtvec [25] ), .ZN(_05876_ ) );
NAND4_X1 _13645_ ( .A1(_05873_ ), .A2(_05874_ ), .A3(_05875_ ), .A4(_05876_ ), .ZN(_05877_ ) );
OAI21_X1 _13646_ ( .A(_05877_ ), .B1(_05231_ ), .B2(_05387_ ), .ZN(_05878_ ) );
BUF_X4 _13647_ ( .A(_03840_ ), .Z(_05879_ ) );
NAND4_X1 _13648_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_05879_ ), .A4(_05401_ ), .ZN(_05880_ ) );
AOI21_X1 _13649_ ( .A(_05454_ ), .B1(_05878_ ), .B2(_05880_ ), .ZN(_05881_ ) );
OAI21_X1 _13650_ ( .A(_05208_ ), .B1(_05872_ ), .B2(_05881_ ), .ZN(_05882_ ) );
NOR2_X1 _13651_ ( .A1(_05871_ ), .A2(_03888_ ), .ZN(_05883_ ) );
BUF_X2 _13652_ ( .A(_05405_ ), .Z(_05884_ ) );
NOR3_X1 _13653_ ( .A1(_03054_ ), .A2(_05884_ ), .A3(_05207_ ), .ZN(_05885_ ) );
NOR2_X1 _13654_ ( .A1(_05883_ ), .A2(_05885_ ), .ZN(_05886_ ) );
AOI21_X1 _13655_ ( .A(_05743_ ), .B1(_05882_ ), .B2(_05886_ ), .ZN(_00148_ ) );
XNOR2_X1 _13656_ ( .A(_05864_ ), .B(\ID_EX_pc [24] ), .ZN(_05887_ ) );
NOR2_X1 _13657_ ( .A1(_05373_ ), .A2(_05887_ ), .ZN(_05888_ ) );
XOR2_X1 _13658_ ( .A(_04024_ ), .B(_04025_ ), .Z(_05889_ ) );
INV_X1 _13659_ ( .A(_05889_ ), .ZN(_05890_ ) );
AOI211_X1 _13660_ ( .A(\ID_EX_typ [3] ), .B(_05888_ ), .C1(_05377_ ), .C2(_05890_ ), .ZN(_05891_ ) );
AND3_X1 _13661_ ( .A1(_05507_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_05246_ ), .ZN(_05892_ ) );
INV_X1 _13662_ ( .A(_05892_ ), .ZN(_05893_ ) );
NAND4_X1 _13663_ ( .A1(_05389_ ), .A2(_05259_ ), .A3(_05390_ ), .A4(\mepc [24] ), .ZN(_05894_ ) );
NAND4_X1 _13664_ ( .A1(_05392_ ), .A2(_05390_ ), .A3(_05394_ ), .A4(\mtvec [24] ), .ZN(_05895_ ) );
NAND4_X1 _13665_ ( .A1(_05364_ ), .A2(_05893_ ), .A3(_05894_ ), .A4(_05895_ ), .ZN(_05896_ ) );
AND3_X1 _13666_ ( .A1(_05397_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_05475_ ), .ZN(_05897_ ) );
OAI22_X1 _13667_ ( .A1(_05896_ ), .A2(_05897_ ), .B1(_05387_ ), .B2(_05231_ ), .ZN(_05898_ ) );
NAND4_X1 _13668_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_05879_ ), .A4(_05401_ ), .ZN(_05899_ ) );
AOI21_X1 _13669_ ( .A(_05454_ ), .B1(_05898_ ), .B2(_05899_ ), .ZN(_05900_ ) );
OAI21_X1 _13670_ ( .A(_05208_ ), .B1(_05891_ ), .B2(_05900_ ), .ZN(_05901_ ) );
NOR4_X1 _13671_ ( .A1(_03055_ ), .A2(_02915_ ), .A3(_05433_ ), .A4(_05206_ ), .ZN(_05902_ ) );
AOI21_X1 _13672_ ( .A(_05902_ ), .B1(_05889_ ), .B2(_05370_ ), .ZN(_05903_ ) );
AOI21_X1 _13673_ ( .A(_05743_ ), .B1(_05901_ ), .B2(_05903_ ), .ZN(_00149_ ) );
NAND3_X1 _13674_ ( .A1(_05286_ ), .A2(\ID_EX_pc [22] ), .A3(_05862_ ), .ZN(_05904_ ) );
XNOR2_X1 _13675_ ( .A(_05904_ ), .B(\ID_EX_pc [23] ), .ZN(_05905_ ) );
OAI21_X1 _13676_ ( .A(_05905_ ), .B1(_05198_ ), .B2(_05201_ ), .ZN(_05906_ ) );
NAND2_X1 _13677_ ( .A1(_05347_ ), .A2(_03934_ ), .ZN(_05907_ ) );
NAND2_X1 _13678_ ( .A1(_05907_ ), .A2(_04021_ ), .ZN(_05908_ ) );
NAND2_X1 _13679_ ( .A1(_05908_ ), .A2(_03930_ ), .ZN(_05909_ ) );
NAND2_X1 _13680_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_05910_ ) );
NAND2_X1 _13681_ ( .A1(_05909_ ), .A2(_05910_ ), .ZN(_05911_ ) );
XNOR2_X1 _13682_ ( .A(_05911_ ), .B(_03929_ ), .ZN(_05912_ ) );
OAI211_X1 _13683_ ( .A(_05283_ ), .B(_05906_ ), .C1(_05297_ ), .C2(_05912_ ), .ZN(_05913_ ) );
NAND3_X1 _13684_ ( .A1(_05321_ ), .A2(\mepc [23] ), .A3(_05258_ ), .ZN(_05914_ ) );
NAND4_X1 _13685_ ( .A1(_05331_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mycsreg.CSReg[0][23] ), .ZN(_05915_ ) );
AND2_X1 _13686_ ( .A1(_05914_ ), .A2(_05915_ ), .ZN(_05916_ ) );
NAND3_X1 _13687_ ( .A1(_05321_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_05323_ ), .ZN(_05917_ ) );
NAND4_X1 _13688_ ( .A1(_05326_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mtvec [23] ), .ZN(_05918_ ) );
AND2_X1 _13689_ ( .A1(_05917_ ), .A2(_05918_ ), .ZN(_05919_ ) );
OAI211_X1 _13690_ ( .A(_05916_ ), .B(_05919_ ), .C1(_05547_ ), .C2(_05536_ ), .ZN(_05920_ ) );
OR3_X1 _13691_ ( .A1(_05547_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_05536_ ), .ZN(_05921_ ) );
NAND2_X1 _13692_ ( .A1(_05920_ ), .A2(_05921_ ), .ZN(_05922_ ) );
INV_X1 _13693_ ( .A(_05922_ ), .ZN(_05923_ ) );
OAI211_X1 _13694_ ( .A(_05913_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05923_ ), .ZN(_05924_ ) );
MUX2_X1 _13695_ ( .A(_05912_ ), .B(_03060_ ), .S(fanout_net_4 ), .Z(_05925_ ) );
OR2_X1 _13696_ ( .A1(_05925_ ), .A2(_05343_ ), .ZN(_05926_ ) );
AOI21_X1 _13697_ ( .A(_05743_ ), .B1(_05924_ ), .B2(_05926_ ), .ZN(_00150_ ) );
XNOR2_X1 _13698_ ( .A(_05863_ ), .B(\ID_EX_pc [22] ), .ZN(_05927_ ) );
XOR2_X1 _13699_ ( .A(_05908_ ), .B(_03930_ ), .Z(_05928_ ) );
INV_X1 _13700_ ( .A(_05928_ ), .ZN(_05929_ ) );
MUX2_X1 _13701_ ( .A(_05927_ ), .B(_05929_ ), .S(_05203_ ), .Z(_05930_ ) );
NAND2_X1 _13702_ ( .A1(_05930_ ), .A2(_05436_ ), .ZN(_05931_ ) );
AND3_X1 _13703_ ( .A1(_05320_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_05322_ ), .ZN(_05932_ ) );
AND4_X1 _13704_ ( .A1(\mtvec [22] ), .A2(_05263_ ), .A3(_05356_ ), .A4(_05357_ ), .ZN(_05933_ ) );
NOR2_X1 _13705_ ( .A1(_05932_ ), .A2(_05933_ ), .ZN(_05934_ ) );
NAND3_X1 _13706_ ( .A1(_05241_ ), .A2(\mepc [22] ), .A3(_05258_ ), .ZN(_05935_ ) );
NAND4_X1 _13707_ ( .A1(_05331_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mycsreg.CSReg[0][22] ), .ZN(_05936_ ) );
NAND4_X1 _13708_ ( .A1(_05934_ ), .A2(_05513_ ), .A3(_05935_ ), .A4(_05936_ ), .ZN(_05937_ ) );
NAND2_X1 _13709_ ( .A1(_05314_ ), .A2(_05937_ ), .ZN(_05938_ ) );
NAND3_X1 _13710_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_05428_ ), .ZN(_05939_ ) );
NAND2_X1 _13711_ ( .A1(_05938_ ), .A2(_05939_ ), .ZN(_05940_ ) );
OAI211_X1 _13712_ ( .A(_05931_ ), .B(_05416_ ), .C1(_05211_ ), .C2(_05940_ ), .ZN(_05941_ ) );
AOI22_X1 _13713_ ( .A1(_03061_ ), .A2(_05371_ ), .B1(_03887_ ), .B2(_05928_ ), .ZN(_05942_ ) );
AOI21_X1 _13714_ ( .A(_03906_ ), .B1(_05941_ ), .B2(_05942_ ), .ZN(_00151_ ) );
INV_X1 _13715_ ( .A(\ID_EX_pc [20] ), .ZN(_05943_ ) );
NOR2_X1 _13716_ ( .A1(_05350_ ), .A2(_05943_ ), .ZN(_05944_ ) );
INV_X1 _13717_ ( .A(\ID_EX_pc [21] ), .ZN(_05945_ ) );
XNOR2_X1 _13718_ ( .A(_05944_ ), .B(_05945_ ), .ZN(_05946_ ) );
NOR2_X1 _13719_ ( .A1(_05203_ ), .A2(_05946_ ), .ZN(_05947_ ) );
AND2_X1 _13720_ ( .A1(_05347_ ), .A2(_03932_ ), .ZN(_05948_ ) );
OR2_X1 _13721_ ( .A1(_05948_ ), .A2(_04020_ ), .ZN(_05949_ ) );
XNOR2_X1 _13722_ ( .A(_05949_ ), .B(_03933_ ), .ZN(_05950_ ) );
AOI211_X1 _13723_ ( .A(\ID_EX_typ [3] ), .B(_05947_ ), .C1(_05377_ ), .C2(_05950_ ), .ZN(_05951_ ) );
NAND4_X1 _13724_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [21] ), .A4(_05327_ ), .ZN(_05952_ ) );
NAND3_X1 _13725_ ( .A1(_05354_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_05322_ ), .ZN(_05953_ ) );
AND3_X1 _13726_ ( .A1(_05952_ ), .A2(_05256_ ), .A3(_05953_ ), .ZN(_05954_ ) );
NAND3_X1 _13727_ ( .A1(_05507_ ), .A2(\mepc [21] ), .A3(_05417_ ), .ZN(_05955_ ) );
NAND3_X1 _13728_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_05261_ ), .ZN(_05956_ ) );
AND2_X1 _13729_ ( .A1(_05955_ ), .A2(_05956_ ), .ZN(_05957_ ) );
NAND3_X1 _13730_ ( .A1(_05745_ ), .A2(_05954_ ), .A3(_05957_ ), .ZN(_05958_ ) );
NOR3_X1 _13731_ ( .A1(_05534_ ), .A2(\EX_LS_result_csreg_mem [21] ), .A3(_05535_ ), .ZN(_05959_ ) );
INV_X1 _13732_ ( .A(_05959_ ), .ZN(_05960_ ) );
AND3_X1 _13733_ ( .A1(_05958_ ), .A2(\ID_EX_typ [3] ), .A3(_05960_ ), .ZN(_05961_ ) );
OAI21_X1 _13734_ ( .A(_05208_ ), .B1(_05951_ ), .B2(_05961_ ), .ZN(_05962_ ) );
NOR3_X1 _13735_ ( .A1(_03016_ ), .A2(_05884_ ), .A3(_05207_ ), .ZN(_05963_ ) );
NOR2_X1 _13736_ ( .A1(_05950_ ), .A2(_03888_ ), .ZN(_05964_ ) );
NOR2_X1 _13737_ ( .A1(_05963_ ), .A2(_05964_ ), .ZN(_05965_ ) );
AOI21_X1 _13738_ ( .A(_03906_ ), .B1(_05962_ ), .B2(_05965_ ), .ZN(_00152_ ) );
INV_X1 _13739_ ( .A(\ID_EX_pc [30] ), .ZN(_05966_ ) );
NOR2_X1 _13740_ ( .A1(_03925_ ), .A2(_05966_ ), .ZN(_05967_ ) );
XNOR2_X1 _13741_ ( .A(_05967_ ), .B(\ID_EX_pc [31] ), .ZN(_05968_ ) );
AND2_X1 _13742_ ( .A1(_05297_ ), .A2(_05968_ ), .ZN(_05969_ ) );
OAI21_X1 _13743_ ( .A(_04043_ ), .B1(_04040_ ), .B2(_04041_ ), .ZN(_05970_ ) );
NAND2_X1 _13744_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_05971_ ) );
AND2_X1 _13745_ ( .A1(_05970_ ), .A2(_05971_ ), .ZN(_05972_ ) );
XNOR2_X1 _13746_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_05973_ ) );
XNOR2_X1 _13747_ ( .A(_05972_ ), .B(_05973_ ), .ZN(_05974_ ) );
AOI211_X1 _13748_ ( .A(\ID_EX_typ [3] ), .B(_05969_ ), .C1(_05450_ ), .C2(_05974_ ), .ZN(_05975_ ) );
AND3_X1 _13749_ ( .A1(_05273_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_05260_ ), .ZN(_05976_ ) );
NAND3_X1 _13750_ ( .A1(_05240_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_05245_ ), .ZN(_05977_ ) );
NAND4_X1 _13751_ ( .A1(_05250_ ), .A2(_05235_ ), .A3(_05260_ ), .A4(\mepc [31] ), .ZN(_05978_ ) );
NAND4_X1 _13752_ ( .A1(_05263_ ), .A2(_05260_ ), .A3(_05267_ ), .A4(\mtvec [31] ), .ZN(_05979_ ) );
NAND3_X1 _13753_ ( .A1(_05977_ ), .A2(_05978_ ), .A3(_05979_ ), .ZN(_05980_ ) );
NOR3_X1 _13754_ ( .A1(_05744_ ), .A2(_05976_ ), .A3(_05980_ ), .ZN(_05981_ ) );
NOR3_X1 _13755_ ( .A1(_05534_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_05535_ ), .ZN(_05982_ ) );
NOR3_X1 _13756_ ( .A1(_05981_ ), .A2(_05210_ ), .A3(_05982_ ), .ZN(_05983_ ) );
OAI21_X1 _13757_ ( .A(_05416_ ), .B1(_05975_ ), .B2(_05983_ ), .ZN(_05984_ ) );
MUX2_X1 _13758_ ( .A(_03007_ ), .B(_05974_ ), .S(_05433_ ), .Z(_05985_ ) );
OAI211_X1 _13759_ ( .A(_05984_ ), .B(_03897_ ), .C1(_05345_ ), .C2(_05985_ ), .ZN(_00153_ ) );
AND3_X1 _13760_ ( .A1(_03903_ ), .A2(\ID_EX_pc [31] ), .A3(_03905_ ), .ZN(_00154_ ) );
AND3_X1 _13761_ ( .A1(_03903_ ), .A2(\ID_EX_pc [30] ), .A3(_03905_ ), .ZN(_00155_ ) );
AND3_X1 _13762_ ( .A1(_03903_ ), .A2(\ID_EX_pc [21] ), .A3(_03905_ ), .ZN(_00156_ ) );
AND3_X1 _13763_ ( .A1(_03903_ ), .A2(\ID_EX_pc [20] ), .A3(_03905_ ), .ZN(_00157_ ) );
AND3_X1 _13764_ ( .A1(_03903_ ), .A2(\ID_EX_pc [19] ), .A3(_03905_ ), .ZN(_00158_ ) );
CLKBUF_X2 _13765_ ( .A(_03894_ ), .Z(_05986_ ) );
CLKBUF_X2 _13766_ ( .A(_03895_ ), .Z(_05987_ ) );
AND3_X1 _13767_ ( .A1(_05986_ ), .A2(\ID_EX_pc [18] ), .A3(_05987_ ), .ZN(_00159_ ) );
AND3_X1 _13768_ ( .A1(_05986_ ), .A2(\ID_EX_pc [17] ), .A3(_05987_ ), .ZN(_00160_ ) );
AND3_X1 _13769_ ( .A1(_05986_ ), .A2(\ID_EX_pc [16] ), .A3(_05987_ ), .ZN(_00161_ ) );
AND3_X1 _13770_ ( .A1(_05986_ ), .A2(\ID_EX_pc [15] ), .A3(_05987_ ), .ZN(_00162_ ) );
AND3_X1 _13771_ ( .A1(_05986_ ), .A2(\ID_EX_pc [14] ), .A3(_05987_ ), .ZN(_00163_ ) );
AND3_X1 _13772_ ( .A1(_05986_ ), .A2(\ID_EX_pc [13] ), .A3(_05987_ ), .ZN(_00164_ ) );
AND3_X1 _13773_ ( .A1(_05986_ ), .A2(\ID_EX_pc [12] ), .A3(_05987_ ), .ZN(_00165_ ) );
AND3_X1 _13774_ ( .A1(_05986_ ), .A2(\ID_EX_pc [29] ), .A3(_05987_ ), .ZN(_00166_ ) );
AND3_X1 _13775_ ( .A1(_05986_ ), .A2(\ID_EX_pc [11] ), .A3(_05987_ ), .ZN(_00167_ ) );
AND3_X1 _13776_ ( .A1(_05986_ ), .A2(\ID_EX_pc [10] ), .A3(_05987_ ), .ZN(_00168_ ) );
CLKBUF_X2 _13777_ ( .A(_03894_ ), .Z(_05988_ ) );
CLKBUF_X2 _13778_ ( .A(_03895_ ), .Z(_05989_ ) );
AND3_X1 _13779_ ( .A1(_05988_ ), .A2(\ID_EX_pc [9] ), .A3(_05989_ ), .ZN(_00169_ ) );
AND3_X1 _13780_ ( .A1(_05988_ ), .A2(\ID_EX_pc [8] ), .A3(_05989_ ), .ZN(_00170_ ) );
AND3_X1 _13781_ ( .A1(_05988_ ), .A2(\ID_EX_pc [7] ), .A3(_05989_ ), .ZN(_00171_ ) );
AND3_X1 _13782_ ( .A1(_05988_ ), .A2(\ID_EX_pc [6] ), .A3(_05989_ ), .ZN(_00172_ ) );
AND3_X1 _13783_ ( .A1(_05988_ ), .A2(\ID_EX_pc [5] ), .A3(_05989_ ), .ZN(_00173_ ) );
AND3_X1 _13784_ ( .A1(_05988_ ), .A2(\ID_EX_pc [4] ), .A3(_05989_ ), .ZN(_00174_ ) );
AND3_X1 _13785_ ( .A1(_05988_ ), .A2(\ID_EX_pc [3] ), .A3(_05989_ ), .ZN(_00175_ ) );
AND3_X1 _13786_ ( .A1(_05988_ ), .A2(\ID_EX_pc [2] ), .A3(_05989_ ), .ZN(_00176_ ) );
AND3_X1 _13787_ ( .A1(_05988_ ), .A2(\ID_EX_pc [28] ), .A3(_05989_ ), .ZN(_00177_ ) );
AND3_X1 _13788_ ( .A1(_05988_ ), .A2(\ID_EX_pc [1] ), .A3(_05989_ ), .ZN(_00178_ ) );
CLKBUF_X2 _13789_ ( .A(_03894_ ), .Z(_05990_ ) );
CLKBUF_X2 _13790_ ( .A(_03895_ ), .Z(_05991_ ) );
AND3_X1 _13791_ ( .A1(_05990_ ), .A2(\ID_EX_pc [0] ), .A3(_05991_ ), .ZN(_00179_ ) );
AND3_X1 _13792_ ( .A1(_05990_ ), .A2(\ID_EX_pc [27] ), .A3(_05991_ ), .ZN(_00180_ ) );
AND3_X1 _13793_ ( .A1(_05990_ ), .A2(\ID_EX_pc [26] ), .A3(_05991_ ), .ZN(_00181_ ) );
AND3_X1 _13794_ ( .A1(_05990_ ), .A2(\ID_EX_pc [25] ), .A3(_05991_ ), .ZN(_00182_ ) );
AND3_X1 _13795_ ( .A1(_05990_ ), .A2(\ID_EX_pc [24] ), .A3(_05991_ ), .ZN(_00183_ ) );
AND3_X1 _13796_ ( .A1(_05990_ ), .A2(\ID_EX_pc [23] ), .A3(_05991_ ), .ZN(_00184_ ) );
AND3_X1 _13797_ ( .A1(_05990_ ), .A2(\ID_EX_pc [22] ), .A3(_05991_ ), .ZN(_00185_ ) );
AND3_X1 _13798_ ( .A1(_05990_ ), .A2(\ID_EX_typ [7] ), .A3(_05991_ ), .ZN(_00186_ ) );
MUX2_X1 _13799_ ( .A(io_master_arready ), .B(_01987_ ), .S(_02072_ ), .Z(_05992_ ) );
CLKBUF_X2 _13800_ ( .A(_01975_ ), .Z(\io_master_arid [1] ) );
AND2_X1 _13801_ ( .A1(_05992_ ), .A2(\io_master_arid [1] ), .ZN(_05993_ ) );
OR2_X1 _13802_ ( .A1(_05993_ ), .A2(_02040_ ), .ZN(_05994_ ) );
INV_X1 _13803_ ( .A(\mylsu.state [4] ), .ZN(_05995_ ) );
INV_X1 _13804_ ( .A(\mylsu.state [0] ), .ZN(_05996_ ) );
NAND2_X1 _13805_ ( .A1(_05995_ ), .A2(_05996_ ), .ZN(_05997_ ) );
INV_X1 _13806_ ( .A(io_master_awready ), .ZN(_05998_ ) );
NAND3_X1 _13807_ ( .A1(_02050_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A3(_05998_ ), .ZN(_05999_ ) );
AND3_X1 _13808_ ( .A1(_05994_ ), .A2(_05997_ ), .A3(_05999_ ), .ZN(_06000_ ) );
AND2_X1 _13809_ ( .A1(_03896_ ), .A2(EXU_valid_LSU ), .ZN(_06001_ ) );
INV_X1 _13810_ ( .A(_06001_ ), .ZN(_06002_ ) );
OAI22_X1 _13811_ ( .A1(_06000_ ), .A2(_06002_ ), .B1(_03883_ ), .B2(_03906_ ), .ZN(_00187_ ) );
AND3_X1 _13812_ ( .A1(_05990_ ), .A2(\ID_EX_typ [6] ), .A3(_05991_ ), .ZN(_00188_ ) );
AND3_X1 _13813_ ( .A1(_05990_ ), .A2(\ID_EX_typ [5] ), .A3(_05991_ ), .ZN(_00189_ ) );
AND3_X1 _13814_ ( .A1(_03902_ ), .A2(\ID_EX_typ [4] ), .A3(_03904_ ), .ZN(_00190_ ) );
AND3_X1 _13815_ ( .A1(_03902_ ), .A2(\ID_EX_typ [3] ), .A3(_03904_ ), .ZN(_00191_ ) );
AND3_X1 _13816_ ( .A1(_03902_ ), .A2(\ID_EX_typ [2] ), .A3(_03904_ ), .ZN(_00192_ ) );
AND3_X1 _13817_ ( .A1(_03902_ ), .A2(\ID_EX_typ [1] ), .A3(_03904_ ), .ZN(_00193_ ) );
AND3_X1 _13818_ ( .A1(_03902_ ), .A2(fanout_net_4 ), .A3(_03904_ ), .ZN(_00194_ ) );
AND2_X1 _13819_ ( .A1(_02062_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _13820_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .ZN(_06003_ ) );
BUF_X2 _13821_ ( .A(_06003_ ), .Z(_06004_ ) );
AND3_X1 _13822_ ( .A1(_02062_ ), .A2(_06004_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00242_ ) );
NAND2_X1 _13823_ ( .A1(_03748_ ), .A2(fanout_net_6 ), .ZN(_06005_ ) );
INV_X1 _13824_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_06006_ ) );
BUF_X4 _13825_ ( .A(_06006_ ), .Z(_06007_ ) );
NOR3_X1 _13826_ ( .A1(_02063_ ), .A2(_06005_ ), .A3(_06007_ ), .ZN(_00243_ ) );
NAND2_X1 _13827_ ( .A1(_03756_ ), .A2(fanout_net_10 ), .ZN(_06008_ ) );
NOR3_X1 _13828_ ( .A1(_02063_ ), .A2(_06008_ ), .A3(_06007_ ), .ZN(_00244_ ) );
AND3_X1 _13829_ ( .A1(_03902_ ), .A2(\EX_LS_pc [2] ), .A3(_03904_ ), .ZN(_00282_ ) );
AND2_X1 _13830_ ( .A1(_03897_ ), .A2(\mylsu.state [3] ), .ZN(_00283_ ) );
INV_X1 _13831_ ( .A(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06009_ ) );
AND2_X1 _13832_ ( .A1(_03896_ ), .A2(_06009_ ), .ZN(_06010_ ) );
NOR2_X1 _13833_ ( .A1(\mylsu.state [3] ), .A2(\mylsu.state [1] ), .ZN(_06011_ ) );
NAND2_X1 _13834_ ( .A1(_06010_ ), .A2(_06011_ ), .ZN(_06012_ ) );
OAI211_X1 _13835_ ( .A(_02049_ ), .B(_02089_ ), .C1(_02086_ ), .C2(_02087_ ), .ZN(_06013_ ) );
AND2_X1 _13836_ ( .A1(_06013_ ), .A2(\EX_LS_flag [2] ), .ZN(_06014_ ) );
NOR3_X1 _13837_ ( .A1(_02042_ ), .A2(_06014_ ), .A3(_02047_ ), .ZN(_06015_ ) );
AOI21_X1 _13838_ ( .A(_06012_ ), .B1(_03850_ ), .B2(_06015_ ), .ZN(_00296_ ) );
INV_X1 _13839_ ( .A(_03853_ ), .ZN(_06016_ ) );
AOI21_X1 _13840_ ( .A(_02083_ ), .B1(_06016_ ), .B2(_06014_ ), .ZN(_06017_ ) );
AOI21_X1 _13841_ ( .A(_06012_ ), .B1(_06017_ ), .B2(_03850_ ), .ZN(_00297_ ) );
NOR2_X1 _13842_ ( .A1(_02088_ ), .A2(_02090_ ), .ZN(_06018_ ) );
AND2_X1 _13843_ ( .A1(_02038_ ), .A2(\EX_LS_flag [2] ), .ZN(_06019_ ) );
AND4_X1 _13844_ ( .A1(_06018_ ), .A2(_06019_ ), .A3(_06011_ ), .A4(_06010_ ), .ZN(_00298_ ) );
AOI21_X1 _13845_ ( .A(_06012_ ), .B1(_03839_ ), .B2(_02048_ ), .ZN(_00299_ ) );
NAND2_X1 _13846_ ( .A1(_06018_ ), .A2(_06019_ ), .ZN(_06020_ ) );
AOI21_X1 _13847_ ( .A(_06012_ ), .B1(_03850_ ), .B2(_06020_ ), .ZN(_00300_ ) );
NAND2_X1 _13848_ ( .A1(_02037_ ), .A2(_02039_ ), .ZN(_06021_ ) );
NOR3_X1 _13849_ ( .A1(_02090_ ), .A2(_02050_ ), .A3(_01941_ ), .ZN(_06022_ ) );
OAI21_X1 _13850_ ( .A(_06022_ ), .B1(_02088_ ), .B2(\EX_LS_flag [1] ), .ZN(_06023_ ) );
AOI21_X1 _13851_ ( .A(_06023_ ), .B1(_05992_ ), .B2(\io_master_arid [1] ), .ZN(_06024_ ) );
OAI221_X1 _13852_ ( .A(_02039_ ), .B1(\EX_LS_typ [4] ), .B2(_06021_ ), .C1(_06024_ ), .C2(_02046_ ), .ZN(_06025_ ) );
INV_X1 _13853_ ( .A(_02052_ ), .ZN(_06026_ ) );
AND3_X1 _13854_ ( .A1(_06025_ ), .A2(_06026_ ), .A3(_06023_ ), .ZN(_06027_ ) );
NOR4_X1 _13855_ ( .A1(_06027_ ), .A2(_03899_ ), .A3(_02058_ ), .A4(_03846_ ), .ZN(_06028_ ) );
AND3_X1 _13856_ ( .A1(_06028_ ), .A2(_03897_ ), .A3(_06011_ ), .ZN(_00301_ ) );
INV_X1 _13857_ ( .A(_00283_ ), .ZN(_06029_ ) );
INV_X1 _13858_ ( .A(_02046_ ), .ZN(_06030_ ) );
OAI211_X1 _13859_ ( .A(EXU_valid_LSU ), .B(_06011_ ), .C1(_06030_ ), .C2(_03836_ ), .ZN(_06031_ ) );
NOR2_X1 _13860_ ( .A1(_03870_ ), .A2(\EX_LS_flag [1] ), .ZN(_06032_ ) );
OAI21_X1 _13861_ ( .A(_03897_ ), .B1(_03841_ ), .B2(_06032_ ), .ZN(_06033_ ) );
OAI21_X1 _13862_ ( .A(_06029_ ), .B1(_06031_ ), .B2(_06033_ ), .ZN(_00302_ ) );
CLKBUF_X2 _13863_ ( .A(_02027_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _13864_ ( .A(_01963_ ), .Z(_06034_ ) );
NOR3_X1 _13865_ ( .A1(_06034_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06035_ ) );
INV_X1 _13866_ ( .A(_01975_ ), .ZN(_06036_ ) );
BUF_X4 _13867_ ( .A(_06036_ ), .Z(_06037_ ) );
BUF_X4 _13868_ ( .A(_06037_ ), .Z(_06038_ ) );
BUF_X2 _13869_ ( .A(_06038_ ), .Z(_06039_ ) );
BUF_X4 _13870_ ( .A(_06039_ ), .Z(_06040_ ) );
BUF_X4 _13871_ ( .A(_06040_ ), .Z(_06041_ ) );
INV_X1 _13872_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06042_ ) );
INV_X1 _13873_ ( .A(_01965_ ), .ZN(_06043_ ) );
AOI211_X1 _13874_ ( .A(_06035_ ), .B(_06041_ ), .C1(_06042_ ), .C2(_06043_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _13875_ ( .A1(_06034_ ), .A2(fanout_net_3 ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06044_ ) );
INV_X1 _13876_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06045_ ) );
AOI211_X1 _13877_ ( .A(_06044_ ), .B(_06040_ ), .C1(_06045_ ), .C2(_06043_ ), .ZN(\io_master_araddr [0] ) );
OR3_X1 _13878_ ( .A1(_06034_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06046_ ) );
BUF_X4 _13879_ ( .A(_01965_ ), .Z(_06047_ ) );
OAI21_X1 _13880_ ( .A(_06046_ ), .B1(_06047_ ), .B2(\mylsu.araddr_tmp [15] ), .ZN(_06048_ ) );
BUF_X4 _13881_ ( .A(_01954_ ), .Z(_06049_ ) );
BUF_X4 _13882_ ( .A(_06049_ ), .Z(_06050_ ) );
BUF_X4 _13883_ ( .A(_06050_ ), .Z(_06051_ ) );
OAI22_X1 _13884_ ( .A1(_06041_ ), .A2(_06048_ ), .B1(_03463_ ), .B2(_06051_ ), .ZN(\io_master_araddr [15] ) );
OAI221_X1 _13885_ ( .A(\IF_ID_pc [14] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_06052_ ) );
OR3_X1 _13886_ ( .A1(_06034_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06053_ ) );
OAI211_X1 _13887_ ( .A(_01959_ ), .B(_06053_ ), .C1(\mylsu.araddr_tmp [14] ), .C2(_06047_ ), .ZN(_06054_ ) );
OAI21_X1 _13888_ ( .A(_06052_ ), .B1(\io_master_arburst [0] ), .B2(_06054_ ), .ZN(\io_master_araddr [14] ) );
NOR3_X1 _13889_ ( .A1(_06034_ ), .A2(_05307_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06055_ ) );
AOI21_X1 _13890_ ( .A(_06055_ ), .B1(_06043_ ), .B2(\mylsu.araddr_tmp [5] ), .ZN(_06056_ ) );
OAI22_X1 _13891_ ( .A1(_06041_ ), .A2(_06056_ ), .B1(_03512_ ), .B2(_06051_ ), .ZN(\io_master_araddr [5] ) );
OR3_X1 _13892_ ( .A1(_06034_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06057_ ) );
OAI21_X1 _13893_ ( .A(_06057_ ), .B1(_06047_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_06058_ ) );
OAI22_X1 _13894_ ( .A1(_06041_ ), .A2(_06058_ ), .B1(_03748_ ), .B2(_06051_ ), .ZN(\io_master_araddr [4] ) );
NOR2_X1 _13895_ ( .A1(_03899_ ), .A2(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06059_ ) );
NAND4_X1 _13896_ ( .A1(_06059_ ), .A2(_05304_ ), .A3(_02038_ ), .A4(_03855_ ), .ZN(_06060_ ) );
OAI21_X1 _13897_ ( .A(_06060_ ), .B1(_06047_ ), .B2(\mylsu.araddr_tmp [3] ), .ZN(_06061_ ) );
OAI22_X1 _13898_ ( .A1(_06041_ ), .A2(_06061_ ), .B1(_03756_ ), .B2(_06051_ ), .ZN(\io_master_araddr [3] ) );
INV_X1 _13899_ ( .A(_01974_ ), .ZN(\io_master_araddr [31] ) );
INV_X1 _13900_ ( .A(_01970_ ), .ZN(\io_master_araddr [30] ) );
INV_X1 _13901_ ( .A(_02008_ ), .ZN(\io_master_araddr [29] ) );
INV_X1 _13902_ ( .A(_01991_ ), .ZN(\io_master_araddr [28] ) );
INV_X1 _13903_ ( .A(_02012_ ), .ZN(\io_master_araddr [27] ) );
INV_X1 _13904_ ( .A(_01995_ ), .ZN(\io_master_araddr [26] ) );
INV_X1 _13905_ ( .A(_01979_ ), .ZN(\io_master_araddr [24] ) );
OR3_X1 _13906_ ( .A1(_06034_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06062_ ) );
OAI21_X1 _13907_ ( .A(_06062_ ), .B1(_06047_ ), .B2(\mylsu.araddr_tmp [13] ), .ZN(_06063_ ) );
OAI22_X1 _13908_ ( .A1(_06041_ ), .A2(_06063_ ), .B1(_03542_ ), .B2(_06051_ ), .ZN(\io_master_araddr [13] ) );
OAI221_X1 _13909_ ( .A(\IF_ID_pc [12] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_06064_ ) );
OR3_X1 _13910_ ( .A1(_06034_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06065_ ) );
OAI211_X1 _13911_ ( .A(_01959_ ), .B(_06065_ ), .C1(\mylsu.araddr_tmp [12] ), .C2(_06047_ ), .ZN(_06066_ ) );
OAI21_X1 _13912_ ( .A(_06064_ ), .B1(\io_master_arburst [0] ), .B2(_06066_ ), .ZN(\io_master_araddr [12] ) );
OAI221_X1 _13913_ ( .A(\IF_ID_pc [11] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_06067_ ) );
OR3_X1 _13914_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [11] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06068_ ) );
OAI211_X1 _13915_ ( .A(_01959_ ), .B(_06068_ ), .C1(\mylsu.araddr_tmp [11] ), .C2(_06047_ ), .ZN(_06069_ ) );
OAI21_X1 _13916_ ( .A(_06067_ ), .B1(\io_master_arburst [0] ), .B2(_06069_ ), .ZN(\io_master_araddr [11] ) );
OAI221_X1 _13917_ ( .A(\IF_ID_pc [10] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01967_ ), .C2(_01968_ ), .ZN(_06070_ ) );
OR3_X1 _13918_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06071_ ) );
OAI211_X1 _13919_ ( .A(_01959_ ), .B(_06071_ ), .C1(\mylsu.araddr_tmp [10] ), .C2(_01965_ ), .ZN(_06072_ ) );
OAI21_X1 _13920_ ( .A(_06070_ ), .B1(\io_master_arburst [0] ), .B2(_06072_ ), .ZN(\io_master_araddr [10] ) );
NOR3_X1 _13921_ ( .A1(_06034_ ), .A2(_03869_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06073_ ) );
AOI21_X1 _13922_ ( .A(_06073_ ), .B1(_06043_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06074_ ) );
OAI22_X1 _13923_ ( .A1(_06041_ ), .A2(_06074_ ), .B1(_03450_ ), .B2(_06051_ ), .ZN(\io_master_araddr [9] ) );
NAND4_X1 _13924_ ( .A1(_06059_ ), .A2(_03873_ ), .A3(_02038_ ), .A4(_03855_ ), .ZN(_06075_ ) );
OAI21_X1 _13925_ ( .A(_06075_ ), .B1(_06047_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_06076_ ) );
OAI22_X1 _13926_ ( .A1(_06041_ ), .A2(_06076_ ), .B1(_01803_ ), .B2(_06051_ ), .ZN(\io_master_araddr [8] ) );
OR3_X1 _13927_ ( .A1(_06034_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06077_ ) );
OAI21_X1 _13928_ ( .A(_06077_ ), .B1(_06047_ ), .B2(\mylsu.araddr_tmp [7] ), .ZN(_06078_ ) );
OAI22_X1 _13929_ ( .A1(_06041_ ), .A2(_06078_ ), .B1(_01852_ ), .B2(_06051_ ), .ZN(\io_master_araddr [7] ) );
NAND4_X1 _13930_ ( .A1(_06059_ ), .A2(_03876_ ), .A3(_02038_ ), .A4(_01941_ ), .ZN(_06079_ ) );
OAI21_X1 _13931_ ( .A(_06079_ ), .B1(_06047_ ), .B2(\mylsu.araddr_tmp [6] ), .ZN(_06080_ ) );
OAI22_X1 _13932_ ( .A1(_06041_ ), .A2(_06080_ ), .B1(_03478_ ), .B2(_06051_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _13933_ ( .A1(_01963_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06081_ ) );
OAI211_X1 _13934_ ( .A(_01959_ ), .B(_06081_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01965_ ), .ZN(_06082_ ) );
NOR2_X1 _13935_ ( .A1(_01953_ ), .A2(_06082_ ), .ZN(_06083_ ) );
BUF_X4 _13936_ ( .A(_06083_ ), .Z(_06084_ ) );
BUF_X4 _13937_ ( .A(_06084_ ), .Z(_06085_ ) );
BUF_X2 _13938_ ( .A(_06085_ ), .Z(\io_master_araddr [2] ) );
AND3_X1 _13939_ ( .A1(_06050_ ), .A2(\EX_LS_typ [3] ), .A3(_01959_ ), .ZN(\io_master_arsize [2] ) );
AND3_X1 _13940_ ( .A1(_06050_ ), .A2(\EX_LS_typ [1] ), .A3(_01959_ ), .ZN(\io_master_arsize [0] ) );
OAI22_X1 _13941_ ( .A1(_01938_ ), .A2(_01939_ ), .B1(_02030_ ), .B2(_01945_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _13942_ ( .A(_02074_ ), .B(_02075_ ), .C1(_02068_ ), .C2(_02071_ ), .ZN(io_master_arvalid ) );
AND2_X1 _13943_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ) );
AND2_X1 _13944_ ( .A1(_02051_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_06086_ ) );
BUF_X4 _13945_ ( .A(_06086_ ), .Z(_06087_ ) );
BUF_X4 _13946_ ( .A(_06087_ ), .Z(_06088_ ) );
MUX2_X1 _13947_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06088_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _13948_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06088_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _13949_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06088_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _13950_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06088_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _13951_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06088_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _13952_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06088_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _13953_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06088_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _13954_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06088_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _13955_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06088_ ), .Z(\io_master_awaddr [15] ) );
BUF_X4 _13956_ ( .A(_06087_ ), .Z(_06089_ ) );
MUX2_X1 _13957_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06089_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _13958_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06089_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _13959_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06089_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _13960_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06089_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _13961_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06089_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _13962_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06089_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _13963_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06089_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _13964_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06089_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _13965_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06089_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _13966_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06089_ ), .Z(\io_master_awaddr [6] ) );
BUF_X4 _13967_ ( .A(_06087_ ), .Z(_06090_ ) );
MUX2_X1 _13968_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06090_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _13969_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06090_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _13970_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06090_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _13971_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06090_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _13972_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06090_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _13973_ ( .A(\mylsu.awaddr_tmp [1] ), .B(\EX_LS_dest_csreg_mem [1] ), .S(_06090_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _13974_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_3 ), .S(_06090_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _13975_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06090_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _13976_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06090_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _13977_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06090_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _13978_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06087_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _13979_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06087_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _13980_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06087_ ), .Z(\io_master_awaddr [22] ) );
AND4_X1 _13981_ ( .A1(\EX_LS_typ [1] ), .A2(_02056_ ), .A3(_03853_ ), .A4(_02033_ ), .ZN(\io_master_awsize [0] ) );
NAND3_X1 _13982_ ( .A1(_02056_ ), .A2(_03853_ ), .A3(_02033_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _13983_ ( .A1(_02048_ ), .A2(_02059_ ), .A3(_06088_ ), .ZN(_06091_ ) );
NAND2_X1 _13984_ ( .A1(_06091_ ), .A2(_05995_ ), .ZN(io_master_awvalid ) );
INV_X1 _13985_ ( .A(\mylsu.state [2] ), .ZN(_06092_ ) );
INV_X1 _13986_ ( .A(\mylsu.state [1] ), .ZN(_06093_ ) );
NAND4_X1 _13987_ ( .A1(_06091_ ), .A2(_06092_ ), .A3(_05995_ ), .A4(_06093_ ), .ZN(io_master_bready ) );
NOR3_X1 _13988_ ( .A1(_01944_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_06094_ ) );
INV_X1 _13989_ ( .A(\mylsu.state [3] ), .ZN(_06095_ ) );
BUF_X2 _13990_ ( .A(_06095_ ), .Z(_06096_ ) );
NOR2_X1 _13991_ ( .A1(_03817_ ), .A2(\io_master_rid [0] ), .ZN(_06097_ ) );
NAND4_X1 _13992_ ( .A1(_06097_ ), .A2(io_master_rlast ), .A3(_03815_ ), .A4(_03816_ ), .ZN(_06098_ ) );
AOI21_X1 _13993_ ( .A(_06040_ ), .B1(_03814_ ), .B2(_06098_ ), .ZN(_06099_ ) );
AOI21_X1 _13994_ ( .A(_06096_ ), .B1(_06099_ ), .B2(_03830_ ), .ZN(_06100_ ) );
INV_X1 _13995_ ( .A(\io_master_bid [0] ), .ZN(_06101_ ) );
OR3_X1 _13996_ ( .A1(_06101_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bresp [1] ), .ZN(_06102_ ) );
INV_X1 _13997_ ( .A(\io_master_bid [2] ), .ZN(_06103_ ) );
INV_X1 _13998_ ( .A(\io_master_bresp [0] ), .ZN(_06104_ ) );
NAND4_X1 _13999_ ( .A1(_06103_ ), .A2(_06104_ ), .A3(\io_master_bid [1] ), .A4(io_master_bvalid ), .ZN(_06105_ ) );
NOR2_X1 _14000_ ( .A1(_06102_ ), .A2(_06105_ ), .ZN(_06106_ ) );
INV_X1 _14001_ ( .A(_06106_ ), .ZN(_06107_ ) );
AOI211_X1 _14002_ ( .A(_06094_ ), .B(_06100_ ), .C1(\mylsu.state [1] ), .C2(_06107_ ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _14003_ ( .A(_02061_ ), .B(_02065_ ), .C1(_02068_ ), .C2(_02071_ ), .ZN(io_master_rready ) );
MUX2_X1 _14004_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_3 ), .Z(_06108_ ) );
CLKBUF_X2 _14005_ ( .A(_05306_ ), .Z(_06109_ ) );
AND2_X1 _14006_ ( .A1(_06108_ ), .A2(_06109_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _14007_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_3 ), .Z(_06110_ ) );
AND2_X1 _14008_ ( .A1(_06110_ ), .A2(_06109_ ), .ZN(\io_master_wdata [14] ) );
INV_X1 _14009_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_06111_ ) );
NOR3_X1 _14010_ ( .A1(_06111_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [5] ) );
INV_X1 _14011_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_06112_ ) );
NOR3_X1 _14012_ ( .A1(_06112_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [4] ) );
INV_X1 _14013_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_06113_ ) );
NOR3_X1 _14014_ ( .A1(_06113_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14015_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_06114_ ) );
NOR3_X1 _14016_ ( .A1(_06114_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14017_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06115_ ) );
NOR3_X1 _14018_ ( .A1(_06115_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14019_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06116_ ) );
NOR3_X1 _14020_ ( .A1(_06116_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14021_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_3 ), .Z(_06117_ ) );
AND2_X1 _14022_ ( .A1(_06117_ ), .A2(_06109_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14023_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_3 ), .Z(_06118_ ) );
AND2_X1 _14024_ ( .A1(_06118_ ), .A2(_06109_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14025_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_3 ), .Z(_06119_ ) );
AND2_X1 _14026_ ( .A1(_06119_ ), .A2(_06109_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14027_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_3 ), .Z(_06120_ ) );
AND2_X1 _14028_ ( .A1(_06120_ ), .A2(_06109_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14029_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_3 ), .Z(_06121_ ) );
AND2_X1 _14030_ ( .A1(_06121_ ), .A2(_06109_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14031_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_3 ), .Z(_06122_ ) );
AND2_X1 _14032_ ( .A1(_06122_ ), .A2(_06109_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14033_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06123_ ) );
NOR3_X1 _14034_ ( .A1(_06123_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [7] ) );
NOR3_X1 _14035_ ( .A1(_05719_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14036_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_3 ), .Z(_06124_ ) );
MUX2_X1 _14037_ ( .A(_06124_ ), .B(_06108_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14038_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_3 ), .Z(_06125_ ) );
MUX2_X1 _14039_ ( .A(_06125_ ), .B(_06110_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [30] ) );
NOR2_X1 _14040_ ( .A1(_05306_ ), .A2(fanout_net_3 ), .ZN(_06126_ ) );
INV_X1 _14041_ ( .A(_06126_ ), .ZN(_06127_ ) );
OAI21_X1 _14042_ ( .A(_05306_ ), .B1(_03879_ ), .B2(\EX_LS_result_csreg_mem [13] ), .ZN(_06128_ ) );
NOR2_X1 _14043_ ( .A1(fanout_net_3 ), .A2(\EX_LS_result_csreg_mem [21] ), .ZN(_06129_ ) );
OAI22_X1 _14044_ ( .A1(_06127_ ), .A2(_06111_ ), .B1(_06128_ ), .B2(_06129_ ), .ZN(\io_master_wdata [21] ) );
OAI21_X1 _14045_ ( .A(_05306_ ), .B1(_03879_ ), .B2(\EX_LS_result_csreg_mem [12] ), .ZN(_06130_ ) );
NOR2_X1 _14046_ ( .A1(fanout_net_3 ), .A2(\EX_LS_result_csreg_mem [20] ), .ZN(_06131_ ) );
OAI22_X1 _14047_ ( .A1(_06127_ ), .A2(_06112_ ), .B1(_06130_ ), .B2(_06131_ ), .ZN(\io_master_wdata [20] ) );
OAI21_X1 _14048_ ( .A(_05306_ ), .B1(_03879_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_06132_ ) );
NOR2_X1 _14049_ ( .A1(fanout_net_3 ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_06133_ ) );
OAI22_X1 _14050_ ( .A1(_06127_ ), .A2(_06113_ ), .B1(_06132_ ), .B2(_06133_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _14051_ ( .A(_05306_ ), .B1(_03879_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_06134_ ) );
NOR2_X1 _14052_ ( .A1(fanout_net_3 ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_06135_ ) );
OAI22_X1 _14053_ ( .A1(_06127_ ), .A2(_06114_ ), .B1(_06134_ ), .B2(_06135_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _14054_ ( .A(_05306_ ), .B1(_03879_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_06136_ ) );
NOR2_X1 _14055_ ( .A1(fanout_net_3 ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_06137_ ) );
OAI22_X1 _14056_ ( .A1(_06127_ ), .A2(_06115_ ), .B1(_06136_ ), .B2(_06137_ ), .ZN(\io_master_wdata [17] ) );
INV_X1 _14057_ ( .A(\EX_LS_result_csreg_mem [16] ), .ZN(_06138_ ) );
INV_X1 _14058_ ( .A(\EX_LS_result_csreg_mem [8] ), .ZN(_06139_ ) );
MUX2_X1 _14059_ ( .A(_06138_ ), .B(_06139_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06140_ ) );
OAI22_X1 _14060_ ( .A1(_06140_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06127_ ), .B2(_06116_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14061_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06141_ ) );
MUX2_X1 _14062_ ( .A(_06141_ ), .B(_06117_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14063_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06142_ ) );
MUX2_X1 _14064_ ( .A(_06142_ ), .B(_06118_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14065_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06143_ ) );
MUX2_X1 _14066_ ( .A(_06143_ ), .B(_06119_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14067_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06144_ ) );
MUX2_X1 _14068_ ( .A(_06144_ ), .B(_06120_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14069_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06145_ ) );
MUX2_X1 _14070_ ( .A(_06145_ ), .B(_06121_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14071_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06146_ ) );
MUX2_X1 _14072_ ( .A(_06146_ ), .B(_06122_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [24] ) );
OAI21_X1 _14073_ ( .A(_05306_ ), .B1(_03879_ ), .B2(\EX_LS_result_csreg_mem [15] ), .ZN(_06147_ ) );
NOR2_X1 _14074_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [23] ), .ZN(_06148_ ) );
OAI22_X1 _14075_ ( .A1(_06127_ ), .A2(_06123_ ), .B1(_06147_ ), .B2(_06148_ ), .ZN(\io_master_wdata [23] ) );
OAI21_X1 _14076_ ( .A(_05306_ ), .B1(_03879_ ), .B2(\EX_LS_result_csreg_mem [14] ), .ZN(_06149_ ) );
NOR2_X1 _14077_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [22] ), .ZN(_06150_ ) );
OAI22_X1 _14078_ ( .A1(_06127_ ), .A2(_05719_ ), .B1(_06149_ ), .B2(_06150_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14079_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06151_ ) );
AND2_X1 _14080_ ( .A1(_06151_ ), .A2(_06109_ ), .ZN(\io_master_wstrb [1] ) );
NOR3_X1 _14081_ ( .A1(_02028_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14082_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06152_ ) );
MUX2_X1 _14083_ ( .A(_06152_ ), .B(_06151_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14084_ ( .A1(_06109_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_06153_ ) );
OAI221_X1 _14085_ ( .A(_06153_ ), .B1(_02053_ ), .B2(_02030_ ), .C1(_06127_ ), .C2(_02028_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _14086_ ( .A1(_06091_ ), .A2(_06092_ ), .ZN(io_master_wvalid ) );
MUX2_X1 _14087_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14088_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14089_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14090_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
INV_X1 _14091_ ( .A(_02060_ ), .ZN(_06154_ ) );
NOR2_X1 _14092_ ( .A1(_06018_ ), .A2(exception_quest_IDU ), .ZN(_06155_ ) );
NOR2_X1 _14093_ ( .A1(_06154_ ), .A2(_06155_ ), .ZN(_06156_ ) );
BUF_X4 _14094_ ( .A(_06156_ ), .Z(_06157_ ) );
MUX2_X1 _14095_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14096_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14097_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14098_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14099_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14100_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14101_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14102_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14103_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14104_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_06157_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14105_ ( .A(_06156_ ), .Z(_06158_ ) );
MUX2_X1 _14106_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14107_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14108_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14109_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14110_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14111_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14112_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14113_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14114_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14115_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_06158_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14116_ ( .A(_06156_ ), .Z(_06159_ ) );
MUX2_X1 _14117_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14118_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14119_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14120_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14121_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14122_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14123_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14124_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14125_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14126_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14127_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_06156_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14128_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_06156_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
XNOR2_X1 _14129_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06160_ ) );
XNOR2_X1 _14130_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06161_ ) );
XNOR2_X1 _14131_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06162_ ) );
XNOR2_X1 _14132_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06163_ ) );
NAND4_X1 _14133_ ( .A1(_06160_ ), .A2(_06161_ ), .A3(_06162_ ), .A4(_06163_ ), .ZN(_06164_ ) );
XNOR2_X1 _14134_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06165_ ) );
XNOR2_X1 _14135_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06166_ ) );
NAND2_X1 _14136_ ( .A1(_06165_ ), .A2(_06166_ ), .ZN(_06167_ ) );
XOR2_X1 _14137_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .Z(_06168_ ) );
XOR2_X1 _14138_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .Z(_06169_ ) );
NOR4_X1 _14139_ ( .A1(_06164_ ), .A2(_06167_ ), .A3(_06168_ ), .A4(_06169_ ), .ZN(_06170_ ) );
XNOR2_X1 _14140_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06171_ ) );
XNOR2_X1 _14141_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06172_ ) );
XNOR2_X1 _14142_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06173_ ) );
XNOR2_X1 _14143_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06174_ ) );
AND4_X1 _14144_ ( .A1(_06171_ ), .A2(_06172_ ), .A3(_06173_ ), .A4(_06174_ ), .ZN(_06175_ ) );
XNOR2_X1 _14145_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06176_ ) );
XNOR2_X1 _14146_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06177_ ) );
XNOR2_X1 _14147_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06178_ ) );
XNOR2_X1 _14148_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06179_ ) );
AND4_X1 _14149_ ( .A1(_06176_ ), .A2(_06177_ ), .A3(_06178_ ), .A4(_06179_ ), .ZN(_06180_ ) );
NAND3_X1 _14150_ ( .A1(_06170_ ), .A2(_06175_ ), .A3(_06180_ ), .ZN(_06181_ ) );
XNOR2_X1 _14151_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_06182_ ) );
XNOR2_X1 _14152_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_06183_ ) );
XNOR2_X1 _14153_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_06184_ ) );
XNOR2_X1 _14154_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_06185_ ) );
NAND4_X1 _14155_ ( .A1(_06182_ ), .A2(_06183_ ), .A3(_06184_ ), .A4(_06185_ ), .ZN(_06186_ ) );
XNOR2_X1 _14156_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06187_ ) );
XNOR2_X1 _14157_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06188_ ) );
NAND2_X1 _14158_ ( .A1(_06187_ ), .A2(_06188_ ), .ZN(_06189_ ) );
XOR2_X1 _14159_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .Z(_06190_ ) );
XOR2_X1 _14160_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .Z(_06191_ ) );
NOR4_X1 _14161_ ( .A1(_06186_ ), .A2(_06189_ ), .A3(_06190_ ), .A4(_06191_ ), .ZN(_06192_ ) );
XNOR2_X1 _14162_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06193_ ) );
XNOR2_X1 _14163_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06194_ ) );
XNOR2_X1 _14164_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06195_ ) );
XNOR2_X1 _14165_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06196_ ) );
NAND4_X1 _14166_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(_06195_ ), .A4(_06196_ ), .ZN(_06197_ ) );
XNOR2_X1 _14167_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06198_ ) );
XNOR2_X1 _14168_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06199_ ) );
XNOR2_X1 _14169_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06200_ ) );
XNOR2_X1 _14170_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06201_ ) );
NAND4_X1 _14171_ ( .A1(_06198_ ), .A2(_06199_ ), .A3(_06200_ ), .A4(_06201_ ), .ZN(_06202_ ) );
NOR2_X1 _14172_ ( .A1(_06197_ ), .A2(_06202_ ), .ZN(_06203_ ) );
NAND2_X1 _14173_ ( .A1(_06192_ ), .A2(_06203_ ), .ZN(_06204_ ) );
NOR3_X1 _14174_ ( .A1(_06181_ ), .A2(_06204_ ), .A3(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06205_ ) );
NAND3_X1 _14175_ ( .A1(_02048_ ), .A2(_02059_ ), .A3(_02091_ ), .ZN(_06206_ ) );
MUX2_X1 _14176_ ( .A(_06205_ ), .B(_06206_ ), .S(_02092_ ), .Z(\myec.state_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _14177_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06207_ ) );
NAND2_X1 _14178_ ( .A1(_06207_ ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06208_ ) );
NOR2_X1 _14179_ ( .A1(_06208_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06209_ ) );
NOR2_X1 _14180_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06210_ ) );
AND3_X1 _14181_ ( .A1(_06210_ ), .A2(\LS_WB_waddr_csreg [9] ), .A3(\LS_WB_waddr_csreg [8] ), .ZN(_06211_ ) );
NOR2_X1 _14182_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_06212_ ) );
AND3_X1 _14183_ ( .A1(_06209_ ), .A2(_06211_ ), .A3(_06212_ ), .ZN(_06213_ ) );
INV_X1 _14184_ ( .A(_06213_ ), .ZN(_06214_ ) );
NOR3_X1 _14185_ ( .A1(reset ), .A2(excp_written ), .A3(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_B ), .ZN(_06215_ ) );
INV_X1 _14186_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_06216_ ) );
NAND3_X1 _14187_ ( .A1(_06215_ ), .A2(_06216_ ), .A3(\LS_WB_waddr_csreg [0] ), .ZN(_06217_ ) );
NOR2_X1 _14188_ ( .A1(_06214_ ), .A2(_06217_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14189_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .A3(\LS_WB_waddr_csreg [5] ), .A4(\LS_WB_waddr_csreg [4] ), .ZN(_06218_ ) );
NOR4_X1 _14190_ ( .A1(\LS_WB_waddr_csreg [1] ), .A2(\LS_WB_waddr_csreg [0] ), .A3(\LS_WB_waddr_csreg [3] ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_06219_ ) );
AND4_X1 _14191_ ( .A1(_06215_ ), .A2(_06211_ ), .A3(_06218_ ), .A4(_06219_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _14192_ ( .A1(_06211_ ), .A2(_06218_ ), .ZN(_06220_ ) );
INV_X1 _14193_ ( .A(\LS_WB_waddr_csreg [2] ), .ZN(_06221_ ) );
NOR4_X1 _14194_ ( .A1(_06220_ ), .A2(_06217_ ), .A3(\LS_WB_waddr_csreg [3] ), .A4(_06221_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND3_X1 _14195_ ( .A1(_01535_ ), .A2(\LS_WB_wen_csreg [7] ), .A3(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06222_ ) );
NOR4_X1 _14196_ ( .A1(_06216_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(\LS_WB_waddr_csreg [3] ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_06223_ ) );
NAND3_X1 _14197_ ( .A1(_06209_ ), .A2(_06211_ ), .A3(_06223_ ), .ZN(_06224_ ) );
AOI21_X1 _14198_ ( .A(_06222_ ), .B1(_06224_ ), .B2(_02078_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NAND2_X1 _14199_ ( .A1(_05809_ ), .A2(_03019_ ), .ZN(_06225_ ) );
AND2_X2 _14200_ ( .A1(_03008_ ), .A2(_03889_ ), .ZN(_06226_ ) );
INV_X1 _14201_ ( .A(_06226_ ), .ZN(_06227_ ) );
BUF_X4 _14202_ ( .A(_06227_ ), .Z(_06228_ ) );
BUF_X4 _14203_ ( .A(_06228_ ), .Z(_06229_ ) );
OAI21_X1 _14204_ ( .A(_06225_ ), .B1(_05248_ ), .B2(_06229_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _14205_ ( .A(_04743_ ), .B(\ID_EX_imm [0] ), .ZN(_06230_ ) );
AND2_X2 _14206_ ( .A1(_03342_ ), .A2(\ID_EX_typ [7] ), .ZN(_06231_ ) );
INV_X1 _14207_ ( .A(_06231_ ), .ZN(_06232_ ) );
BUF_X4 _14208_ ( .A(_06232_ ), .Z(_06233_ ) );
BUF_X4 _14209_ ( .A(_06233_ ), .Z(_06234_ ) );
NAND2_X1 _14210_ ( .A1(_06230_ ), .A2(_06234_ ), .ZN(_06235_ ) );
BUF_X4 _14211_ ( .A(_06227_ ), .Z(_06236_ ) );
BUF_X4 _14212_ ( .A(_06236_ ), .Z(_06237_ ) );
MUX2_X1 _14213_ ( .A(\ID_EX_csr [0] ), .B(_06235_ ), .S(_06237_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
BUF_X4 _14214_ ( .A(_06232_ ), .Z(_06238_ ) );
AND2_X1 _14215_ ( .A1(_05642_ ), .A2(_06238_ ), .ZN(_06239_ ) );
MUX2_X1 _14216_ ( .A(\ID_EX_csr [10] ), .B(_06239_ ), .S(_06237_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
NOR4_X1 _14217_ ( .A1(_03343_ ), .A2(_03898_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [9] ), .ZN(_06240_ ) );
AOI21_X1 _14218_ ( .A(_06240_ ), .B1(_05663_ ), .B2(_03019_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR2_X1 _14219_ ( .A1(_05681_ ), .A2(_06231_ ), .ZN(_06241_ ) );
MUX2_X1 _14220_ ( .A(\ID_EX_csr [8] ), .B(_06241_ ), .S(_06237_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _14221_ ( .A1(_05704_ ), .A2(_03019_ ), .ZN(_06242_ ) );
OAI21_X1 _14222_ ( .A(_06242_ ), .B1(_05234_ ), .B2(_06229_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
NOR2_X1 _14223_ ( .A1(_05723_ ), .A2(_03008_ ), .ZN(_06243_ ) );
BUF_X4 _14224_ ( .A(_06226_ ), .Z(_06244_ ) );
BUF_X4 _14225_ ( .A(_06244_ ), .Z(_06245_ ) );
AOI21_X1 _14226_ ( .A(_06243_ ), .B1(_05302_ ), .B2(_06245_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14227_ ( .A1(_05741_ ), .A2(_03019_ ), .ZN(_06246_ ) );
OAI21_X1 _14228_ ( .A(_06246_ ), .B1(_05252_ ), .B2(_06229_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
AND2_X1 _14229_ ( .A1(_05761_ ), .A2(_06233_ ), .ZN(_06247_ ) );
MUX2_X1 _14230_ ( .A(\ID_EX_csr [4] ), .B(_06247_ ), .S(_06237_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _14231_ ( .A1(_05778_ ), .A2(_03018_ ), .ZN(_06248_ ) );
BUF_X4 _14232_ ( .A(_06236_ ), .Z(_06249_ ) );
OAI21_X1 _14233_ ( .A(_06248_ ), .B1(_05242_ ), .B2(_06249_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _14234_ ( .A1(_05794_ ), .A2(_03018_ ), .ZN(_06250_ ) );
OAI21_X1 _14235_ ( .A(_06250_ ), .B1(_05243_ ), .B2(_06249_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
AND2_X1 _14236_ ( .A1(_05605_ ), .A2(_06233_ ), .ZN(_06251_ ) );
MUX2_X1 _14237_ ( .A(\ID_EX_csr [11] ), .B(_06251_ ), .S(_06228_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X2 _14238_ ( .A(_06227_ ), .Z(_06252_ ) );
NAND2_X1 _14239_ ( .A1(_02357_ ), .A2(fanout_net_4 ), .ZN(_06253_ ) );
AND2_X1 _14240_ ( .A1(_05958_ ), .A2(_05960_ ), .ZN(_06254_ ) );
OAI221_X1 _14241_ ( .A(_06253_ ), .B1(_06254_ ), .B2(_04869_ ), .C1(fanout_net_4 ), .C2(_04477_ ), .ZN(_06255_ ) );
NOR2_X1 _14242_ ( .A1(_04867_ ), .A2(\ID_EX_typ [2] ), .ZN(_06256_ ) );
BUF_X2 _14243_ ( .A(_06256_ ), .Z(_06257_ ) );
NAND3_X1 _14244_ ( .A1(_05958_ ), .A2(_06257_ ), .A3(_05960_ ), .ZN(_06258_ ) );
AOI21_X1 _14245_ ( .A(_06252_ ), .B1(_06255_ ), .B2(_06258_ ), .ZN(_06259_ ) );
AND3_X1 _14246_ ( .A1(_03342_ ), .A2(_05945_ ), .A3(\ID_EX_typ [7] ), .ZN(_06260_ ) );
AOI211_X1 _14247_ ( .A(_06244_ ), .B(_06260_ ), .C1(_04476_ ), .C2(_06234_ ), .ZN(_06261_ ) );
OR2_X1 _14248_ ( .A1(_06259_ ), .A2(_06261_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
INV_X2 _14249_ ( .A(_06256_ ), .ZN(_06262_ ) );
BUF_X2 _14250_ ( .A(_06262_ ), .Z(_06263_ ) );
AOI21_X1 _14251_ ( .A(_06263_ ), .B1(_05366_ ), .B2(_05367_ ), .ZN(_06264_ ) );
NAND3_X1 _14252_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_05428_ ), .ZN(_06265_ ) );
AND2_X1 _14253_ ( .A1(_05366_ ), .A2(_06265_ ), .ZN(_06266_ ) );
AOI22_X1 _14254_ ( .A1(_06266_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02383_ ), .ZN(_06267_ ) );
NAND3_X1 _14255_ ( .A1(_02380_ ), .A2(_02381_ ), .A3(_05406_ ), .ZN(_06268_ ) );
AOI211_X1 _14256_ ( .A(_06252_ ), .B(_06264_ ), .C1(_06267_ ), .C2(_06268_ ), .ZN(_06269_ ) );
MUX2_X1 _14257_ ( .A(_05943_ ), .B(_04452_ ), .S(_06238_ ), .Z(_06270_ ) );
AOI21_X1 _14258_ ( .A(_06269_ ), .B1(_06229_ ), .B2(_06270_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
OR3_X1 _14259_ ( .A1(_05547_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_05535_ ), .ZN(_06271_ ) );
NAND3_X1 _14260_ ( .A1(_05321_ ), .A2(\mepc [19] ), .A3(_05389_ ), .ZN(_06272_ ) );
NAND4_X1 _14261_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [19] ), .A4(_05444_ ), .ZN(_06273_ ) );
NAND4_X1 _14262_ ( .A1(_05835_ ), .A2(_06272_ ), .A3(_05388_ ), .A4(_06273_ ), .ZN(_06274_ ) );
INV_X1 _14263_ ( .A(_05398_ ), .ZN(_06275_ ) );
OAI21_X1 _14264_ ( .A(_06275_ ), .B1(_05547_ ), .B2(_05536_ ), .ZN(_06276_ ) );
OAI21_X1 _14265_ ( .A(_06271_ ), .B1(_06274_ ), .B2(_06276_ ), .ZN(_06277_ ) );
AOI22_X1 _14266_ ( .A1(_06277_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02430_ ), .ZN(_06278_ ) );
BUF_X4 _14267_ ( .A(_06226_ ), .Z(_06279_ ) );
OAI211_X1 _14268_ ( .A(_06278_ ), .B(_06279_ ), .C1(fanout_net_4 ), .C2(_04330_ ), .ZN(_06280_ ) );
OR3_X1 _14269_ ( .A1(_06277_ ), .A2(_06263_ ), .A3(_06236_ ), .ZN(_06281_ ) );
MUX2_X1 _14270_ ( .A(_04010_ ), .B(_04328_ ), .S(_06233_ ), .Z(_06282_ ) );
OAI211_X1 _14271_ ( .A(_06280_ ), .B(_06281_ ), .C1(_06245_ ), .C2(_06282_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
NAND4_X1 _14272_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_03840_ ), .A4(_05401_ ), .ZN(_06283_ ) );
AOI21_X1 _14273_ ( .A(_06263_ ), .B1(_05426_ ), .B2(_06283_ ), .ZN(_06284_ ) );
NOR2_X1 _14274_ ( .A1(_05405_ ), .A2(\ID_EX_imm [18] ), .ZN(_06285_ ) );
AOI21_X1 _14275_ ( .A(_06285_ ), .B1(_05430_ ), .B2(\ID_EX_typ [2] ), .ZN(_06286_ ) );
NAND3_X1 _14276_ ( .A1(_02404_ ), .A2(_02405_ ), .A3(_05406_ ), .ZN(_06287_ ) );
AOI211_X1 _14277_ ( .A(_06252_ ), .B(_06284_ ), .C1(_06286_ ), .C2(_06287_ ), .ZN(_06288_ ) );
MUX2_X1 _14278_ ( .A(_05410_ ), .B(_04305_ ), .S(_06238_ ), .Z(_06289_ ) );
AOI21_X1 _14279_ ( .A(_06288_ ), .B1(_06229_ ), .B2(_06289_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
AOI21_X1 _14280_ ( .A(fanout_net_4 ), .B1(_02455_ ), .B2(_02457_ ), .ZN(_06290_ ) );
AND2_X1 _14281_ ( .A1(fanout_net_4 ), .A2(\ID_EX_imm [17] ), .ZN(_06291_ ) );
BUF_X4 _14282_ ( .A(_04869_ ), .Z(_06292_ ) );
OAI221_X1 _14283_ ( .A(_06244_ ), .B1(_06290_ ), .B2(_06291_ ), .C1(_05449_ ), .C2(_06292_ ), .ZN(_06293_ ) );
NAND4_X1 _14284_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_05736_ ), .A4(_05401_ ), .ZN(_06294_ ) );
AOI21_X1 _14285_ ( .A(_06236_ ), .B1(_05446_ ), .B2(_06294_ ), .ZN(_06295_ ) );
NAND2_X1 _14286_ ( .A1(_06295_ ), .A2(_06257_ ), .ZN(_06296_ ) );
AND3_X1 _14287_ ( .A1(_03342_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_typ [7] ), .ZN(_06297_ ) );
AOI21_X1 _14288_ ( .A(_06297_ ), .B1(_04356_ ), .B2(_06234_ ), .ZN(_06298_ ) );
OAI211_X1 _14289_ ( .A(_06293_ ), .B(_06296_ ), .C1(_06245_ ), .C2(_06298_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _14290_ ( .A1(_05320_ ), .A2(\mepc [16] ), .A3(_05417_ ), .ZN(_06299_ ) );
NAND4_X1 _14291_ ( .A1(_05330_ ), .A2(_05327_ ), .A3(_05393_ ), .A4(\mycsreg.CSReg[0][16] ), .ZN(_06300_ ) );
AND3_X1 _14292_ ( .A1(_05470_ ), .A2(_06299_ ), .A3(_06300_ ), .ZN(_06301_ ) );
NAND4_X1 _14293_ ( .A1(_05326_ ), .A2(_05474_ ), .A3(_05441_ ), .A4(\mtvec [16] ), .ZN(_06302_ ) );
NAND3_X1 _14294_ ( .A1(_06301_ ), .A2(_05513_ ), .A3(_06302_ ), .ZN(_06303_ ) );
NAND2_X1 _14295_ ( .A1(_05314_ ), .A2(_06303_ ), .ZN(_06304_ ) );
NAND3_X1 _14296_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [16] ), .A3(_05428_ ), .ZN(_06305_ ) );
AOI21_X1 _14297_ ( .A(_06262_ ), .B1(_06304_ ), .B2(_06305_ ), .ZN(_06306_ ) );
AND2_X1 _14298_ ( .A1(_06304_ ), .A2(_06305_ ), .ZN(_06307_ ) );
AOI22_X1 _14299_ ( .A1(_06307_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02481_ ), .ZN(_06308_ ) );
NAND3_X1 _14300_ ( .A1(_02478_ ), .A2(_02479_ ), .A3(_05406_ ), .ZN(_06309_ ) );
AOI211_X1 _14301_ ( .A(_06252_ ), .B(_06306_ ), .C1(_06308_ ), .C2(_06309_ ), .ZN(_06310_ ) );
MUX2_X1 _14302_ ( .A(_05458_ ), .B(_04378_ ), .S(_06238_ ), .Z(_06311_ ) );
AOI21_X1 _14303_ ( .A(_06310_ ), .B1(_06229_ ), .B2(_06311_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
NAND4_X1 _14304_ ( .A1(_05400_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_03840_ ), .A4(_05401_ ), .ZN(_06312_ ) );
AOI21_X1 _14305_ ( .A(_06263_ ), .B1(_05499_ ), .B2(_06312_ ), .ZN(_06313_ ) );
NOR2_X1 _14306_ ( .A1(_05433_ ), .A2(\ID_EX_imm [15] ), .ZN(_06314_ ) );
AOI21_X1 _14307_ ( .A(_06314_ ), .B1(_05501_ ), .B2(\ID_EX_typ [2] ), .ZN(_06315_ ) );
NAND3_X1 _14308_ ( .A1(_02501_ ), .A2(_05623_ ), .A3(_02502_ ), .ZN(_06316_ ) );
AOI211_X1 _14309_ ( .A(_06228_ ), .B(_06313_ ), .C1(_06315_ ), .C2(_06316_ ), .ZN(_06317_ ) );
AND4_X1 _14310_ ( .A1(\ID_EX_pc [15] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06318_ ) );
AOI211_X1 _14311_ ( .A(_06244_ ), .B(_06318_ ), .C1(_05138_ ), .C2(_06234_ ), .ZN(_06319_ ) );
NOR2_X1 _14312_ ( .A1(_06317_ ), .A2(_06319_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _14313_ ( .A(_06263_ ), .B1(_05516_ ), .B2(_05517_ ), .ZN(_06320_ ) );
AOI22_X1 _14314_ ( .A1(_05518_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02527_ ), .ZN(_06321_ ) );
NAND3_X1 _14315_ ( .A1(_02523_ ), .A2(_02524_ ), .A3(_05884_ ), .ZN(_06322_ ) );
AOI211_X1 _14316_ ( .A(_06228_ ), .B(_06320_ ), .C1(_06321_ ), .C2(_06322_ ), .ZN(_06323_ ) );
AND4_X1 _14317_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06324_ ) );
AOI211_X1 _14318_ ( .A(_06244_ ), .B(_06324_ ), .C1(_04622_ ), .C2(_06234_ ), .ZN(_06325_ ) );
NOR2_X1 _14319_ ( .A1(_06323_ ), .A2(_06325_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OR3_X1 _14320_ ( .A1(_05547_ ), .A2(\EX_LS_result_csreg_mem [13] ), .A3(_05536_ ), .ZN(_06326_ ) );
OAI211_X1 _14321_ ( .A(_06257_ ), .B(_06326_ ), .C1(_05537_ ), .C2(_05545_ ), .ZN(_06327_ ) );
OAI22_X1 _14322_ ( .A1(_05549_ ), .A2(_06292_ ), .B1(_05433_ ), .B2(\ID_EX_imm [13] ), .ZN(_06328_ ) );
AND3_X1 _14323_ ( .A1(_02549_ ), .A2(_05433_ ), .A3(_02550_ ), .ZN(_06329_ ) );
OAI211_X1 _14324_ ( .A(_06244_ ), .B(_06327_ ), .C1(_06328_ ), .C2(_06329_ ), .ZN(_06330_ ) );
NAND4_X1 _14325_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06331_ ) );
OAI211_X1 _14326_ ( .A(_06228_ ), .B(_06331_ ), .C1(_04668_ ), .C2(_06231_ ), .ZN(_06332_ ) );
AND2_X1 _14327_ ( .A1(_06330_ ), .A2(_06332_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AOI21_X1 _14328_ ( .A(_06262_ ), .B1(_05572_ ), .B2(_05573_ ), .ZN(_06333_ ) );
AOI22_X1 _14329_ ( .A1(_05574_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02575_ ), .ZN(_06334_ ) );
NAND3_X1 _14330_ ( .A1(_02572_ ), .A2(_02573_ ), .A3(_05406_ ), .ZN(_06335_ ) );
AOI211_X1 _14331_ ( .A(_06252_ ), .B(_06333_ ), .C1(_06334_ ), .C2(_06335_ ), .ZN(_06336_ ) );
MUX2_X1 _14332_ ( .A(_05561_ ), .B(_04645_ ), .S(_06238_ ), .Z(_06337_ ) );
AOI21_X1 _14333_ ( .A(_06336_ ), .B1(_06229_ ), .B2(_06337_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
INV_X1 _14334_ ( .A(_05277_ ), .ZN(_06338_ ) );
AOI22_X1 _14335_ ( .A1(_06338_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02173_ ), .ZN(_06339_ ) );
OAI211_X1 _14336_ ( .A(_06279_ ), .B(_06339_ ), .C1(_05187_ ), .C2(fanout_net_4 ), .ZN(_06340_ ) );
BUF_X4 _14337_ ( .A(_06226_ ), .Z(_06341_ ) );
NAND3_X1 _14338_ ( .A1(_05277_ ), .A2(_06257_ ), .A3(_06341_ ), .ZN(_06342_ ) );
MUX2_X1 _14339_ ( .A(_05966_ ), .B(_04102_ ), .S(_06233_ ), .Z(_06343_ ) );
OAI211_X1 _14340_ ( .A(_06340_ ), .B(_06342_ ), .C1(_06245_ ), .C2(_06343_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
AOI21_X1 _14341_ ( .A(_06263_ ), .B1(_05586_ ), .B2(_05587_ ), .ZN(_06344_ ) );
AOI22_X1 _14342_ ( .A1(_05588_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02671_ ), .ZN(_06345_ ) );
NAND3_X1 _14343_ ( .A1(_02668_ ), .A2(_02669_ ), .A3(_05884_ ), .ZN(_06346_ ) );
AOI211_X1 _14344_ ( .A(_06228_ ), .B(_06344_ ), .C1(_06345_ ), .C2(_06346_ ), .ZN(_06347_ ) );
AND4_X1 _14345_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06348_ ) );
AOI211_X1 _14346_ ( .A(_06244_ ), .B(_06348_ ), .C1(_04526_ ), .C2(_06234_ ), .ZN(_06349_ ) );
NOR2_X1 _14347_ ( .A1(_06347_ ), .A2(_06349_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _14348_ ( .A(_06262_ ), .B1(_05638_ ), .B2(_05639_ ), .ZN(_06350_ ) );
NAND3_X1 _14349_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_05428_ ), .ZN(_06351_ ) );
AND2_X1 _14350_ ( .A1(_05638_ ), .A2(_06351_ ), .ZN(_06352_ ) );
AOI22_X1 _14351_ ( .A1(_06352_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_4 ), .B2(_02648_ ), .ZN(_06353_ ) );
NAND3_X1 _14352_ ( .A1(_02645_ ), .A2(_02646_ ), .A3(_05433_ ), .ZN(_06354_ ) );
AOI211_X1 _14353_ ( .A(_06252_ ), .B(_06350_ ), .C1(_06353_ ), .C2(_06354_ ), .ZN(_06355_ ) );
MUX2_X1 _14354_ ( .A(_05626_ ), .B(_04503_ ), .S(_06238_ ), .Z(_06356_ ) );
AOI21_X1 _14355_ ( .A(_06355_ ), .B1(_06229_ ), .B2(_06356_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
AOI21_X1 _14356_ ( .A(_06262_ ), .B1(_05650_ ), .B2(_05651_ ), .ZN(_06357_ ) );
AOI21_X1 _14357_ ( .A(_06357_ ), .B1(fanout_net_4 ), .B2(\ID_EX_imm [9] ), .ZN(_06358_ ) );
NAND2_X1 _14358_ ( .A1(_02624_ ), .A2(_05405_ ), .ZN(_06359_ ) );
AOI221_X4 _14359_ ( .A(_06227_ ), .B1(\ID_EX_typ [2] ), .B2(_05652_ ), .C1(_06358_ ), .C2(_06359_ ), .ZN(_06360_ ) );
NOR4_X1 _14360_ ( .A1(_03343_ ), .A2(_03898_ ), .A3(_03889_ ), .A4(\ID_EX_pc [9] ), .ZN(_06361_ ) );
AOI211_X1 _14361_ ( .A(_06226_ ), .B(_06361_ ), .C1(_04571_ ), .C2(_06238_ ), .ZN(_06362_ ) );
OR2_X1 _14362_ ( .A1(_06360_ ), .A2(_06362_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
NAND2_X1 _14363_ ( .A1(_02601_ ), .A2(fanout_net_4 ), .ZN(_06363_ ) );
OAI221_X1 _14364_ ( .A(_06363_ ), .B1(fanout_net_4 ), .B2(_02600_ ), .C1(_05675_ ), .C2(_06292_ ), .ZN(_06364_ ) );
OR2_X1 _14365_ ( .A1(_05674_ ), .A2(_06263_ ), .ZN(_06365_ ) );
NAND3_X1 _14366_ ( .A1(_06364_ ), .A2(_06279_ ), .A3(_06365_ ), .ZN(_06366_ ) );
NAND4_X1 _14367_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06367_ ) );
OAI211_X1 _14368_ ( .A(_06228_ ), .B(_06367_ ), .C1(_04549_ ), .C2(_06231_ ), .ZN(_06368_ ) );
AND2_X1 _14369_ ( .A1(_06366_ ), .A2(_06368_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
AOI22_X1 _14370_ ( .A1(_05692_ ), .A2(_06257_ ), .B1(fanout_net_4 ), .B2(\ID_EX_imm [7] ), .ZN(_06369_ ) );
INV_X1 _14371_ ( .A(_02816_ ), .ZN(_06370_ ) );
OAI21_X1 _14372_ ( .A(_06369_ ), .B1(_06370_ ), .B2(\ID_EX_typ [0] ), .ZN(_06371_ ) );
BUF_X4 _14373_ ( .A(_06244_ ), .Z(_06372_ ) );
OAI211_X1 _14374_ ( .A(_06371_ ), .B(_06372_ ), .C1(_06292_ ), .C2(_05692_ ), .ZN(_06373_ ) );
BUF_X4 _14375_ ( .A(_06236_ ), .Z(_06374_ ) );
OR4_X1 _14376_ ( .A1(\ID_EX_pc [7] ), .A2(_03343_ ), .A3(_03898_ ), .A4(_03889_ ), .ZN(_06375_ ) );
OAI211_X1 _14377_ ( .A(_06374_ ), .B(_06375_ ), .C1(_04814_ ), .C2(_06231_ ), .ZN(_06376_ ) );
NAND2_X1 _14378_ ( .A1(_06373_ ), .A2(_06376_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _14379_ ( .A1(_05721_ ), .A2(_04869_ ), .B1(_05405_ ), .B2(\ID_EX_imm [6] ), .ZN(_06377_ ) );
AOI21_X1 _14380_ ( .A(_06377_ ), .B1(_05623_ ), .B2(_02870_ ), .ZN(_06378_ ) );
NOR3_X1 _14381_ ( .A1(_05718_ ), .A2(_06263_ ), .A3(_05720_ ), .ZN(_06379_ ) );
OAI21_X1 _14382_ ( .A(_06372_ ), .B1(_06378_ ), .B2(_06379_ ), .ZN(_06380_ ) );
MUX2_X1 _14383_ ( .A(_05709_ ), .B(_04836_ ), .S(_06238_ ), .Z(_06381_ ) );
OAI21_X1 _14384_ ( .A(_06380_ ), .B1(_06245_ ), .B2(_06381_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
AND3_X1 _14385_ ( .A1(_05354_ ), .A2(\mepc [5] ), .A3(_05257_ ), .ZN(_06382_ ) );
INV_X1 _14386_ ( .A(_06382_ ), .ZN(_06383_ ) );
NAND4_X1 _14387_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [5] ), .A4(_05265_ ), .ZN(_06384_ ) );
NAND4_X1 _14388_ ( .A1(_06383_ ), .A2(_05542_ ), .A3(_05730_ ), .A4(_06384_ ), .ZN(_06385_ ) );
NOR3_X1 _14389_ ( .A1(_06385_ ), .A2(_05744_ ), .A3(_05734_ ), .ZN(_06386_ ) );
NOR3_X1 _14390_ ( .A1(_05547_ ), .A2(\EX_LS_result_csreg_mem [5] ), .A3(_05536_ ), .ZN(_06387_ ) );
NOR2_X1 _14391_ ( .A1(_06386_ ), .A2(_06387_ ), .ZN(_06388_ ) );
OAI22_X1 _14392_ ( .A1(_06388_ ), .A2(_04869_ ), .B1(_05405_ ), .B2(\ID_EX_imm [5] ), .ZN(_06389_ ) );
AOI21_X1 _14393_ ( .A(_06389_ ), .B1(_05623_ ), .B2(_02875_ ), .ZN(_06390_ ) );
OR3_X1 _14394_ ( .A1(_06386_ ), .A2(_06262_ ), .A3(_06387_ ), .ZN(_06391_ ) );
INV_X1 _14395_ ( .A(_06391_ ), .ZN(_06392_ ) );
OAI21_X1 _14396_ ( .A(_06341_ ), .B1(_06390_ ), .B2(_06392_ ), .ZN(_06393_ ) );
AND4_X1 _14397_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06394_ ) );
AOI21_X1 _14398_ ( .A(_06394_ ), .B1(_04860_ ), .B2(_06234_ ), .ZN(_06395_ ) );
OAI21_X1 _14399_ ( .A(_06393_ ), .B1(_06245_ ), .B2(_06395_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14400_ ( .A(\ID_EX_pc [4] ), .B(_04718_ ), .S(_06233_ ), .Z(_06396_ ) );
NAND3_X1 _14401_ ( .A1(_05752_ ), .A2(_06257_ ), .A3(_05753_ ), .ZN(_06397_ ) );
OAI22_X1 _14402_ ( .A1(_05754_ ), .A2(_04869_ ), .B1(_05433_ ), .B2(\ID_EX_imm [4] ), .ZN(_06398_ ) );
AND3_X1 _14403_ ( .A1(_02861_ ), .A2(_05405_ ), .A3(_02862_ ), .ZN(_06399_ ) );
OAI21_X1 _14404_ ( .A(_06397_ ), .B1(_06398_ ), .B2(_06399_ ), .ZN(_06400_ ) );
MUX2_X1 _14405_ ( .A(_06396_ ), .B(_06400_ ), .S(_06279_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
AND3_X1 _14406_ ( .A1(_05769_ ), .A2(_05770_ ), .A3(_06226_ ), .ZN(_06401_ ) );
NAND2_X1 _14407_ ( .A1(_06401_ ), .A2(_06257_ ), .ZN(_06402_ ) );
AND4_X1 _14408_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06403_ ) );
AOI21_X1 _14409_ ( .A(_06403_ ), .B1(_04695_ ), .B2(_06234_ ), .ZN(_06404_ ) );
OAI221_X1 _14410_ ( .A(_06279_ ), .B1(_05623_ ), .B2(\ID_EX_imm [3] ), .C1(_05771_ ), .C2(_06292_ ), .ZN(_06405_ ) );
AND3_X1 _14411_ ( .A1(_02764_ ), .A2(_05884_ ), .A3(_02765_ ), .ZN(_06406_ ) );
OAI221_X1 _14412_ ( .A(_06402_ ), .B1(_06372_ ), .B2(_06404_ ), .C1(_06405_ ), .C2(_06406_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
NAND3_X1 _14413_ ( .A1(_05335_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_05337_ ), .ZN(_06407_ ) );
AND2_X1 _14414_ ( .A1(_05790_ ), .A2(_06407_ ), .ZN(_06408_ ) );
INV_X1 _14415_ ( .A(_06408_ ), .ZN(_06409_ ) );
OAI22_X1 _14416_ ( .A1(_06409_ ), .A2(_04869_ ), .B1(_05405_ ), .B2(\ID_EX_imm [2] ), .ZN(_06410_ ) );
AOI211_X1 _14417_ ( .A(_06236_ ), .B(_06410_ ), .C1(_05884_ ), .C2(_05047_ ), .ZN(_06411_ ) );
AOI21_X1 _14418_ ( .A(_06227_ ), .B1(_05790_ ), .B2(_05791_ ), .ZN(_06412_ ) );
AND2_X1 _14419_ ( .A1(_06412_ ), .A2(_06257_ ), .ZN(_06413_ ) );
MUX2_X1 _14420_ ( .A(\ID_EX_pc [2] ), .B(_04741_ ), .S(_06232_ ), .Z(_06414_ ) );
AND2_X1 _14421_ ( .A1(_06414_ ), .A2(_06227_ ), .ZN(_06415_ ) );
OR3_X1 _14422_ ( .A1(_06411_ ), .A2(_06413_ ), .A3(_06415_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
NAND4_X1 _14423_ ( .A1(_04039_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06416_ ) );
OAI211_X1 _14424_ ( .A(_06237_ ), .B(_06416_ ), .C1(_04173_ ), .C2(_06231_ ), .ZN(_06417_ ) );
NAND3_X1 _14425_ ( .A1(_05334_ ), .A2(_06256_ ), .A3(_05339_ ), .ZN(_06418_ ) );
OAI21_X1 _14426_ ( .A(_06418_ ), .B1(_05884_ ), .B2(_02200_ ), .ZN(_06419_ ) );
AOI21_X1 _14427_ ( .A(_06419_ ), .B1(_05623_ ), .B2(_02199_ ), .ZN(_06420_ ) );
OAI21_X1 _14428_ ( .A(_06341_ ), .B1(_05340_ ), .B2(_06292_ ), .ZN(_06421_ ) );
OAI21_X1 _14429_ ( .A(_06417_ ), .B1(_06420_ ), .B2(_06421_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
NAND3_X1 _14430_ ( .A1(_05354_ ), .A2(\mepc [1] ), .A3(_05257_ ), .ZN(_06422_ ) );
NAND4_X1 _14431_ ( .A1(_05264_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mtvec [1] ), .ZN(_06423_ ) );
NAND4_X1 _14432_ ( .A1(_05330_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mycsreg.CSReg[0][1] ), .ZN(_06424_ ) );
AND4_X1 _14433_ ( .A1(_06422_ ), .A2(_05800_ ), .A3(_06423_ ), .A4(_06424_ ), .ZN(_06425_ ) );
OR2_X1 _14434_ ( .A1(_05313_ ), .A2(_06425_ ), .ZN(_06426_ ) );
NAND3_X1 _14435_ ( .A1(_05335_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_05337_ ), .ZN(_06427_ ) );
AOI21_X1 _14436_ ( .A(_06262_ ), .B1(_06426_ ), .B2(_06427_ ), .ZN(_06428_ ) );
AND2_X1 _14437_ ( .A1(_06426_ ), .A2(_06427_ ), .ZN(_06429_ ) );
AOI22_X1 _14438_ ( .A1(_06429_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02718_ ), .ZN(_06430_ ) );
NAND3_X1 _14439_ ( .A1(_02715_ ), .A2(_02716_ ), .A3(_05433_ ), .ZN(_06431_ ) );
AOI211_X1 _14440_ ( .A(_06236_ ), .B(_06428_ ), .C1(_06430_ ), .C2(_06431_ ), .ZN(_06432_ ) );
NAND2_X1 _14441_ ( .A1(_04787_ ), .A2(_06234_ ), .ZN(_06433_ ) );
OAI21_X1 _14442_ ( .A(_06433_ ), .B1(\ID_EX_pc [1] ), .B2(_06234_ ), .ZN(_06434_ ) );
AOI21_X1 _14443_ ( .A(_06432_ ), .B1(_06229_ ), .B2(_06434_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
OAI21_X1 _14444_ ( .A(_05833_ ), .B1(_05839_ ), .B2(_05841_ ), .ZN(_06435_ ) );
AOI22_X1 _14445_ ( .A1(_06435_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02720_ ), .ZN(_06436_ ) );
OAI211_X1 _14446_ ( .A(_06436_ ), .B(_06341_ ), .C1(_04743_ ), .C2(\ID_EX_typ [0] ), .ZN(_06437_ ) );
AND3_X1 _14447_ ( .A1(_04762_ ), .A2(_04763_ ), .A3(_06233_ ), .ZN(_06438_ ) );
AND3_X1 _14448_ ( .A1(_03342_ ), .A2(\ID_EX_pc [0] ), .A3(\ID_EX_typ [7] ), .ZN(_06439_ ) );
OAI21_X1 _14449_ ( .A(_06374_ ), .B1(_06438_ ), .B2(_06439_ ), .ZN(_06440_ ) );
OR3_X1 _14450_ ( .A1(_06435_ ), .A2(_06263_ ), .A3(_06236_ ), .ZN(_06441_ ) );
NAND3_X1 _14451_ ( .A1(_06437_ ), .A2(_06440_ ), .A3(_06441_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
NAND4_X1 _14452_ ( .A1(_05607_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06442_ ) );
OAI211_X1 _14453_ ( .A(_06237_ ), .B(_06442_ ), .C1(_04151_ ), .C2(_06231_ ), .ZN(_06443_ ) );
NAND3_X1 _14454_ ( .A1(_05617_ ), .A2(_06256_ ), .A3(_05620_ ), .ZN(_06444_ ) );
INV_X1 _14455_ ( .A(\ID_EX_imm [28] ), .ZN(_06445_ ) );
OAI21_X1 _14456_ ( .A(_06444_ ), .B1(_05884_ ), .B2(_06445_ ), .ZN(_06446_ ) );
AOI21_X1 _14457_ ( .A(_06446_ ), .B1(_05623_ ), .B2(_02226_ ), .ZN(_06447_ ) );
OAI21_X1 _14458_ ( .A(_06341_ ), .B1(_05621_ ), .B2(_06292_ ), .ZN(_06448_ ) );
OAI21_X1 _14459_ ( .A(_06443_ ), .B1(_06447_ ), .B2(_06448_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND4_X1 _14460_ ( .A1(_05331_ ), .A2(_05265_ ), .A3(_05268_ ), .A4(\mycsreg.CSReg[0][27] ), .ZN(_06449_ ) );
NAND4_X1 _14461_ ( .A1(_05326_ ), .A2(_05265_ ), .A3(_05268_ ), .A4(\mtvec [27] ), .ZN(_06450_ ) );
AND4_X1 _14462_ ( .A1(_05819_ ), .A2(_05820_ ), .A3(_06449_ ), .A4(_06450_ ), .ZN(_06451_ ) );
NAND3_X1 _14463_ ( .A1(_05315_ ), .A2(_05319_ ), .A3(_06451_ ), .ZN(_06452_ ) );
OAI211_X1 _14464_ ( .A(_06452_ ), .B(_06256_ ), .C1(\EX_LS_result_csreg_mem [27] ), .C2(_05315_ ), .ZN(_06453_ ) );
OAI21_X1 _14465_ ( .A(_06453_ ), .B1(_05884_ ), .B2(_02249_ ), .ZN(_06454_ ) );
AOI21_X1 _14466_ ( .A(\ID_EX_typ [0] ), .B1(_02246_ ), .B2(_02247_ ), .ZN(_06455_ ) );
OAI221_X1 _14467_ ( .A(_06279_ ), .B1(_06292_ ), .B2(_05826_ ), .C1(_06454_ ), .C2(_06455_ ), .ZN(_06456_ ) );
MUX2_X1 _14468_ ( .A(_05291_ ), .B(_04200_ ), .S(_06238_ ), .Z(_06457_ ) );
OAI21_X1 _14469_ ( .A(_06456_ ), .B1(_06245_ ), .B2(_06457_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
NAND3_X1 _14470_ ( .A1(_05354_ ), .A2(\mepc [26] ), .A3(_05257_ ), .ZN(_06458_ ) );
NAND4_X1 _14471_ ( .A1(_05264_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mtvec [26] ), .ZN(_06459_ ) );
NAND4_X1 _14472_ ( .A1(_05330_ ), .A2(_05356_ ), .A3(_05357_ ), .A4(\mycsreg.CSReg[0][26] ), .ZN(_06460_ ) );
AND4_X1 _14473_ ( .A1(_06458_ ), .A2(_05851_ ), .A3(_06459_ ), .A4(_06460_ ), .ZN(_06461_ ) );
OR2_X1 _14474_ ( .A1(_05313_ ), .A2(_06461_ ), .ZN(_06462_ ) );
NAND3_X1 _14475_ ( .A1(_05335_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_05337_ ), .ZN(_06463_ ) );
AOI21_X1 _14476_ ( .A(_06262_ ), .B1(_06462_ ), .B2(_06463_ ), .ZN(_06464_ ) );
AND2_X1 _14477_ ( .A1(_06462_ ), .A2(_06463_ ), .ZN(_06465_ ) );
AOI22_X1 _14478_ ( .A1(_06465_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02966_ ), .ZN(_06466_ ) );
NAND3_X1 _14479_ ( .A1(_02962_ ), .A2(_02963_ ), .A3(_05433_ ), .ZN(_06467_ ) );
AOI211_X1 _14480_ ( .A(_06236_ ), .B(_06464_ ), .C1(_06466_ ), .C2(_06467_ ), .ZN(_06468_ ) );
MUX2_X1 _14481_ ( .A(_05292_ ), .B(_05179_ ), .S(_06238_ ), .Z(_06469_ ) );
AOI21_X1 _14482_ ( .A(_06468_ ), .B1(_06229_ ), .B2(_06469_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
INV_X1 _14483_ ( .A(_02940_ ), .ZN(_06470_ ) );
NAND3_X1 _14484_ ( .A1(_05241_ ), .A2(\mepc [25] ), .A3(_05258_ ), .ZN(_06471_ ) );
NAND4_X1 _14485_ ( .A1(_05543_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [25] ), .A4(_05265_ ), .ZN(_06472_ ) );
AND4_X1 _14486_ ( .A1(_06471_ ), .A2(_06472_ ), .A3(_05873_ ), .A4(_05874_ ), .ZN(_06473_ ) );
NAND2_X1 _14487_ ( .A1(_06473_ ), .A2(_05745_ ), .ZN(_06474_ ) );
OR3_X1 _14488_ ( .A1(_05534_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_05535_ ), .ZN(_06475_ ) );
NAND2_X1 _14489_ ( .A1(_06474_ ), .A2(_06475_ ), .ZN(_06476_ ) );
AOI22_X1 _14490_ ( .A1(_06470_ ), .A2(_05406_ ), .B1(\ID_EX_typ [2] ), .B2(_06476_ ), .ZN(_06477_ ) );
OAI211_X1 _14491_ ( .A(_06477_ ), .B(_06279_ ), .C1(_05623_ ), .C2(\ID_EX_imm [25] ), .ZN(_06478_ ) );
NAND4_X1 _14492_ ( .A1(_06474_ ), .A2(_06257_ ), .A3(_06475_ ), .A4(_06244_ ), .ZN(_06479_ ) );
MUX2_X1 _14493_ ( .A(_04028_ ), .B(_05176_ ), .S(_06233_ ), .Z(_06480_ ) );
OAI211_X1 _14494_ ( .A(_06478_ ), .B(_06479_ ), .C1(_06245_ ), .C2(_06480_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
AND4_X1 _14495_ ( .A1(\mtvec [24] ), .A2(_05264_ ), .A3(_05261_ ), .A4(_05268_ ), .ZN(_06481_ ) );
NOR2_X1 _14496_ ( .A1(_05892_ ), .A2(_06481_ ), .ZN(_06482_ ) );
NAND3_X1 _14497_ ( .A1(_05321_ ), .A2(\mepc [24] ), .A3(_05389_ ), .ZN(_06483_ ) );
NAND4_X1 _14498_ ( .A1(_05331_ ), .A2(_05444_ ), .A3(_05394_ ), .A4(\mycsreg.CSReg[0][24] ), .ZN(_06484_ ) );
NAND4_X1 _14499_ ( .A1(_06482_ ), .A2(_05513_ ), .A3(_06483_ ), .A4(_06484_ ), .ZN(_06485_ ) );
NAND2_X1 _14500_ ( .A1(_05315_ ), .A2(_06485_ ), .ZN(_06486_ ) );
NAND3_X1 _14501_ ( .A1(_05427_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_05428_ ), .ZN(_06487_ ) );
NAND2_X1 _14502_ ( .A1(_06486_ ), .A2(_06487_ ), .ZN(_06488_ ) );
AND2_X1 _14503_ ( .A1(_06486_ ), .A2(_06487_ ), .ZN(_06489_ ) );
OAI22_X1 _14504_ ( .A1(_06489_ ), .A2(_06263_ ), .B1(_05884_ ), .B2(_02272_ ), .ZN(_06490_ ) );
AOI21_X1 _14505_ ( .A(\ID_EX_typ [0] ), .B1(_02269_ ), .B2(_02270_ ), .ZN(_06491_ ) );
OAI221_X1 _14506_ ( .A(_06372_ ), .B1(_06292_ ), .B2(_06488_ ), .C1(_06490_ ), .C2(_06491_ ), .ZN(_06492_ ) );
NAND4_X1 _14507_ ( .A1(_05865_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06493_ ) );
OAI211_X1 _14508_ ( .A(_06374_ ), .B(_06493_ ), .C1(_04270_ ), .C2(_06231_ ), .ZN(_06494_ ) );
NAND2_X1 _14509_ ( .A1(_06492_ ), .A2(_06494_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
AOI22_X1 _14510_ ( .A1(_05922_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02308_ ), .ZN(_06495_ ) );
OAI211_X1 _14511_ ( .A(_06495_ ), .B(_06279_ ), .C1(_02307_ ), .C2(\ID_EX_typ [0] ), .ZN(_06496_ ) );
AND3_X1 _14512_ ( .A1(_05920_ ), .A2(_05921_ ), .A3(_06226_ ), .ZN(_06497_ ) );
NAND2_X1 _14513_ ( .A1(_06497_ ), .A2(_06257_ ), .ZN(_06498_ ) );
MUX2_X1 _14514_ ( .A(_04008_ ), .B(_04405_ ), .S(_06233_ ), .Z(_06499_ ) );
OAI211_X1 _14515_ ( .A(_06496_ ), .B(_06498_ ), .C1(_06245_ ), .C2(_06499_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
AOI22_X1 _14516_ ( .A1(_05940_ ), .A2(_06256_ ), .B1(\ID_EX_typ [0] ), .B2(\ID_EX_imm [22] ), .ZN(_06500_ ) );
INV_X1 _14517_ ( .A(_02333_ ), .ZN(_06501_ ) );
OAI21_X1 _14518_ ( .A(_06500_ ), .B1(\ID_EX_typ [0] ), .B2(_06501_ ), .ZN(_06502_ ) );
OAI211_X1 _14519_ ( .A(_06502_ ), .B(_06372_ ), .C1(_06292_ ), .C2(_05940_ ), .ZN(_06503_ ) );
OR4_X1 _14520_ ( .A1(\ID_EX_pc [22] ), .A2(_03343_ ), .A3(_03898_ ), .A4(_03889_ ), .ZN(_06504_ ) );
OAI211_X1 _14521_ ( .A(_06374_ ), .B(_06504_ ), .C1(_04429_ ), .C2(_06231_ ), .ZN(_06505_ ) );
NAND2_X1 _14522_ ( .A1(_06503_ ), .A2(_06505_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14523_ ( .A(\ID_EX_pc [31] ), .B(_04127_ ), .S(_06233_ ), .Z(_06506_ ) );
NOR2_X1 _14524_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06507_ ) );
INV_X1 _14525_ ( .A(_06507_ ), .ZN(_06508_ ) );
MUX2_X1 _14526_ ( .A(_04883_ ), .B(_04878_ ), .S(_03886_ ), .Z(_06509_ ) );
NOR3_X1 _14527_ ( .A1(_06509_ ), .A2(_05981_ ), .A3(_05982_ ), .ZN(_06510_ ) );
NAND2_X1 _14528_ ( .A1(_06510_ ), .A2(_06262_ ), .ZN(_06511_ ) );
INV_X1 _14529_ ( .A(_06511_ ), .ZN(_06512_ ) );
OR2_X1 _14530_ ( .A1(_05981_ ), .A2(_05982_ ), .ZN(_06513_ ) );
AOI21_X1 _14531_ ( .A(_06262_ ), .B1(_06509_ ), .B2(_06513_ ), .ZN(_06514_ ) );
OAI21_X1 _14532_ ( .A(_06508_ ), .B1(_06512_ ), .B2(_06514_ ), .ZN(_06515_ ) );
OAI21_X1 _14533_ ( .A(_06515_ ), .B1(_06508_ ), .B2(_06509_ ), .ZN(_06516_ ) );
MUX2_X1 _14534_ ( .A(_06506_ ), .B(_06516_ ), .S(_06244_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
NAND3_X1 _14535_ ( .A1(_05958_ ), .A2(_05960_ ), .A3(_06341_ ), .ZN(_06517_ ) );
BUF_X4 _14536_ ( .A(_05206_ ), .Z(_06518_ ) );
NOR3_X1 _14537_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_06519_ ) );
AND2_X1 _14538_ ( .A1(\ID_EX_typ [3] ), .A2(\ID_EX_typ [2] ), .ZN(_06520_ ) );
AND2_X1 _14539_ ( .A1(_06519_ ), .A2(_06520_ ), .ZN(_06521_ ) );
INV_X1 _14540_ ( .A(_06521_ ), .ZN(_06522_ ) );
BUF_X2 _14541_ ( .A(_06522_ ), .Z(_06523_ ) );
NOR3_X1 _14542_ ( .A1(_04867_ ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_06524_ ) );
AND2_X1 _14543_ ( .A1(_06524_ ), .A2(_06520_ ), .ZN(_06525_ ) );
INV_X1 _14544_ ( .A(_06525_ ), .ZN(_06526_ ) );
BUF_X4 _14545_ ( .A(_06526_ ), .Z(_06527_ ) );
OAI22_X1 _14546_ ( .A1(_05950_ ), .A2(_06523_ ), .B1(_02357_ ), .B2(_06527_ ), .ZN(_06528_ ) );
NAND2_X1 _14547_ ( .A1(_05150_ ), .A2(_04381_ ), .ZN(_06529_ ) );
AND2_X1 _14548_ ( .A1(_06529_ ), .A2(_05159_ ), .ZN(_06530_ ) );
INV_X1 _14549_ ( .A(_04454_ ), .ZN(_06531_ ) );
NOR2_X1 _14550_ ( .A1(_06530_ ), .A2(_06531_ ), .ZN(_06532_ ) );
NOR2_X1 _14551_ ( .A1(_06532_ ), .A2(_05167_ ), .ZN(_06533_ ) );
XNOR2_X1 _14552_ ( .A(_06533_ ), .B(_04480_ ), .ZN(_06534_ ) );
AND3_X1 _14553_ ( .A1(_04045_ ), .A2(\ID_EX_typ [3] ), .A3(_04869_ ), .ZN(_06535_ ) );
AND2_X1 _14554_ ( .A1(_06535_ ), .A2(_04881_ ), .ZN(_06536_ ) );
BUF_X4 _14555_ ( .A(_06536_ ), .Z(_06537_ ) );
AOI21_X1 _14556_ ( .A(_06528_ ), .B1(_06534_ ), .B2(_06537_ ), .ZN(_06538_ ) );
NOR2_X1 _14557_ ( .A1(_03889_ ), .A2(\ID_EX_typ [6] ), .ZN(_06539_ ) );
AND2_X2 _14558_ ( .A1(_06539_ ), .A2(_03343_ ), .ZN(_06540_ ) );
INV_X2 _14559_ ( .A(_06540_ ), .ZN(_06541_ ) );
BUF_X4 _14560_ ( .A(_06541_ ), .Z(_06542_ ) );
BUF_X4 _14561_ ( .A(_06542_ ), .Z(_06543_ ) );
OAI21_X1 _14562_ ( .A(_06518_ ), .B1(_06538_ ), .B2(_06543_ ), .ZN(_06544_ ) );
INV_X1 _14563_ ( .A(_04955_ ), .ZN(_06545_ ) );
AND2_X1 _14564_ ( .A1(_04995_ ), .A2(_04999_ ), .ZN(_06546_ ) );
INV_X1 _14565_ ( .A(_06546_ ), .ZN(_06547_ ) );
AND2_X1 _14566_ ( .A1(_05033_ ), .A2(_02766_ ), .ZN(_06548_ ) );
INV_X1 _14567_ ( .A(_06548_ ), .ZN(_06549_ ) );
NOR2_X1 _14568_ ( .A1(_05028_ ), .A2(_05047_ ), .ZN(_06550_ ) );
INV_X1 _14569_ ( .A(_06550_ ), .ZN(_06551_ ) );
INV_X1 _14570_ ( .A(_04743_ ), .ZN(_06552_ ) );
NOR2_X1 _14571_ ( .A1(_05044_ ), .A2(_06552_ ), .ZN(_06553_ ) );
INV_X1 _14572_ ( .A(_06553_ ), .ZN(_06554_ ) );
NOR3_X2 _14573_ ( .A1(_06554_ ), .A2(_05041_ ), .A3(_05039_ ), .ZN(_06555_ ) );
NOR2_X1 _14574_ ( .A1(_06555_ ), .A2(_05041_ ), .ZN(_06556_ ) );
INV_X1 _14575_ ( .A(_05029_ ), .ZN(_06557_ ) );
OAI211_X4 _14576_ ( .A(_06549_ ), .B(_06551_ ), .C1(_06556_ ), .C2(_06557_ ), .ZN(_06558_ ) );
NOR2_X1 _14577_ ( .A1(_05033_ ), .A2(_02766_ ), .ZN(_06559_ ) );
INV_X1 _14578_ ( .A(_06559_ ), .ZN(_06560_ ) );
AND2_X1 _14579_ ( .A1(_05004_ ), .A2(_05009_ ), .ZN(_06561_ ) );
AND2_X1 _14580_ ( .A1(_05019_ ), .A2(_05052_ ), .ZN(_06562_ ) );
NAND4_X1 _14581_ ( .A1(_06558_ ), .A2(_06560_ ), .A3(_06561_ ), .A4(_06562_ ), .ZN(_06563_ ) );
NOR2_X1 _14582_ ( .A1(_05003_ ), .A2(_06370_ ), .ZN(_06564_ ) );
NOR2_X1 _14583_ ( .A1(_05008_ ), .A2(_02870_ ), .ZN(_06565_ ) );
NOR2_X1 _14584_ ( .A1(_05018_ ), .A2(_02841_ ), .ZN(_06566_ ) );
AND2_X1 _14585_ ( .A1(_05018_ ), .A2(_02841_ ), .ZN(_06567_ ) );
INV_X1 _14586_ ( .A(_06567_ ), .ZN(_06568_ ) );
AND2_X1 _14587_ ( .A1(_05014_ ), .A2(_02863_ ), .ZN(_06569_ ) );
INV_X1 _14588_ ( .A(_06569_ ), .ZN(_06570_ ) );
AOI21_X1 _14589_ ( .A(_06566_ ), .B1(_06568_ ), .B2(_06570_ ), .ZN(_06571_ ) );
AOI221_X2 _14590_ ( .A(_06564_ ), .B1(_05004_ ), .B2(_06565_ ), .C1(_06571_ ), .C2(_06561_ ), .ZN(_06572_ ) );
AOI21_X2 _14591_ ( .A(_06547_ ), .B1(_06563_ ), .B2(_06572_ ), .ZN(_06573_ ) );
AND3_X1 _14592_ ( .A1(_04967_ ), .A2(_04968_ ), .A3(_04962_ ), .ZN(_06574_ ) );
AND2_X1 _14593_ ( .A1(_04973_ ), .A2(_04978_ ), .ZN(_06575_ ) );
AND2_X1 _14594_ ( .A1(_04984_ ), .A2(_04989_ ), .ZN(_06576_ ) );
NAND4_X1 _14595_ ( .A1(_06573_ ), .A2(_06574_ ), .A3(_06575_ ), .A4(_06576_ ), .ZN(_06577_ ) );
INV_X1 _14596_ ( .A(_05063_ ), .ZN(_06578_ ) );
INV_X1 _14597_ ( .A(_02599_ ), .ZN(_06579_ ) );
NOR2_X1 _14598_ ( .A1(_04998_ ), .A2(_06579_ ), .ZN(_06580_ ) );
AOI21_X1 _14599_ ( .A(_05064_ ), .B1(_06578_ ), .B2(_06580_ ), .ZN(_06581_ ) );
NOR3_X1 _14600_ ( .A1(_06581_ ), .A2(_04985_ ), .A3(_04990_ ), .ZN(_06582_ ) );
NOR2_X1 _14601_ ( .A1(_04983_ ), .A2(_05068_ ), .ZN(_06583_ ) );
INV_X1 _14602_ ( .A(_02647_ ), .ZN(_06584_ ) );
NOR2_X1 _14603_ ( .A1(_04988_ ), .A2(_06584_ ), .ZN(_06585_ ) );
AND2_X1 _14604_ ( .A1(_04984_ ), .A2(_06585_ ), .ZN(_06586_ ) );
NOR3_X2 _14605_ ( .A1(_06582_ ), .A2(_06583_ ), .A3(_06586_ ), .ZN(_06587_ ) );
NAND3_X1 _14606_ ( .A1(_05056_ ), .A2(_04962_ ), .A3(_06575_ ), .ZN(_06588_ ) );
OR2_X1 _14607_ ( .A1(_06587_ ), .A2(_06588_ ), .ZN(_06589_ ) );
NOR2_X1 _14608_ ( .A1(_04961_ ), .A2(_05057_ ), .ZN(_06590_ ) );
NAND3_X1 _14609_ ( .A1(_04967_ ), .A2(_04968_ ), .A3(_06590_ ), .ZN(_06591_ ) );
INV_X1 _14610_ ( .A(_02552_ ), .ZN(_06592_ ) );
NOR2_X1 _14611_ ( .A1(_04972_ ), .A2(_06592_ ), .ZN(_06593_ ) );
NOR2_X1 _14612_ ( .A1(_04977_ ), .A2(_05072_ ), .ZN(_06594_ ) );
AOI21_X1 _14613_ ( .A(_06593_ ), .B1(_04973_ ), .B2(_06594_ ), .ZN(_06595_ ) );
INV_X1 _14614_ ( .A(_06595_ ), .ZN(_06596_ ) );
NAND3_X1 _14615_ ( .A1(_05056_ ), .A2(_04962_ ), .A3(_06596_ ), .ZN(_06597_ ) );
AND4_X2 _14616_ ( .A1(_04967_ ), .A2(_06589_ ), .A3(_06591_ ), .A4(_06597_ ), .ZN(_06598_ ) );
AND2_X1 _14617_ ( .A1(_06577_ ), .A2(_06598_ ), .ZN(_06599_ ) );
INV_X1 _14618_ ( .A(_06599_ ), .ZN(_06600_ ) );
AND2_X1 _14619_ ( .A1(_05080_ ), .A2(_05081_ ), .ZN(_06601_ ) );
NAND4_X2 _14620_ ( .A1(_06600_ ), .A2(_04943_ ), .A3(_04948_ ), .A4(_06601_ ), .ZN(_06602_ ) );
INV_X1 _14621_ ( .A(_02480_ ), .ZN(_06603_ ) );
NOR2_X1 _14622_ ( .A1(_04930_ ), .A2(_06603_ ), .ZN(_06604_ ) );
AOI21_X1 _14623_ ( .A(_04936_ ), .B1(_05080_ ), .B2(_06604_ ), .ZN(_06605_ ) );
NOR3_X1 _14624_ ( .A1(_06605_ ), .A2(_04944_ ), .A3(_04949_ ), .ZN(_06606_ ) );
NOR2_X1 _14625_ ( .A1(_04942_ ), .A2(_04952_ ), .ZN(_06607_ ) );
INV_X1 _14626_ ( .A(_02406_ ), .ZN(_06608_ ) );
NOR2_X1 _14627_ ( .A1(_04947_ ), .A2(_06608_ ), .ZN(_06609_ ) );
AND2_X1 _14628_ ( .A1(_04943_ ), .A2(_06609_ ), .ZN(_06610_ ) );
NOR3_X1 _14629_ ( .A1(_06606_ ), .A2(_06607_ ), .A3(_06610_ ), .ZN(_06611_ ) );
AOI21_X1 _14630_ ( .A(_06545_ ), .B1(_06602_ ), .B2(_06611_ ), .ZN(_06612_ ) );
INV_X1 _14631_ ( .A(_02382_ ), .ZN(_06613_ ) );
NOR2_X1 _14632_ ( .A1(_04918_ ), .A2(_06613_ ), .ZN(_06614_ ) );
OR3_X1 _14633_ ( .A1(_06612_ ), .A2(_06614_ ), .A3(_04956_ ), .ZN(_06615_ ) );
NOR2_X1 _14634_ ( .A1(_04866_ ), .A2(_06508_ ), .ZN(_06616_ ) );
BUF_X2 _14635_ ( .A(_06616_ ), .Z(_06617_ ) );
OAI21_X1 _14636_ ( .A(_04956_ ), .B1(_06612_ ), .B2(_06614_ ), .ZN(_06618_ ) );
NAND3_X1 _14637_ ( .A1(_06615_ ), .A2(_06617_ ), .A3(_06618_ ), .ZN(_06619_ ) );
AND2_X2 _14638_ ( .A1(_05193_ ), .A2(\ID_EX_typ [2] ), .ZN(_06620_ ) );
BUF_X4 _14639_ ( .A(_06620_ ), .Z(_06621_ ) );
AND2_X1 _14640_ ( .A1(_05044_ ), .A2(_05040_ ), .ZN(_06622_ ) );
AND2_X2 _14641_ ( .A1(_06622_ ), .A2(_05028_ ), .ZN(_06623_ ) );
INV_X1 _14642_ ( .A(_05033_ ), .ZN(_06624_ ) );
BUF_X4 _14643_ ( .A(_06624_ ), .Z(_06625_ ) );
AND2_X1 _14644_ ( .A1(_06623_ ), .A2(_06625_ ), .ZN(_06626_ ) );
BUF_X2 _14645_ ( .A(_05013_ ), .Z(_06627_ ) );
AND2_X2 _14646_ ( .A1(_06626_ ), .A2(_06627_ ), .ZN(_06628_ ) );
INV_X1 _14647_ ( .A(_06628_ ), .ZN(_06629_ ) );
NOR4_X1 _14648_ ( .A1(_04965_ ), .A2(_04961_ ), .A3(_04933_ ), .A4(_04930_ ), .ZN(_06630_ ) );
INV_X1 _14649_ ( .A(_04972_ ), .ZN(_06631_ ) );
INV_X1 _14650_ ( .A(_04988_ ), .ZN(_06632_ ) );
AOI22_X1 _14651_ ( .A1(_04997_ ), .A2(_04996_ ), .B1(_05001_ ), .B2(_05002_ ), .ZN(_06633_ ) );
AOI22_X1 _14652_ ( .A1(_04993_ ), .A2(_04992_ ), .B1(_05006_ ), .B2(_05007_ ), .ZN(_06634_ ) );
AND4_X1 _14653_ ( .A1(_06631_ ), .A2(_06632_ ), .A3(_06633_ ), .A4(_06634_ ), .ZN(_06635_ ) );
AND4_X1 _14654_ ( .A1(_05073_ ), .A2(_06630_ ), .A3(_05069_ ), .A4(_06635_ ), .ZN(_06636_ ) );
NOR4_X1 _14655_ ( .A1(_04921_ ), .A2(_04918_ ), .A3(_04942_ ), .A4(_04947_ ), .ZN(_06637_ ) );
NAND4_X1 _14656_ ( .A1(_06629_ ), .A2(_06636_ ), .A3(_05018_ ), .A4(_06637_ ), .ZN(_06638_ ) );
AND4_X1 _14657_ ( .A1(_05003_ ), .A2(_05018_ ), .A3(_05008_ ), .A4(_06627_ ), .ZN(_06639_ ) );
NAND3_X1 _14658_ ( .A1(_06623_ ), .A2(_06639_ ), .A3(_06624_ ), .ZN(_06640_ ) );
NAND4_X1 _14659_ ( .A1(_05003_ ), .A2(_05016_ ), .A3(_05008_ ), .A4(_05017_ ), .ZN(_06641_ ) );
NAND2_X1 _14660_ ( .A1(_06640_ ), .A2(_06641_ ), .ZN(_06642_ ) );
NAND4_X1 _14661_ ( .A1(_04965_ ), .A2(_04972_ ), .A3(_04961_ ), .A4(_04977_ ), .ZN(_06643_ ) );
NAND2_X1 _14662_ ( .A1(_04998_ ), .A2(_04994_ ), .ZN(_06644_ ) );
OR3_X1 _14663_ ( .A1(_06644_ ), .A2(_05069_ ), .A3(_06632_ ), .ZN(_06645_ ) );
NOR2_X1 _14664_ ( .A1(_06643_ ), .A2(_06645_ ), .ZN(_06646_ ) );
AND2_X1 _14665_ ( .A1(_04921_ ), .A2(_04918_ ), .ZN(_06647_ ) );
AND2_X1 _14666_ ( .A1(_04933_ ), .A2(_04930_ ), .ZN(_06648_ ) );
AND4_X1 _14667_ ( .A1(_04942_ ), .A2(_06647_ ), .A3(_04947_ ), .A4(_06648_ ), .ZN(_06649_ ) );
AND3_X1 _14668_ ( .A1(_06642_ ), .A2(_06646_ ), .A3(_06649_ ), .ZN(_06650_ ) );
INV_X1 _14669_ ( .A(_06650_ ), .ZN(_06651_ ) );
OR3_X1 _14670_ ( .A1(_06650_ ), .A2(_04905_ ), .A3(_04911_ ), .ZN(_06652_ ) );
AND2_X1 _14671_ ( .A1(_04911_ ), .A2(_04905_ ), .ZN(_06653_ ) );
NAND2_X1 _14672_ ( .A1(_06650_ ), .A2(_06653_ ), .ZN(_06654_ ) );
AOI221_X4 _14673_ ( .A(_04878_ ), .B1(_06638_ ), .B2(_06651_ ), .C1(_06652_ ), .C2(_06654_ ), .ZN(_06655_ ) );
INV_X1 _14674_ ( .A(_04893_ ), .ZN(_06656_ ) );
NAND4_X1 _14675_ ( .A1(_05116_ ), .A2(_05096_ ), .A3(_05101_ ), .A4(_06656_ ), .ZN(_06657_ ) );
NAND3_X1 _14676_ ( .A1(_05087_ ), .A2(_05091_ ), .A3(_04885_ ), .ZN(_06658_ ) );
NOR3_X1 _14677_ ( .A1(_06657_ ), .A2(_04876_ ), .A3(_06658_ ), .ZN(_06659_ ) );
NAND3_X1 _14678_ ( .A1(_06650_ ), .A2(_06653_ ), .A3(_06659_ ), .ZN(_06660_ ) );
NOR4_X1 _14679_ ( .A1(_05116_ ), .A2(_05096_ ), .A3(_05101_ ), .A4(_06656_ ), .ZN(_06661_ ) );
NAND4_X1 _14680_ ( .A1(_06661_ ), .A2(_05085_ ), .A3(_05086_ ), .A4(_04876_ ), .ZN(_06662_ ) );
OR3_X1 _14681_ ( .A1(_06662_ ), .A2(_05091_ ), .A3(_04885_ ), .ZN(_06663_ ) );
AND2_X1 _14682_ ( .A1(_06650_ ), .A2(_06653_ ), .ZN(_06664_ ) );
OAI21_X1 _14683_ ( .A(_06660_ ), .B1(_06663_ ), .B2(_06664_ ), .ZN(_06665_ ) );
AND2_X2 _14684_ ( .A1(_06655_ ), .A2(_06665_ ), .ZN(_06666_ ) );
XNOR2_X1 _14685_ ( .A(_06628_ ), .B(_05018_ ), .ZN(_06667_ ) );
NAND2_X1 _14686_ ( .A1(_06666_ ), .A2(_06667_ ), .ZN(_06668_ ) );
XNOR2_X1 _14687_ ( .A(_06626_ ), .B(_06627_ ), .ZN(_06669_ ) );
NOR2_X1 _14688_ ( .A1(_06669_ ), .A2(_05018_ ), .ZN(_06670_ ) );
INV_X1 _14689_ ( .A(_06670_ ), .ZN(_06671_ ) );
AND2_X1 _14690_ ( .A1(_06668_ ), .A2(_06671_ ), .ZN(_06672_ ) );
BUF_X4 _14691_ ( .A(_05048_ ), .Z(_06673_ ) );
XNOR2_X1 _14692_ ( .A(_06622_ ), .B(_06673_ ), .ZN(_06674_ ) );
INV_X1 _14693_ ( .A(_06674_ ), .ZN(_06675_ ) );
NAND2_X1 _14694_ ( .A1(_06666_ ), .A2(_06675_ ), .ZN(_06676_ ) );
BUF_X2 _14695_ ( .A(_06665_ ), .Z(_06677_ ) );
BUF_X4 _14696_ ( .A(_05044_ ), .Z(_06678_ ) );
BUF_X4 _14697_ ( .A(_06678_ ), .Z(_06679_ ) );
BUF_X4 _14698_ ( .A(_06679_ ), .Z(_06680_ ) );
BUF_X4 _14699_ ( .A(_05040_ ), .Z(_06681_ ) );
BUF_X4 _14700_ ( .A(_06681_ ), .Z(_06682_ ) );
BUF_X4 _14701_ ( .A(_06682_ ), .Z(_06683_ ) );
XNOR2_X1 _14702_ ( .A(_06680_ ), .B(_06683_ ), .ZN(_06684_ ) );
NAND3_X1 _14703_ ( .A1(_06655_ ), .A2(_06677_ ), .A3(_06684_ ), .ZN(_06685_ ) );
NAND2_X1 _14704_ ( .A1(_06676_ ), .A2(_06685_ ), .ZN(_06686_ ) );
XNOR2_X1 _14705_ ( .A(_06623_ ), .B(_05033_ ), .ZN(_06687_ ) );
INV_X1 _14706_ ( .A(_06687_ ), .ZN(_06688_ ) );
BUF_X2 _14707_ ( .A(_06688_ ), .Z(_06689_ ) );
NAND2_X1 _14708_ ( .A1(_06686_ ), .A2(_06689_ ), .ZN(_06690_ ) );
INV_X1 _14709_ ( .A(_06669_ ), .ZN(_06691_ ) );
AOI21_X1 _14710_ ( .A(_06672_ ), .B1(_06690_ ), .B2(_06691_ ), .ZN(_06692_ ) );
BUF_X4 _14711_ ( .A(_06673_ ), .Z(_06693_ ) );
INV_X1 _14712_ ( .A(_05044_ ), .ZN(_06694_ ) );
NAND3_X1 _14713_ ( .A1(_02160_ ), .A2(_06694_ ), .A3(_02171_ ), .ZN(_06695_ ) );
NAND2_X1 _14714_ ( .A1(_06679_ ), .A2(_04894_ ), .ZN(_06696_ ) );
NAND3_X1 _14715_ ( .A1(_06695_ ), .A2(_06683_ ), .A3(_06696_ ), .ZN(_06697_ ) );
INV_X2 _14716_ ( .A(_05040_ ), .ZN(_06698_ ) );
BUF_X4 _14717_ ( .A(_06698_ ), .Z(_06699_ ) );
BUF_X4 _14718_ ( .A(_06699_ ), .Z(_06700_ ) );
NAND3_X1 _14719_ ( .A1(_06700_ ), .A2(_03005_ ), .A3(_06680_ ), .ZN(_06701_ ) );
AOI21_X1 _14720_ ( .A(_06693_ ), .B1(_06697_ ), .B2(_06701_ ), .ZN(_06702_ ) );
BUF_X2 _14721_ ( .A(_05048_ ), .Z(_06703_ ) );
BUF_X4 _14722_ ( .A(_05042_ ), .Z(_06704_ ) );
BUF_X4 _14723_ ( .A(_06704_ ), .Z(_06705_ ) );
BUF_X4 _14724_ ( .A(_05043_ ), .Z(_06706_ ) );
BUF_X4 _14725_ ( .A(_06706_ ), .Z(_06707_ ) );
AOI21_X1 _14726_ ( .A(_02248_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06708_ ) );
AOI211_X1 _14727_ ( .A(_06681_ ), .B(_06708_ ), .C1(_02976_ ), .C2(_06694_ ), .ZN(_06709_ ) );
BUF_X4 _14728_ ( .A(_05044_ ), .Z(_06710_ ) );
NOR2_X1 _14729_ ( .A1(_06710_ ), .A2(_02965_ ), .ZN(_06711_ ) );
AOI21_X1 _14730_ ( .A(_02940_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06712_ ) );
NOR3_X1 _14731_ ( .A1(_06711_ ), .A2(_06699_ ), .A3(_06712_ ), .ZN(_06713_ ) );
OAI21_X1 _14732_ ( .A(_06703_ ), .B1(_06709_ ), .B2(_06713_ ), .ZN(_06714_ ) );
BUF_X2 _14733_ ( .A(_06682_ ), .Z(_06715_ ) );
NOR2_X1 _14734_ ( .A1(_06679_ ), .A2(_02333_ ), .ZN(_06716_ ) );
AOI21_X1 _14735_ ( .A(_04477_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06717_ ) );
OAI21_X1 _14736_ ( .A(_06715_ ), .B1(_06716_ ), .B2(_06717_ ), .ZN(_06718_ ) );
BUF_X4 _14737_ ( .A(_06699_ ), .Z(_06719_ ) );
NOR2_X1 _14738_ ( .A1(_06679_ ), .A2(_02271_ ), .ZN(_06720_ ) );
AOI21_X1 _14739_ ( .A(_02307_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06721_ ) );
OAI21_X1 _14740_ ( .A(_06719_ ), .B1(_06720_ ), .B2(_06721_ ), .ZN(_06722_ ) );
BUF_X4 _14741_ ( .A(_05028_ ), .Z(_06723_ ) );
BUF_X4 _14742_ ( .A(_06723_ ), .Z(_06724_ ) );
NAND3_X1 _14743_ ( .A1(_06718_ ), .A2(_06722_ ), .A3(_06724_ ), .ZN(_06725_ ) );
NAND2_X1 _14744_ ( .A1(_06714_ ), .A2(_06725_ ), .ZN(_06726_ ) );
BUF_X4 _14745_ ( .A(_06625_ ), .Z(_06727_ ) );
MUX2_X1 _14746_ ( .A(_06702_ ), .B(_06726_ ), .S(_06727_ ), .Z(_06728_ ) );
BUF_X2 _14747_ ( .A(_06627_ ), .Z(_06729_ ) );
BUF_X2 _14748_ ( .A(_06729_ ), .Z(_06730_ ) );
BUF_X2 _14749_ ( .A(_06730_ ), .Z(_06731_ ) );
AND2_X1 _14750_ ( .A1(_06728_ ), .A2(_06731_ ), .ZN(_06732_ ) );
OAI21_X1 _14751_ ( .A(_06621_ ), .B1(_06692_ ), .B2(_06732_ ), .ZN(_06733_ ) );
BUF_X2 _14752_ ( .A(_06627_ ), .Z(_06734_ ) );
BUF_X2 _14753_ ( .A(_06734_ ), .Z(_06735_ ) );
AND2_X1 _14754_ ( .A1(_04868_ ), .A2(\ID_EX_typ [2] ), .ZN(_06736_ ) );
BUF_X2 _14755_ ( .A(_06736_ ), .Z(_06737_ ) );
AND3_X1 _14756_ ( .A1(_06728_ ), .A2(_06735_ ), .A3(_06737_ ), .ZN(_06738_ ) );
BUF_X2 _14757_ ( .A(_05191_ ), .Z(_06739_ ) );
INV_X1 _14758_ ( .A(_06739_ ), .ZN(_06740_ ) );
BUF_X2 _14759_ ( .A(_06724_ ), .Z(_06741_ ) );
NOR2_X1 _14760_ ( .A1(_06710_ ), .A2(_02526_ ), .ZN(_06742_ ) );
BUF_X4 _14761_ ( .A(_05042_ ), .Z(_06743_ ) );
BUF_X4 _14762_ ( .A(_05043_ ), .Z(_06744_ ) );
AOI21_X1 _14763_ ( .A(_02503_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06745_ ) );
BUF_X4 _14764_ ( .A(_06681_ ), .Z(_06746_ ) );
BUF_X4 _14765_ ( .A(_06746_ ), .Z(_06747_ ) );
OR3_X1 _14766_ ( .A1(_06742_ ), .A2(_06745_ ), .A3(_06747_ ), .ZN(_06748_ ) );
NOR2_X1 _14767_ ( .A1(_06678_ ), .A2(_02480_ ), .ZN(_06749_ ) );
BUF_X4 _14768_ ( .A(_06698_ ), .Z(_06750_ ) );
BUF_X2 _14769_ ( .A(_06750_ ), .Z(_06751_ ) );
AOI21_X1 _14770_ ( .A(_02458_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06752_ ) );
OR3_X1 _14771_ ( .A1(_06749_ ), .A2(_06751_ ), .A3(_06752_ ), .ZN(_06753_ ) );
AOI21_X1 _14772_ ( .A(_06741_ ), .B1(_06748_ ), .B2(_06753_ ), .ZN(_06754_ ) );
NOR2_X1 _14773_ ( .A1(_06679_ ), .A2(_02382_ ), .ZN(_06755_ ) );
OAI21_X1 _14774_ ( .A(_06747_ ), .B1(_06755_ ), .B2(_06717_ ), .ZN(_06756_ ) );
NOR2_X1 _14775_ ( .A1(_06678_ ), .A2(_02406_ ), .ZN(_06757_ ) );
AOI21_X1 _14776_ ( .A(_04330_ ), .B1(_06704_ ), .B2(_06706_ ), .ZN(_06758_ ) );
OAI21_X1 _14777_ ( .A(_06751_ ), .B1(_06757_ ), .B2(_06758_ ), .ZN(_06759_ ) );
BUF_X2 _14778_ ( .A(_06723_ ), .Z(_06760_ ) );
AND3_X1 _14779_ ( .A1(_06756_ ), .A2(_06759_ ), .A3(_06760_ ), .ZN(_06761_ ) );
BUF_X4 _14780_ ( .A(_05033_ ), .Z(_06762_ ) );
BUF_X4 _14781_ ( .A(_06762_ ), .Z(_06763_ ) );
OR3_X1 _14782_ ( .A1(_06754_ ), .A2(_06761_ ), .A3(_06763_ ), .ZN(_06764_ ) );
BUF_X2 _14783_ ( .A(_06734_ ), .Z(_06765_ ) );
BUF_X4 _14784_ ( .A(_06762_ ), .Z(_06766_ ) );
BUF_X4 _14785_ ( .A(_06766_ ), .Z(_06767_ ) );
NOR2_X1 _14786_ ( .A1(_06678_ ), .A2(_02647_ ), .ZN(_06768_ ) );
AOI21_X1 _14787_ ( .A(_02670_ ), .B1(_06704_ ), .B2(_06706_ ), .ZN(_06769_ ) );
OR3_X1 _14788_ ( .A1(_06768_ ), .A2(_06715_ ), .A3(_06769_ ), .ZN(_06770_ ) );
NOR2_X1 _14789_ ( .A1(_06710_ ), .A2(_02574_ ), .ZN(_06771_ ) );
AOI21_X1 _14790_ ( .A(_02552_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06772_ ) );
OR3_X1 _14791_ ( .A1(_06771_ ), .A2(_06719_ ), .A3(_06772_ ), .ZN(_06773_ ) );
AND3_X1 _14792_ ( .A1(_06770_ ), .A2(_06773_ ), .A3(_06760_ ), .ZN(_06774_ ) );
NOR2_X1 _14793_ ( .A1(_06678_ ), .A2(_02600_ ), .ZN(_06775_ ) );
AOI21_X1 _14794_ ( .A(_02624_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06776_ ) );
OAI21_X1 _14795_ ( .A(_06747_ ), .B1(_06775_ ), .B2(_06776_ ), .ZN(_06777_ ) );
NOR2_X1 _14796_ ( .A1(_05044_ ), .A2(_02792_ ), .ZN(_06778_ ) );
AOI21_X1 _14797_ ( .A(_02816_ ), .B1(_06704_ ), .B2(_06706_ ), .ZN(_06779_ ) );
OAI21_X1 _14798_ ( .A(_06751_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06780_ ) );
AOI21_X1 _14799_ ( .A(_06760_ ), .B1(_06777_ ), .B2(_06780_ ), .ZN(_06781_ ) );
OAI21_X1 _14800_ ( .A(_06767_ ), .B1(_06774_ ), .B2(_06781_ ), .ZN(_06782_ ) );
NAND3_X1 _14801_ ( .A1(_06764_ ), .A2(_06765_ ), .A3(_06782_ ), .ZN(_06783_ ) );
AOI21_X1 _14802_ ( .A(_02841_ ), .B1(_06704_ ), .B2(_06706_ ), .ZN(_06784_ ) );
NOR2_X1 _14803_ ( .A1(_06678_ ), .A2(_02864_ ), .ZN(_06785_ ) );
NOR3_X1 _14804_ ( .A1(_06784_ ), .A2(_06785_ ), .A3(_06751_ ), .ZN(_06786_ ) );
NOR2_X1 _14805_ ( .A1(_06678_ ), .A2(_02695_ ), .ZN(_06787_ ) );
AOI21_X1 _14806_ ( .A(_02766_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06788_ ) );
NOR3_X1 _14807_ ( .A1(_06787_ ), .A2(_06747_ ), .A3(_06788_ ), .ZN(_06789_ ) );
BUF_X2 _14808_ ( .A(_06673_ ), .Z(_06790_ ) );
OR3_X1 _14809_ ( .A1(_06786_ ), .A2(_06789_ ), .A3(_06790_ ), .ZN(_06791_ ) );
BUF_X4 _14810_ ( .A(_05015_ ), .Z(_06792_ ) );
BUF_X4 _14811_ ( .A(_06792_ ), .Z(_06793_ ) );
BUF_X4 _14812_ ( .A(_06625_ ), .Z(_06794_ ) );
BUF_X2 _14813_ ( .A(_06794_ ), .Z(_06795_ ) );
BUF_X2 _14814_ ( .A(_06795_ ), .Z(_06796_ ) );
NOR2_X1 _14815_ ( .A1(_06680_ ), .A2(_04743_ ), .ZN(_06797_ ) );
AOI21_X1 _14816_ ( .A(_02717_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06798_ ) );
NOR3_X1 _14817_ ( .A1(_06797_ ), .A2(_06751_ ), .A3(_06798_ ), .ZN(_06799_ ) );
OR2_X1 _14818_ ( .A1(_06799_ ), .A2(_06760_ ), .ZN(_06800_ ) );
NAND4_X1 _14819_ ( .A1(_06791_ ), .A2(_06793_ ), .A3(_06796_ ), .A4(_06800_ ), .ZN(_06801_ ) );
AOI21_X1 _14820_ ( .A(_06740_ ), .B1(_06783_ ), .B2(_06801_ ), .ZN(_06802_ ) );
NOR3_X1 _14821_ ( .A1(_04923_ ), .A2(_04924_ ), .A3(_05195_ ), .ZN(_06803_ ) );
INV_X1 _14822_ ( .A(_04866_ ), .ZN(_06804_ ) );
OR3_X1 _14823_ ( .A1(_04921_ ), .A2(_04922_ ), .A3(_06804_ ), .ZN(_06805_ ) );
OAI21_X1 _14824_ ( .A(_06805_ ), .B1(_04923_ ), .B2(_04871_ ), .ZN(_06806_ ) );
NOR4_X1 _14825_ ( .A1(_06738_ ), .A2(_06802_ ), .A3(_06803_ ), .A4(_06806_ ), .ZN(_06807_ ) );
NAND3_X1 _14826_ ( .A1(_06619_ ), .A2(_06733_ ), .A3(_06807_ ), .ZN(_06808_ ) );
INV_X1 _14827_ ( .A(_06536_ ), .ZN(_06809_ ) );
NAND3_X1 _14828_ ( .A1(_06809_ ), .A2(_06522_ ), .A3(_06526_ ), .ZN(_06810_ ) );
AND4_X1 _14829_ ( .A1(\ID_EX_typ [3] ), .A2(_04869_ ), .A3(_04867_ ), .A4(\ID_EX_typ [0] ), .ZN(_06811_ ) );
MUX2_X1 _14830_ ( .A(_06811_ ), .B(_06535_ ), .S(\ID_EX_typ [4] ), .Z(_06812_ ) );
NOR2_X1 _14831_ ( .A1(_06810_ ), .A2(_06812_ ), .ZN(_06813_ ) );
NOR2_X1 _14832_ ( .A1(_06813_ ), .A2(_06541_ ), .ZN(_06814_ ) );
INV_X2 _14833_ ( .A(_06814_ ), .ZN(_06815_ ) );
BUF_X4 _14834_ ( .A(_06815_ ), .Z(_06816_ ) );
AOI21_X1 _14835_ ( .A(_06544_ ), .B1(_06808_ ), .B2(_06816_ ), .ZN(_06817_ ) );
OAI21_X1 _14836_ ( .A(_06374_ ), .B1(_05946_ ), .B2(_05506_ ), .ZN(_06818_ ) );
OAI21_X1 _14837_ ( .A(_06517_ ), .B1(_06817_ ), .B2(_06818_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
OR2_X1 _14838_ ( .A1(_06266_ ), .A2(_06228_ ), .ZN(_06819_ ) );
BUF_X2 _14839_ ( .A(_06536_ ), .Z(_06820_ ) );
OAI21_X1 _14840_ ( .A(_06820_ ), .B1(_06530_ ), .B2(_06531_ ), .ZN(_06821_ ) );
AOI21_X1 _14841_ ( .A(_06821_ ), .B1(_06531_ ), .B2(_06530_ ), .ZN(_06822_ ) );
BUF_X4 _14842_ ( .A(_06521_ ), .Z(_06823_ ) );
BUF_X2 _14843_ ( .A(_06823_ ), .Z(_06824_ ) );
AND2_X1 _14844_ ( .A1(_05348_ ), .A2(_06824_ ), .ZN(_06825_ ) );
AND3_X1 _14845_ ( .A1(_06524_ ), .A2(\ID_EX_imm [20] ), .A3(_06520_ ), .ZN(_06826_ ) );
NOR3_X1 _14846_ ( .A1(_06822_ ), .A2(_06825_ ), .A3(_06826_ ), .ZN(_06827_ ) );
OAI21_X1 _14847_ ( .A(_06518_ ), .B1(_06827_ ), .B2(_06543_ ), .ZN(_06828_ ) );
NAND3_X1 _14848_ ( .A1(_06655_ ), .A2(_06622_ ), .A3(_06677_ ), .ZN(_06829_ ) );
NAND2_X1 _14849_ ( .A1(_06676_ ), .A2(_06829_ ), .ZN(_06830_ ) );
NAND2_X1 _14850_ ( .A1(_06830_ ), .A2(_06689_ ), .ZN(_06831_ ) );
AOI21_X1 _14851_ ( .A(_06672_ ), .B1(_06831_ ), .B2(_06691_ ), .ZN(_06832_ ) );
NOR2_X1 _14852_ ( .A1(_05044_ ), .A2(_02940_ ), .ZN(_06833_ ) );
AOI21_X1 _14853_ ( .A(_02271_ ), .B1(_06704_ ), .B2(_06706_ ), .ZN(_06834_ ) );
NOR2_X1 _14854_ ( .A1(_06833_ ), .A2(_06834_ ), .ZN(_06835_ ) );
NOR2_X1 _14855_ ( .A1(_06835_ ), .A2(_06698_ ), .ZN(_06836_ ) );
INV_X1 _14856_ ( .A(_02248_ ), .ZN(_06837_ ) );
NAND3_X1 _14857_ ( .A1(_06837_ ), .A2(_06704_ ), .A3(_06706_ ), .ZN(_06838_ ) );
AOI21_X1 _14858_ ( .A(_02965_ ), .B1(_05042_ ), .B2(_05043_ ), .ZN(_06839_ ) );
INV_X1 _14859_ ( .A(_06839_ ), .ZN(_06840_ ) );
AOI21_X1 _14860_ ( .A(_05040_ ), .B1(_06838_ ), .B2(_06840_ ), .ZN(_06841_ ) );
OR3_X1 _14861_ ( .A1(_06836_ ), .A2(_05028_ ), .A3(_06841_ ), .ZN(_06842_ ) );
NOR2_X1 _14862_ ( .A1(_06710_ ), .A2(_04477_ ), .ZN(_06843_ ) );
AOI21_X1 _14863_ ( .A(_02382_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06844_ ) );
OAI21_X1 _14864_ ( .A(_06682_ ), .B1(_06843_ ), .B2(_06844_ ), .ZN(_06845_ ) );
NOR2_X1 _14865_ ( .A1(_06710_ ), .A2(_02307_ ), .ZN(_06846_ ) );
AOI21_X1 _14866_ ( .A(_02333_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06847_ ) );
OAI21_X1 _14867_ ( .A(_06699_ ), .B1(_06846_ ), .B2(_06847_ ), .ZN(_06848_ ) );
BUF_X2 _14868_ ( .A(_05028_ ), .Z(_06849_ ) );
NAND3_X1 _14869_ ( .A1(_06845_ ), .A2(_06848_ ), .A3(_06849_ ), .ZN(_06850_ ) );
NAND2_X1 _14870_ ( .A1(_06842_ ), .A2(_06850_ ), .ZN(_06851_ ) );
NAND2_X1 _14871_ ( .A1(_02976_ ), .A2(_05044_ ), .ZN(_06852_ ) );
NAND3_X1 _14872_ ( .A1(_04894_ ), .A2(_06704_ ), .A3(_06706_ ), .ZN(_06853_ ) );
AND3_X1 _14873_ ( .A1(_06852_ ), .A2(_05040_ ), .A3(_06853_ ), .ZN(_06854_ ) );
AND3_X1 _14874_ ( .A1(_02160_ ), .A2(_02171_ ), .A3(_05044_ ), .ZN(_06855_ ) );
AOI21_X1 _14875_ ( .A(_06855_ ), .B1(_04878_ ), .B2(_06694_ ), .ZN(_06856_ ) );
AOI21_X1 _14876_ ( .A(_06854_ ), .B1(_06856_ ), .B2(_06699_ ), .ZN(_06857_ ) );
NOR2_X1 _14877_ ( .A1(_06857_ ), .A2(_06673_ ), .ZN(_06858_ ) );
MUX2_X1 _14878_ ( .A(_06851_ ), .B(_06858_ ), .S(_06762_ ), .Z(_06859_ ) );
AND2_X1 _14879_ ( .A1(_06859_ ), .A2(_06730_ ), .ZN(_06860_ ) );
OAI21_X1 _14880_ ( .A(_06620_ ), .B1(_06832_ ), .B2(_06860_ ), .ZN(_06861_ ) );
AOI21_X1 _14881_ ( .A(_06552_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06862_ ) );
AND2_X1 _14882_ ( .A1(_06862_ ), .A2(_06715_ ), .ZN(_06863_ ) );
INV_X1 _14883_ ( .A(_06863_ ), .ZN(_06864_ ) );
NOR2_X1 _14884_ ( .A1(_06710_ ), .A2(_02717_ ), .ZN(_06865_ ) );
AOI21_X1 _14885_ ( .A(_02695_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06866_ ) );
NOR3_X1 _14886_ ( .A1(_06865_ ), .A2(_06683_ ), .A3(_06866_ ), .ZN(_06867_ ) );
NOR2_X1 _14887_ ( .A1(_06678_ ), .A2(_02766_ ), .ZN(_06868_ ) );
AOI21_X1 _14888_ ( .A(_02864_ ), .B1(_06704_ ), .B2(_06706_ ), .ZN(_06869_ ) );
NOR3_X1 _14889_ ( .A1(_06868_ ), .A2(_06700_ ), .A3(_06869_ ), .ZN(_06870_ ) );
NOR2_X1 _14890_ ( .A1(_06867_ ), .A2(_06870_ ), .ZN(_06871_ ) );
BUF_X4 _14891_ ( .A(_06723_ ), .Z(_06872_ ) );
MUX2_X1 _14892_ ( .A(_06864_ ), .B(_06871_ ), .S(_06872_ ), .Z(_06873_ ) );
NOR2_X1 _14893_ ( .A1(_06873_ ), .A2(_06763_ ), .ZN(_06874_ ) );
NOR2_X1 _14894_ ( .A1(_06710_ ), .A2(_02624_ ), .ZN(_06875_ ) );
AOI21_X1 _14895_ ( .A(_02647_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06876_ ) );
NOR3_X1 _14896_ ( .A1(_06875_ ), .A2(_06876_ ), .A3(_06683_ ), .ZN(_06877_ ) );
NOR2_X1 _14897_ ( .A1(_06678_ ), .A2(_02670_ ), .ZN(_06878_ ) );
AOI21_X1 _14898_ ( .A(_02574_ ), .B1(_06704_ ), .B2(_06706_ ), .ZN(_06879_ ) );
NOR3_X1 _14899_ ( .A1(_06878_ ), .A2(_06700_ ), .A3(_06879_ ), .ZN(_06880_ ) );
OAI21_X1 _14900_ ( .A(_06724_ ), .B1(_06877_ ), .B2(_06880_ ), .ZN(_06881_ ) );
NOR2_X1 _14901_ ( .A1(_06679_ ), .A2(_02841_ ), .ZN(_06882_ ) );
AOI21_X1 _14902_ ( .A(_02792_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06883_ ) );
NOR3_X1 _14903_ ( .A1(_06882_ ), .A2(_06683_ ), .A3(_06883_ ), .ZN(_06884_ ) );
NOR2_X1 _14904_ ( .A1(_06710_ ), .A2(_02816_ ), .ZN(_06885_ ) );
AOI21_X1 _14905_ ( .A(_02600_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06886_ ) );
NOR3_X1 _14906_ ( .A1(_06885_ ), .A2(_06700_ ), .A3(_06886_ ), .ZN(_06887_ ) );
OAI21_X1 _14907_ ( .A(_06693_ ), .B1(_06884_ ), .B2(_06887_ ), .ZN(_06888_ ) );
NAND2_X1 _14908_ ( .A1(_06881_ ), .A2(_06888_ ), .ZN(_06889_ ) );
AOI21_X1 _14909_ ( .A(_02526_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06890_ ) );
INV_X1 _14910_ ( .A(_06890_ ), .ZN(_06891_ ) );
OAI211_X1 _14911_ ( .A(_06891_ ), .B(_06700_ ), .C1(_02552_ ), .C2(_06680_ ), .ZN(_06892_ ) );
AOI21_X1 _14912_ ( .A(_02480_ ), .B1(_06705_ ), .B2(_06707_ ), .ZN(_06893_ ) );
INV_X1 _14913_ ( .A(_06893_ ), .ZN(_06894_ ) );
OAI211_X1 _14914_ ( .A(_06894_ ), .B(_06746_ ), .C1(_02503_ ), .C2(_06680_ ), .ZN(_06895_ ) );
AND3_X1 _14915_ ( .A1(_06892_ ), .A2(_06895_ ), .A3(_06703_ ), .ZN(_06896_ ) );
NOR2_X1 _14916_ ( .A1(_06710_ ), .A2(_02458_ ), .ZN(_06897_ ) );
AOI21_X1 _14917_ ( .A(_02406_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06898_ ) );
OAI21_X1 _14918_ ( .A(_06719_ ), .B1(_06897_ ), .B2(_06898_ ), .ZN(_06899_ ) );
NOR2_X1 _14919_ ( .A1(_06678_ ), .A2(_04330_ ), .ZN(_06900_ ) );
OAI21_X1 _14920_ ( .A(_06715_ ), .B1(_06900_ ), .B2(_06844_ ), .ZN(_06901_ ) );
AOI21_X1 _14921_ ( .A(_06703_ ), .B1(_06899_ ), .B2(_06901_ ), .ZN(_06902_ ) );
NOR2_X1 _14922_ ( .A1(_06896_ ), .A2(_06902_ ), .ZN(_06903_ ) );
MUX2_X1 _14923_ ( .A(_06889_ ), .B(_06903_ ), .S(_06727_ ), .Z(_06904_ ) );
MUX2_X1 _14924_ ( .A(_06874_ ), .B(_06904_ ), .S(_06730_ ), .Z(_06905_ ) );
NAND2_X1 _14925_ ( .A1(_06905_ ), .A2(_06739_ ), .ZN(_06906_ ) );
BUF_X2 _14926_ ( .A(_06737_ ), .Z(_06907_ ) );
NAND3_X1 _14927_ ( .A1(_06859_ ), .A2(_06731_ ), .A3(_06907_ ), .ZN(_06908_ ) );
NAND3_X1 _14928_ ( .A1(_06861_ ), .A2(_06906_ ), .A3(_06908_ ), .ZN(_06909_ ) );
AND2_X2 _14929_ ( .A1(_06602_ ), .A2(_06611_ ), .ZN(_06910_ ) );
OAI21_X1 _14930_ ( .A(_06616_ ), .B1(_06910_ ), .B2(_06545_ ), .ZN(_06911_ ) );
AOI21_X1 _14931_ ( .A(_06911_ ), .B1(_06545_ ), .B2(_06910_ ), .ZN(_06912_ ) );
BUF_X2 _14932_ ( .A(_05194_ ), .Z(_06913_ ) );
AND2_X1 _14933_ ( .A1(_04955_ ), .A2(_06913_ ), .ZN(_06914_ ) );
NOR3_X1 _14934_ ( .A1(_04918_ ), .A2(_06613_ ), .A3(_06804_ ), .ZN(_06915_ ) );
AOI21_X1 _14935_ ( .A(_04871_ ), .B1(_04918_ ), .B2(_06613_ ), .ZN(_06916_ ) );
OR3_X1 _14936_ ( .A1(_06914_ ), .A2(_06915_ ), .A3(_06916_ ), .ZN(_06917_ ) );
OR3_X1 _14937_ ( .A1(_06909_ ), .A2(_06912_ ), .A3(_06917_ ), .ZN(_06918_ ) );
AOI21_X1 _14938_ ( .A(_06828_ ), .B1(_06918_ ), .B2(_06816_ ), .ZN(_06919_ ) );
OAI21_X1 _14939_ ( .A(_06374_ ), .B1(_05351_ ), .B2(_05506_ ), .ZN(_06920_ ) );
OAI21_X1 _14940_ ( .A(_06819_ ), .B1(_06919_ ), .B2(_06920_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
CLKBUF_X2 _14941_ ( .A(_06227_ ), .Z(_06921_ ) );
OR2_X1 _14942_ ( .A1(_06277_ ), .A2(_06921_ ), .ZN(_06922_ ) );
BUF_X4 _14943_ ( .A(_06525_ ), .Z(_06923_ ) );
AOI22_X1 _14944_ ( .A1(_05408_ ), .A2(_06824_ ), .B1(\ID_EX_imm [19] ), .B2(_06923_ ), .ZN(_06924_ ) );
NAND3_X1 _14945_ ( .A1(_05150_ ), .A2(_04357_ ), .A3(_04380_ ), .ZN(_06925_ ) );
NAND2_X1 _14946_ ( .A1(_06925_ ), .A2(_05157_ ), .ZN(_06926_ ) );
AND2_X1 _14947_ ( .A1(_06926_ ), .A2(_04306_ ), .ZN(_06927_ ) );
OR3_X1 _14948_ ( .A1(_06927_ ), .A2(_04331_ ), .A3(_05152_ ), .ZN(_06928_ ) );
OAI21_X1 _14949_ ( .A(_04331_ ), .B1(_06927_ ), .B2(_05152_ ), .ZN(_06929_ ) );
NAND3_X1 _14950_ ( .A1(_06928_ ), .A2(_06820_ ), .A3(_06929_ ), .ZN(_06930_ ) );
AOI21_X1 _14951_ ( .A(_06542_ ), .B1(_06924_ ), .B2(_06930_ ), .ZN(_06931_ ) );
CLKBUF_X2 _14952_ ( .A(_03885_ ), .Z(_06932_ ) );
OR2_X1 _14953_ ( .A1(_06931_ ), .A2(_06932_ ), .ZN(_06933_ ) );
INV_X1 _14954_ ( .A(_06616_ ), .ZN(_06934_ ) );
BUF_X2 _14955_ ( .A(_06934_ ), .Z(_06935_ ) );
NAND2_X1 _14956_ ( .A1(_06600_ ), .A2(_06601_ ), .ZN(_06936_ ) );
AOI21_X1 _14957_ ( .A(_04949_ ), .B1(_06936_ ), .B2(_06605_ ), .ZN(_06937_ ) );
OR3_X1 _14958_ ( .A1(_06937_ ), .A2(_04944_ ), .A3(_06609_ ), .ZN(_06938_ ) );
OAI21_X1 _14959_ ( .A(_04944_ ), .B1(_06937_ ), .B2(_06609_ ), .ZN(_06939_ ) );
AOI21_X1 _14960_ ( .A(_06935_ ), .B1(_06938_ ), .B2(_06939_ ), .ZN(_06940_ ) );
NOR3_X1 _14961_ ( .A1(_06716_ ), .A2(_06746_ ), .A3(_06717_ ), .ZN(_06941_ ) );
NOR3_X1 _14962_ ( .A1(_06755_ ), .A2(_06750_ ), .A3(_06758_ ), .ZN(_06942_ ) );
NOR3_X1 _14963_ ( .A1(_06941_ ), .A2(_06942_ ), .A3(_06673_ ), .ZN(_06943_ ) );
NOR3_X1 _14964_ ( .A1(_06720_ ), .A2(_06750_ ), .A3(_06721_ ), .ZN(_06944_ ) );
NOR3_X1 _14965_ ( .A1(_06711_ ), .A2(_06712_ ), .A3(_06746_ ), .ZN(_06945_ ) );
NOR3_X1 _14966_ ( .A1(_06944_ ), .A2(_06945_ ), .A3(_06723_ ), .ZN(_06946_ ) );
NOR2_X1 _14967_ ( .A1(_06943_ ), .A2(_06946_ ), .ZN(_06947_ ) );
NAND4_X1 _14968_ ( .A1(_06703_ ), .A2(_03005_ ), .A3(_06715_ ), .A4(_06680_ ), .ZN(_06948_ ) );
AOI211_X1 _14969_ ( .A(_06699_ ), .B(_06708_ ), .C1(_02976_ ), .C2(_06694_ ), .ZN(_06949_ ) );
AND3_X1 _14970_ ( .A1(_06695_ ), .A2(_06750_ ), .A3(_06696_ ), .ZN(_06950_ ) );
NOR2_X1 _14971_ ( .A1(_06949_ ), .A2(_06950_ ), .ZN(_06951_ ) );
OAI21_X1 _14972_ ( .A(_06948_ ), .B1(_06951_ ), .B2(_06693_ ), .ZN(_06952_ ) );
MUX2_X1 _14973_ ( .A(_06947_ ), .B(_06952_ ), .S(_06762_ ), .Z(_06953_ ) );
NAND3_X1 _14974_ ( .A1(_06953_ ), .A2(_06731_ ), .A3(_06907_ ), .ZN(_06954_ ) );
BUF_X4 _14975_ ( .A(_04870_ ), .Z(_06955_ ) );
OAI21_X1 _14976_ ( .A(_06955_ ), .B1(_04953_ ), .B2(_04330_ ), .ZN(_06956_ ) );
NAND2_X1 _14977_ ( .A1(_06954_ ), .A2(_06956_ ), .ZN(_06957_ ) );
NOR3_X1 _14978_ ( .A1(_06787_ ), .A2(_06698_ ), .A3(_06788_ ), .ZN(_06958_ ) );
AOI21_X1 _14979_ ( .A(_06798_ ), .B1(_06694_ ), .B2(_06552_ ), .ZN(_06959_ ) );
AOI21_X1 _14980_ ( .A(_06958_ ), .B1(_06750_ ), .B2(_06959_ ), .ZN(_06960_ ) );
NOR2_X1 _14981_ ( .A1(_06960_ ), .A2(_06673_ ), .ZN(_06961_ ) );
AND2_X1 _14982_ ( .A1(_06961_ ), .A2(_06625_ ), .ZN(_06962_ ) );
OAI21_X1 _14983_ ( .A(_06739_ ), .B1(_06962_ ), .B2(_06627_ ), .ZN(_06963_ ) );
NOR3_X1 _14984_ ( .A1(_06749_ ), .A2(_06752_ ), .A3(_06681_ ), .ZN(_06964_ ) );
NOR3_X1 _14985_ ( .A1(_06757_ ), .A2(_06698_ ), .A3(_06758_ ), .ZN(_06965_ ) );
NOR2_X1 _14986_ ( .A1(_06964_ ), .A2(_06965_ ), .ZN(_06966_ ) );
NAND2_X1 _14987_ ( .A1(_06966_ ), .A2(_06849_ ), .ZN(_06967_ ) );
OAI21_X1 _14988_ ( .A(_06682_ ), .B1(_06742_ ), .B2(_06745_ ), .ZN(_06968_ ) );
OAI21_X1 _14989_ ( .A(_06698_ ), .B1(_06771_ ), .B2(_06772_ ), .ZN(_06969_ ) );
NAND2_X1 _14990_ ( .A1(_06968_ ), .A2(_06969_ ), .ZN(_06970_ ) );
NAND2_X1 _14991_ ( .A1(_06970_ ), .A2(_05048_ ), .ZN(_06971_ ) );
NAND2_X1 _14992_ ( .A1(_06967_ ), .A2(_06971_ ), .ZN(_06972_ ) );
NOR3_X1 _14993_ ( .A1(_06784_ ), .A2(_06785_ ), .A3(_06681_ ), .ZN(_06973_ ) );
NOR3_X1 _14994_ ( .A1(_06778_ ), .A2(_06698_ ), .A3(_06779_ ), .ZN(_06974_ ) );
OR3_X1 _14995_ ( .A1(_06973_ ), .A2(_06974_ ), .A3(_05028_ ), .ZN(_06975_ ) );
NOR3_X1 _14996_ ( .A1(_06775_ ), .A2(_06681_ ), .A3(_06776_ ), .ZN(_06976_ ) );
NOR3_X1 _14997_ ( .A1(_06768_ ), .A2(_06698_ ), .A3(_06769_ ), .ZN(_06977_ ) );
NOR2_X1 _14998_ ( .A1(_06976_ ), .A2(_06977_ ), .ZN(_06978_ ) );
NAND2_X1 _14999_ ( .A1(_06978_ ), .A2(_06849_ ), .ZN(_06979_ ) );
NAND2_X1 _15000_ ( .A1(_06975_ ), .A2(_06979_ ), .ZN(_06980_ ) );
MUX2_X1 _15001_ ( .A(_06972_ ), .B(_06980_ ), .S(_05033_ ), .Z(_06981_ ) );
AOI21_X1 _15002_ ( .A(_06963_ ), .B1(_06729_ ), .B2(_06981_ ), .ZN(_06982_ ) );
BUF_X4 _15003_ ( .A(_04866_ ), .Z(_06983_ ) );
AOI221_X4 _15004_ ( .A(_06982_ ), .B1(_06607_ ), .B2(_06983_ ), .C1(_04943_ ), .C2(_05194_ ), .ZN(_06984_ ) );
BUF_X2 _15005_ ( .A(_06666_ ), .Z(_06985_ ) );
BUF_X2 _15006_ ( .A(_06675_ ), .Z(_06986_ ) );
AND4_X1 _15007_ ( .A1(_06689_ ), .A2(_06985_ ), .A3(_06986_ ), .A4(_06667_ ), .ZN(_06987_ ) );
AND2_X1 _15008_ ( .A1(_06953_ ), .A2(_06734_ ), .ZN(_06988_ ) );
AND2_X1 _15009_ ( .A1(_06667_ ), .A2(_06669_ ), .ZN(_06989_ ) );
AND2_X1 _15010_ ( .A1(_06666_ ), .A2(_06989_ ), .ZN(_06990_ ) );
NOR3_X1 _15011_ ( .A1(_06987_ ), .A2(_06988_ ), .A3(_06990_ ), .ZN(_06991_ ) );
INV_X1 _15012_ ( .A(_06620_ ), .ZN(_06992_ ) );
BUF_X4 _15013_ ( .A(_06992_ ), .Z(_06993_ ) );
OAI21_X1 _15014_ ( .A(_06984_ ), .B1(_06991_ ), .B2(_06993_ ), .ZN(_06994_ ) );
OR3_X1 _15015_ ( .A1(_06940_ ), .A2(_06957_ ), .A3(_06994_ ), .ZN(_06995_ ) );
AOI21_X1 _15016_ ( .A(_06933_ ), .B1(_06995_ ), .B2(_06816_ ), .ZN(_06996_ ) );
OAI21_X1 _15017_ ( .A(_06374_ ), .B1(_05375_ ), .B2(_05506_ ), .ZN(_06997_ ) );
OAI21_X1 _15018_ ( .A(_06922_ ), .B1(_06996_ ), .B2(_06997_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
OR2_X1 _15019_ ( .A1(_05430_ ), .A2(_06921_ ), .ZN(_06998_ ) );
AOI22_X1 _15020_ ( .A1(_05413_ ), .A2(_06824_ ), .B1(\ID_EX_imm [18] ), .B2(_06923_ ), .ZN(_06999_ ) );
BUF_X2 _15021_ ( .A(_06809_ ), .Z(_07000_ ) );
AOI21_X1 _15022_ ( .A(_07000_ ), .B1(_06926_ ), .B2(_04306_ ), .ZN(_07001_ ) );
OAI21_X1 _15023_ ( .A(_07001_ ), .B1(_04306_ ), .B2(_06926_ ), .ZN(_07002_ ) );
AOI21_X1 _15024_ ( .A(_06542_ ), .B1(_06999_ ), .B2(_07002_ ), .ZN(_07003_ ) );
OR2_X1 _15025_ ( .A1(_07003_ ), .A2(_06932_ ), .ZN(_07004_ ) );
AND3_X1 _15026_ ( .A1(_06985_ ), .A2(_06688_ ), .A3(_06675_ ), .ZN(_07005_ ) );
NOR2_X1 _15027_ ( .A1(_06751_ ), .A2(_06680_ ), .ZN(_07006_ ) );
INV_X1 _15028_ ( .A(_07006_ ), .ZN(_07007_ ) );
NAND2_X1 _15029_ ( .A1(_07005_ ), .A2(_07007_ ), .ZN(_07008_ ) );
AOI21_X1 _15030_ ( .A(_06672_ ), .B1(_07008_ ), .B2(_06691_ ), .ZN(_07009_ ) );
OAI21_X1 _15031_ ( .A(_06750_ ), .B1(_06843_ ), .B2(_06844_ ), .ZN(_07010_ ) );
OAI21_X1 _15032_ ( .A(_06746_ ), .B1(_06900_ ), .B2(_06898_ ), .ZN(_07011_ ) );
AOI21_X1 _15033_ ( .A(_06693_ ), .B1(_07010_ ), .B2(_07011_ ), .ZN(_07012_ ) );
OAI21_X1 _15034_ ( .A(_06682_ ), .B1(_06846_ ), .B2(_06847_ ), .ZN(_07013_ ) );
OAI21_X1 _15035_ ( .A(_06699_ ), .B1(_06833_ ), .B2(_06834_ ), .ZN(_07014_ ) );
AOI21_X1 _15036_ ( .A(_06724_ ), .B1(_07013_ ), .B2(_07014_ ), .ZN(_07015_ ) );
NOR2_X1 _15037_ ( .A1(_07012_ ), .A2(_07015_ ), .ZN(_07016_ ) );
AOI21_X1 _15038_ ( .A(_06681_ ), .B1(_06852_ ), .B2(_06853_ ), .ZN(_07017_ ) );
AOI21_X1 _15039_ ( .A(_06698_ ), .B1(_06838_ ), .B2(_06840_ ), .ZN(_07018_ ) );
OAI21_X1 _15040_ ( .A(_06724_ ), .B1(_07017_ ), .B2(_07018_ ), .ZN(_07019_ ) );
AND2_X1 _15041_ ( .A1(_06856_ ), .A2(_06715_ ), .ZN(_07020_ ) );
OAI21_X1 _15042_ ( .A(_07019_ ), .B1(_07020_ ), .B2(_06872_ ), .ZN(_07021_ ) );
INV_X1 _15043_ ( .A(_07021_ ), .ZN(_07022_ ) );
MUX2_X1 _15044_ ( .A(_07016_ ), .B(_07022_ ), .S(_06766_ ), .Z(_07023_ ) );
AND2_X1 _15045_ ( .A1(_07023_ ), .A2(_06765_ ), .ZN(_07024_ ) );
OAI21_X1 _15046_ ( .A(_06621_ ), .B1(_07009_ ), .B2(_07024_ ), .ZN(_07025_ ) );
OR3_X1 _15047_ ( .A1(_06897_ ), .A2(_06700_ ), .A3(_06898_ ), .ZN(_07026_ ) );
OAI211_X1 _15048_ ( .A(_06894_ ), .B(_06719_ ), .C1(_02503_ ), .C2(_06680_ ), .ZN(_07027_ ) );
NAND3_X1 _15049_ ( .A1(_07026_ ), .A2(_06872_ ), .A3(_07027_ ), .ZN(_07028_ ) );
OR3_X1 _15050_ ( .A1(_06878_ ), .A2(_06681_ ), .A3(_06879_ ), .ZN(_07029_ ) );
OAI211_X1 _15051_ ( .A(_06891_ ), .B(_06682_ ), .C1(_02552_ ), .C2(_06679_ ), .ZN(_07030_ ) );
NAND3_X1 _15052_ ( .A1(_07029_ ), .A2(_07030_ ), .A3(_06790_ ), .ZN(_07031_ ) );
AND2_X1 _15053_ ( .A1(_07028_ ), .A2(_07031_ ), .ZN(_07032_ ) );
OR2_X1 _15054_ ( .A1(_07032_ ), .A2(_06763_ ), .ZN(_07033_ ) );
NOR3_X1 _15055_ ( .A1(_06885_ ), .A2(_06682_ ), .A3(_06886_ ), .ZN(_07034_ ) );
NOR3_X1 _15056_ ( .A1(_06875_ ), .A2(_06699_ ), .A3(_06876_ ), .ZN(_07035_ ) );
NOR2_X1 _15057_ ( .A1(_07034_ ), .A2(_07035_ ), .ZN(_07036_ ) );
NOR2_X1 _15058_ ( .A1(_07036_ ), .A2(_06790_ ), .ZN(_07037_ ) );
BUF_X2 _15059_ ( .A(_06794_ ), .Z(_07038_ ) );
OR3_X1 _15060_ ( .A1(_06868_ ), .A2(_06681_ ), .A3(_06869_ ), .ZN(_07039_ ) );
INV_X1 _15061_ ( .A(_06883_ ), .ZN(_07040_ ) );
OAI211_X1 _15062_ ( .A(_07040_ ), .B(_06681_ ), .C1(_02841_ ), .C2(_06710_ ), .ZN(_07041_ ) );
AOI21_X1 _15063_ ( .A(_06872_ ), .B1(_07039_ ), .B2(_07041_ ), .ZN(_07042_ ) );
OR3_X1 _15064_ ( .A1(_07037_ ), .A2(_07038_ ), .A3(_07042_ ), .ZN(_07043_ ) );
AND3_X1 _15065_ ( .A1(_07033_ ), .A2(_06765_ ), .A3(_07043_ ), .ZN(_07044_ ) );
OAI21_X1 _15066_ ( .A(_06682_ ), .B1(_06865_ ), .B2(_06866_ ), .ZN(_07045_ ) );
OAI21_X1 _15067_ ( .A(_07045_ ), .B1(_06682_ ), .B2(_06862_ ), .ZN(_07046_ ) );
BUF_X2 _15068_ ( .A(_06790_ ), .Z(_07047_ ) );
NOR4_X1 _15069_ ( .A1(_07046_ ), .A2(_06730_ ), .A3(_06767_ ), .A4(_07047_ ), .ZN(_07048_ ) );
OAI21_X1 _15070_ ( .A(_06739_ ), .B1(_07044_ ), .B2(_07048_ ), .ZN(_07049_ ) );
BUF_X2 _15071_ ( .A(_05194_ ), .Z(_07050_ ) );
BUF_X4 _15072_ ( .A(_06983_ ), .Z(_07051_ ) );
AOI22_X1 _15073_ ( .A1(_04948_ ), .A2(_07050_ ), .B1(_06609_ ), .B2(_07051_ ), .ZN(_07052_ ) );
AND3_X1 _15074_ ( .A1(_07025_ ), .A2(_07049_ ), .A3(_07052_ ), .ZN(_07053_ ) );
AND3_X1 _15075_ ( .A1(_06936_ ), .A2(_04949_ ), .A3(_06605_ ), .ZN(_07054_ ) );
OR3_X1 _15076_ ( .A1(_07054_ ), .A2(_06937_ ), .A3(_06935_ ), .ZN(_07055_ ) );
BUF_X4 _15077_ ( .A(_04871_ ), .Z(_07056_ ) );
AOI21_X1 _15078_ ( .A(_07056_ ), .B1(_04947_ ), .B2(_06608_ ), .ZN(_07057_ ) );
AOI21_X1 _15079_ ( .A(_07057_ ), .B1(_07024_ ), .B2(_06907_ ), .ZN(_07058_ ) );
NAND3_X1 _15080_ ( .A1(_07053_ ), .A2(_07055_ ), .A3(_07058_ ), .ZN(_07059_ ) );
AOI21_X1 _15081_ ( .A(_07004_ ), .B1(_07059_ ), .B2(_06816_ ), .ZN(_07060_ ) );
BUF_X4 _15082_ ( .A(_06236_ ), .Z(_07061_ ) );
BUF_X4 _15083_ ( .A(_05207_ ), .Z(_07062_ ) );
OAI21_X1 _15084_ ( .A(_07061_ ), .B1(_05411_ ), .B2(_07062_ ), .ZN(_07063_ ) );
OAI21_X1 _15085_ ( .A(_06998_ ), .B1(_07060_ ), .B2(_07063_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
INV_X1 _15086_ ( .A(_06295_ ), .ZN(_07064_ ) );
AOI22_X1 _15087_ ( .A1(_05452_ ), .A2(_06824_ ), .B1(\ID_EX_imm [17] ), .B2(_06923_ ), .ZN(_07065_ ) );
INV_X1 _15088_ ( .A(_04380_ ), .ZN(_07066_ ) );
AOI21_X1 _15089_ ( .A(_07066_ ), .B1(_05136_ ), .B2(_05148_ ), .ZN(_07067_ ) );
OR3_X1 _15090_ ( .A1(_07067_ ), .A2(_04357_ ), .A3(_05155_ ), .ZN(_07068_ ) );
OAI21_X1 _15091_ ( .A(_04357_ ), .B1(_07067_ ), .B2(_05155_ ), .ZN(_07069_ ) );
NAND3_X1 _15092_ ( .A1(_07068_ ), .A2(_06820_ ), .A3(_07069_ ), .ZN(_07070_ ) );
AOI21_X1 _15093_ ( .A(_06542_ ), .B1(_07065_ ), .B2(_07070_ ), .ZN(_07071_ ) );
OR2_X1 _15094_ ( .A1(_07071_ ), .A2(_06932_ ), .ZN(_07072_ ) );
AND4_X1 _15095_ ( .A1(_05003_ ), .A2(_05008_ ), .A3(_04942_ ), .A4(_04947_ ), .ZN(_07073_ ) );
AND4_X1 _15096_ ( .A1(_06646_ ), .A2(_07073_ ), .A3(_06648_ ), .A4(_06647_ ), .ZN(_07074_ ) );
INV_X1 _15097_ ( .A(_05018_ ), .ZN(_07075_ ) );
OAI21_X1 _15098_ ( .A(_07074_ ), .B1(_07075_ ), .B2(_06628_ ), .ZN(_07076_ ) );
NOR4_X1 _15099_ ( .A1(_05003_ ), .A2(_05008_ ), .A3(_04942_ ), .A4(_04947_ ), .ZN(_07077_ ) );
NOR4_X1 _15100_ ( .A1(_04965_ ), .A2(_04972_ ), .A3(_04961_ ), .A4(_04977_ ), .ZN(_07078_ ) );
NOR4_X1 _15101_ ( .A1(_04921_ ), .A2(_04918_ ), .A3(_04933_ ), .A4(_04930_ ), .ZN(_07079_ ) );
NOR4_X1 _15102_ ( .A1(_04983_ ), .A2(_04988_ ), .A3(_04994_ ), .A4(_04998_ ), .ZN(_07080_ ) );
AND4_X1 _15103_ ( .A1(_07077_ ), .A2(_07078_ ), .A3(_07079_ ), .A4(_07080_ ), .ZN(_07081_ ) );
NAND3_X1 _15104_ ( .A1(_06629_ ), .A2(_07081_ ), .A3(_05018_ ), .ZN(_07082_ ) );
AOI221_X4 _15105_ ( .A(_04878_ ), .B1(_07076_ ), .B2(_07082_ ), .C1(_06654_ ), .C2(_06652_ ), .ZN(_07083_ ) );
AND2_X1 _15106_ ( .A1(_07083_ ), .A2(_06677_ ), .ZN(_07084_ ) );
NAND4_X1 _15107_ ( .A1(_07084_ ), .A2(_06689_ ), .A3(_06986_ ), .A4(_06684_ ), .ZN(_07085_ ) );
AOI22_X1 _15108_ ( .A1(_07085_ ), .A2(_06691_ ), .B1(_06671_ ), .B2(_06668_ ), .ZN(_07086_ ) );
OR3_X1 _15109_ ( .A1(_06709_ ), .A2(_06713_ ), .A3(_05048_ ), .ZN(_07087_ ) );
NAND3_X1 _15110_ ( .A1(_06697_ ), .A2(_06703_ ), .A3(_06701_ ), .ZN(_07088_ ) );
NAND3_X1 _15111_ ( .A1(_07087_ ), .A2(_06763_ ), .A3(_07088_ ), .ZN(_07089_ ) );
NAND3_X1 _15112_ ( .A1(_06718_ ), .A2(_06722_ ), .A3(_06693_ ), .ZN(_07090_ ) );
OAI21_X1 _15113_ ( .A(_06715_ ), .B1(_06757_ ), .B2(_06752_ ), .ZN(_07091_ ) );
OAI21_X1 _15114_ ( .A(_06719_ ), .B1(_06755_ ), .B2(_06758_ ), .ZN(_07092_ ) );
NAND3_X1 _15115_ ( .A1(_07091_ ), .A2(_07092_ ), .A3(_06724_ ), .ZN(_07093_ ) );
NAND2_X1 _15116_ ( .A1(_07090_ ), .A2(_07093_ ), .ZN(_07094_ ) );
BUF_X2 _15117_ ( .A(_06727_ ), .Z(_07095_ ) );
NAND2_X1 _15118_ ( .A1(_07094_ ), .A2(_07095_ ), .ZN(_07096_ ) );
AOI21_X1 _15119_ ( .A(_06792_ ), .B1(_07089_ ), .B2(_07096_ ), .ZN(_07097_ ) );
OAI21_X1 _15120_ ( .A(_06620_ ), .B1(_07086_ ), .B2(_07097_ ), .ZN(_07098_ ) );
BUF_X2 _15121_ ( .A(_06804_ ), .Z(_07099_ ) );
NOR3_X1 _15122_ ( .A1(_04933_ ), .A2(_04934_ ), .A3(_07099_ ), .ZN(_07100_ ) );
AOI21_X1 _15123_ ( .A(_07100_ ), .B1(_05080_ ), .B2(_07050_ ), .ZN(_07101_ ) );
OR3_X1 _15124_ ( .A1(_06786_ ), .A2(_06789_ ), .A3(_06760_ ), .ZN(_07102_ ) );
BUF_X4 _15125_ ( .A(_06763_ ), .Z(_07103_ ) );
NAND2_X1 _15126_ ( .A1(_06777_ ), .A2(_06780_ ), .ZN(_07104_ ) );
NAND2_X1 _15127_ ( .A1(_07104_ ), .A2(_06741_ ), .ZN(_07105_ ) );
NAND3_X1 _15128_ ( .A1(_07102_ ), .A2(_07103_ ), .A3(_07105_ ), .ZN(_07106_ ) );
NAND3_X1 _15129_ ( .A1(_06748_ ), .A2(_06741_ ), .A3(_06753_ ), .ZN(_07107_ ) );
BUF_X2 _15130_ ( .A(_06693_ ), .Z(_07108_ ) );
NAND3_X1 _15131_ ( .A1(_06770_ ), .A2(_06773_ ), .A3(_07108_ ), .ZN(_07109_ ) );
BUF_X2 _15132_ ( .A(_07038_ ), .Z(_07110_ ) );
NAND3_X1 _15133_ ( .A1(_07107_ ), .A2(_07109_ ), .A3(_07110_ ), .ZN(_07111_ ) );
AND3_X1 _15134_ ( .A1(_07106_ ), .A2(_06765_ ), .A3(_07111_ ), .ZN(_07112_ ) );
BUF_X4 _15135_ ( .A(_06747_ ), .Z(_07113_ ) );
AND3_X1 _15136_ ( .A1(_06959_ ), .A2(_06741_ ), .A3(_07113_ ), .ZN(_07114_ ) );
AND2_X1 _15137_ ( .A1(_07114_ ), .A2(_07110_ ), .ZN(_07115_ ) );
OAI21_X1 _15138_ ( .A(_06739_ ), .B1(_07115_ ), .B2(_06735_ ), .ZN(_07116_ ) );
OAI211_X1 _15139_ ( .A(_07098_ ), .B(_07101_ ), .C1(_07112_ ), .C2(_07116_ ), .ZN(_07117_ ) );
INV_X1 _15140_ ( .A(_05081_ ), .ZN(_07118_ ) );
AOI21_X1 _15141_ ( .A(_07118_ ), .B1(_06577_ ), .B2(_06598_ ), .ZN(_07119_ ) );
OR3_X1 _15142_ ( .A1(_07119_ ), .A2(_05080_ ), .A3(_06604_ ), .ZN(_07120_ ) );
OAI21_X1 _15143_ ( .A(_05080_ ), .B1(_07119_ ), .B2(_06604_ ), .ZN(_07121_ ) );
AND3_X1 _15144_ ( .A1(_07120_ ), .A2(_06617_ ), .A3(_07121_ ), .ZN(_07122_ ) );
NAND2_X1 _15145_ ( .A1(_07089_ ), .A2(_07096_ ), .ZN(_07123_ ) );
NAND3_X1 _15146_ ( .A1(_07123_ ), .A2(_06735_ ), .A3(_06737_ ), .ZN(_07124_ ) );
OAI21_X1 _15147_ ( .A(_07124_ ), .B1(_04935_ ), .B2(_07056_ ), .ZN(_07125_ ) );
OR3_X1 _15148_ ( .A1(_07117_ ), .A2(_07122_ ), .A3(_07125_ ), .ZN(_07126_ ) );
AOI21_X1 _15149_ ( .A(_07072_ ), .B1(_07126_ ), .B2(_06816_ ), .ZN(_07127_ ) );
NAND2_X1 _15150_ ( .A1(_05460_ ), .A2(_05280_ ), .ZN(_07128_ ) );
NAND2_X1 _15151_ ( .A1(_07128_ ), .A2(_06249_ ), .ZN(_07129_ ) );
OAI21_X1 _15152_ ( .A(_07064_ ), .B1(_07127_ ), .B2(_07129_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
OR2_X1 _15153_ ( .A1(_06307_ ), .A2(_06921_ ), .ZN(_07130_ ) );
OAI22_X1 _15154_ ( .A1(_05468_ ), .A2(_06523_ ), .B1(_02481_ ), .B2(_06527_ ), .ZN(_07131_ ) );
OAI21_X1 _15155_ ( .A(_06820_ ), .B1(_05149_ ), .B2(_07066_ ), .ZN(_07132_ ) );
AOI21_X1 _15156_ ( .A(_07132_ ), .B1(_07066_ ), .B2(_05149_ ), .ZN(_07133_ ) );
OAI21_X1 _15157_ ( .A(_06540_ ), .B1(_07131_ ), .B2(_07133_ ), .ZN(_07134_ ) );
NAND2_X1 _15158_ ( .A1(_07134_ ), .A2(_05343_ ), .ZN(_07135_ ) );
INV_X1 _15159_ ( .A(_06626_ ), .ZN(_07136_ ) );
AOI21_X1 _15160_ ( .A(_06668_ ), .B1(_06731_ ), .B2(_07136_ ), .ZN(_07137_ ) );
AOI21_X1 _15161_ ( .A(_06849_ ), .B1(_06845_ ), .B2(_06848_ ), .ZN(_07138_ ) );
OAI21_X1 _15162_ ( .A(_06682_ ), .B1(_06897_ ), .B2(_06893_ ), .ZN(_07139_ ) );
OAI21_X1 _15163_ ( .A(_06699_ ), .B1(_06900_ ), .B2(_06898_ ), .ZN(_07140_ ) );
AOI21_X1 _15164_ ( .A(_05048_ ), .B1(_07139_ ), .B2(_07140_ ), .ZN(_07141_ ) );
NOR2_X1 _15165_ ( .A1(_07138_ ), .A2(_07141_ ), .ZN(_07142_ ) );
OR3_X1 _15166_ ( .A1(_06836_ ), .A2(_05048_ ), .A3(_06841_ ), .ZN(_07143_ ) );
OAI21_X1 _15167_ ( .A(_07143_ ), .B1(_06857_ ), .B2(_06849_ ), .ZN(_07144_ ) );
MUX2_X1 _15168_ ( .A(_07142_ ), .B(_07144_ ), .S(_05033_ ), .Z(_07145_ ) );
AND2_X1 _15169_ ( .A1(_07145_ ), .A2(_06731_ ), .ZN(_07146_ ) );
OAI21_X1 _15170_ ( .A(_06621_ ), .B1(_07137_ ), .B2(_07146_ ), .ZN(_07147_ ) );
NOR2_X1 _15171_ ( .A1(_07119_ ), .A2(_06935_ ), .ZN(_07148_ ) );
OAI21_X1 _15172_ ( .A(_07148_ ), .B1(_05081_ ), .B2(_06600_ ), .ZN(_07149_ ) );
AND3_X1 _15173_ ( .A1(_06862_ ), .A2(_06741_ ), .A3(_07113_ ), .ZN(_07150_ ) );
NAND2_X1 _15174_ ( .A1(_07150_ ), .A2(_07110_ ), .ZN(_07151_ ) );
AOI21_X1 _15175_ ( .A(_06740_ ), .B1(_07151_ ), .B2(_06793_ ), .ZN(_07152_ ) );
NOR2_X1 _15176_ ( .A1(_06877_ ), .A2(_06880_ ), .ZN(_07153_ ) );
AND2_X1 _15177_ ( .A1(_06892_ ), .A2(_06895_ ), .ZN(_07154_ ) );
MUX2_X1 _15178_ ( .A(_07153_ ), .B(_07154_ ), .S(_06872_ ), .Z(_07155_ ) );
OAI21_X1 _15179_ ( .A(_06765_ ), .B1(_07155_ ), .B2(_07103_ ), .ZN(_07156_ ) );
OAI21_X1 _15180_ ( .A(_07047_ ), .B1(_06867_ ), .B2(_06870_ ), .ZN(_07157_ ) );
BUF_X4 _15181_ ( .A(_06760_ ), .Z(_07158_ ) );
OAI21_X1 _15182_ ( .A(_07158_ ), .B1(_06884_ ), .B2(_06887_ ), .ZN(_07159_ ) );
AOI21_X1 _15183_ ( .A(_07110_ ), .B1(_07157_ ), .B2(_07159_ ), .ZN(_07160_ ) );
OAI21_X1 _15184_ ( .A(_07152_ ), .B1(_07156_ ), .B2(_07160_ ), .ZN(_07161_ ) );
OR3_X1 _15185_ ( .A1(_04930_ ), .A2(_06603_ ), .A3(_07099_ ), .ZN(_07162_ ) );
OAI211_X1 _15186_ ( .A(_07161_ ), .B(_07162_ ), .C1(_07118_ ), .C2(_05195_ ), .ZN(_07163_ ) );
AND3_X1 _15187_ ( .A1(_07145_ ), .A2(_06735_ ), .A3(_06737_ ), .ZN(_07164_ ) );
AOI21_X1 _15188_ ( .A(_07056_ ), .B1(_04930_ ), .B2(_06603_ ), .ZN(_07165_ ) );
NOR3_X1 _15189_ ( .A1(_07163_ ), .A2(_07164_ ), .A3(_07165_ ), .ZN(_07166_ ) );
NAND3_X1 _15190_ ( .A1(_07147_ ), .A2(_07149_ ), .A3(_07166_ ), .ZN(_07167_ ) );
AOI21_X1 _15191_ ( .A(_07135_ ), .B1(_07167_ ), .B2(_06816_ ), .ZN(_07168_ ) );
OAI21_X1 _15192_ ( .A(_07061_ ), .B1(_05465_ ), .B2(_07062_ ), .ZN(_07169_ ) );
OAI21_X1 _15193_ ( .A(_07130_ ), .B1(_07168_ ), .B2(_07169_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OR2_X1 _15194_ ( .A1(_05501_ ), .A2(_06921_ ), .ZN(_07170_ ) );
INV_X1 _15195_ ( .A(_04647_ ), .ZN(_07171_ ) );
INV_X1 _15196_ ( .A(_04671_ ), .ZN(_07172_ ) );
NAND2_X1 _15197_ ( .A1(_05135_ ), .A2(_04575_ ), .ZN(_07173_ ) );
AOI211_X1 _15198_ ( .A(_07171_ ), .B(_07172_ ), .C1(_07173_ ), .C2(_05143_ ), .ZN(_07174_ ) );
OAI21_X1 _15199_ ( .A(_04623_ ), .B1(_07174_ ), .B2(_05147_ ), .ZN(_07175_ ) );
NAND2_X1 _15200_ ( .A1(_02526_ ), .A2(_04621_ ), .ZN(_07176_ ) );
AND2_X1 _15201_ ( .A1(_07175_ ), .A2(_07176_ ), .ZN(_07177_ ) );
XNOR2_X1 _15202_ ( .A(_07177_ ), .B(_04600_ ), .ZN(_07178_ ) );
NAND2_X1 _15203_ ( .A1(_07178_ ), .A2(_06537_ ), .ZN(_07179_ ) );
AOI22_X1 _15204_ ( .A1(_05491_ ), .A2(_06824_ ), .B1(\ID_EX_imm [15] ), .B2(_06923_ ), .ZN(_07180_ ) );
AOI21_X1 _15205_ ( .A(_06542_ ), .B1(_07179_ ), .B2(_07180_ ), .ZN(_07181_ ) );
OR2_X1 _15206_ ( .A1(_07181_ ), .A2(_06932_ ), .ZN(_07182_ ) );
INV_X1 _15207_ ( .A(_04962_ ), .ZN(_07183_ ) );
NAND2_X1 _15208_ ( .A1(_06573_ ), .A2(_06576_ ), .ZN(_07184_ ) );
AOI211_X1 _15209_ ( .A(_04974_ ), .B(_04979_ ), .C1(_07184_ ), .C2(_06587_ ), .ZN(_07185_ ) );
INV_X1 _15210_ ( .A(_07185_ ), .ZN(_07186_ ) );
AOI21_X1 _15211_ ( .A(_07183_ ), .B1(_07186_ ), .B2(_06595_ ), .ZN(_07187_ ) );
OR3_X1 _15212_ ( .A1(_07187_ ), .A2(_05056_ ), .A3(_06590_ ), .ZN(_07188_ ) );
OAI21_X1 _15213_ ( .A(_05056_ ), .B1(_07187_ ), .B2(_06590_ ), .ZN(_07189_ ) );
AND3_X1 _15214_ ( .A1(_07188_ ), .A2(_06617_ ), .A3(_07189_ ), .ZN(_07190_ ) );
AOI22_X1 _15215_ ( .A1(_05056_ ), .A2(_07050_ ), .B1(_04968_ ), .B2(_06955_ ), .ZN(_07191_ ) );
OAI21_X1 _15216_ ( .A(_07191_ ), .B1(_04967_ ), .B2(_07099_ ), .ZN(_07192_ ) );
BUF_X4 _15217_ ( .A(_06989_ ), .Z(_07193_ ) );
NAND2_X1 _15218_ ( .A1(_06985_ ), .A2(_07193_ ), .ZN(_07194_ ) );
OAI21_X1 _15219_ ( .A(_06703_ ), .B1(_06941_ ), .B2(_06942_ ), .ZN(_07195_ ) );
OAI21_X1 _15220_ ( .A(_06683_ ), .B1(_06749_ ), .B2(_06745_ ), .ZN(_07196_ ) );
OAI21_X1 _15221_ ( .A(_06700_ ), .B1(_06757_ ), .B2(_06752_ ), .ZN(_07197_ ) );
NAND2_X1 _15222_ ( .A1(_07196_ ), .A2(_07197_ ), .ZN(_07198_ ) );
OAI211_X1 _15223_ ( .A(_07195_ ), .B(_06794_ ), .C1(_06693_ ), .C2(_07198_ ), .ZN(_07199_ ) );
OAI21_X1 _15224_ ( .A(_06703_ ), .B1(_06949_ ), .B2(_06950_ ), .ZN(_07200_ ) );
OAI21_X1 _15225_ ( .A(_06723_ ), .B1(_06944_ ), .B2(_06945_ ), .ZN(_07201_ ) );
NAND2_X1 _15226_ ( .A1(_07200_ ), .A2(_07201_ ), .ZN(_07202_ ) );
OAI211_X1 _15227_ ( .A(_06627_ ), .B(_07199_ ), .C1(_07202_ ), .C2(_06727_ ), .ZN(_07203_ ) );
NAND4_X1 _15228_ ( .A1(_06623_ ), .A2(_03005_ ), .A3(_05015_ ), .A4(_06727_ ), .ZN(_07204_ ) );
AND2_X1 _15229_ ( .A1(_07203_ ), .A2(_07204_ ), .ZN(_07205_ ) );
AOI21_X1 _15230_ ( .A(_06992_ ), .B1(_07194_ ), .B2(_07205_ ), .ZN(_07206_ ) );
INV_X1 _15231_ ( .A(_06736_ ), .ZN(_07207_ ) );
BUF_X2 _15232_ ( .A(_07207_ ), .Z(_07208_ ) );
AOI21_X1 _15233_ ( .A(_07208_ ), .B1(_07203_ ), .B2(_07204_ ), .ZN(_07209_ ) );
NOR2_X1 _15234_ ( .A1(_06973_ ), .A2(_06974_ ), .ZN(_07210_ ) );
MUX2_X1 _15235_ ( .A(_07210_ ), .B(_06960_ ), .S(_06703_ ), .Z(_07211_ ) );
NAND2_X1 _15236_ ( .A1(_07211_ ), .A2(_06766_ ), .ZN(_07212_ ) );
NAND2_X1 _15237_ ( .A1(_06978_ ), .A2(_06790_ ), .ZN(_07213_ ) );
NAND2_X1 _15238_ ( .A1(_06970_ ), .A2(_06872_ ), .ZN(_07214_ ) );
NAND2_X1 _15239_ ( .A1(_07213_ ), .A2(_07214_ ), .ZN(_07215_ ) );
NAND2_X1 _15240_ ( .A1(_07215_ ), .A2(_07038_ ), .ZN(_07216_ ) );
AND2_X1 _15241_ ( .A1(_06627_ ), .A2(_05191_ ), .ZN(_07217_ ) );
AND3_X1 _15242_ ( .A1(_07212_ ), .A2(_07216_ ), .A3(_07217_ ), .ZN(_07218_ ) );
OR3_X1 _15243_ ( .A1(_07206_ ), .A2(_07209_ ), .A3(_07218_ ), .ZN(_07219_ ) );
OR3_X1 _15244_ ( .A1(_07190_ ), .A2(_07192_ ), .A3(_07219_ ), .ZN(_07220_ ) );
AOI21_X1 _15245_ ( .A(_07182_ ), .B1(_07220_ ), .B2(_06816_ ), .ZN(_07221_ ) );
OAI21_X1 _15246_ ( .A(_07061_ ), .B1(_05483_ ), .B2(_07062_ ), .ZN(_07222_ ) );
OAI21_X1 _15247_ ( .A(_07170_ ), .B1(_07221_ ), .B2(_07222_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
OR2_X1 _15248_ ( .A1(_05518_ ), .A2(_06921_ ), .ZN(_07223_ ) );
OR3_X1 _15249_ ( .A1(_07174_ ), .A2(_04623_ ), .A3(_05147_ ), .ZN(_07224_ ) );
NAND3_X1 _15250_ ( .A1(_07224_ ), .A2(_06537_ ), .A3(_07175_ ), .ZN(_07225_ ) );
AOI22_X1 _15251_ ( .A1(_05521_ ), .A2(_06824_ ), .B1(\ID_EX_imm [14] ), .B2(_06923_ ), .ZN(_07226_ ) );
AOI21_X1 _15252_ ( .A(_06542_ ), .B1(_07225_ ), .B2(_07226_ ), .ZN(_07227_ ) );
OR2_X1 _15253_ ( .A1(_07227_ ), .A2(_06932_ ), .ZN(_07228_ ) );
OAI211_X1 _15254_ ( .A(_06655_ ), .B(_06677_ ), .C1(_06790_ ), .C2(_07007_ ), .ZN(_07229_ ) );
INV_X1 _15255_ ( .A(_06666_ ), .ZN(_07230_ ) );
BUF_X4 _15256_ ( .A(_06687_ ), .Z(_07231_ ) );
OAI21_X1 _15257_ ( .A(_07229_ ), .B1(_07230_ ), .B2(_07231_ ), .ZN(_07232_ ) );
NAND2_X1 _15258_ ( .A1(_07232_ ), .A2(_07193_ ), .ZN(_07233_ ) );
NAND3_X1 _15259_ ( .A1(_07011_ ), .A2(_07010_ ), .A3(_06673_ ), .ZN(_07234_ ) );
NOR2_X1 _15260_ ( .A1(_06679_ ), .A2(_02503_ ), .ZN(_07235_ ) );
OAI21_X1 _15261_ ( .A(_06746_ ), .B1(_07235_ ), .B2(_06890_ ), .ZN(_07236_ ) );
OAI21_X1 _15262_ ( .A(_06750_ ), .B1(_06897_ ), .B2(_06893_ ), .ZN(_07237_ ) );
NAND3_X1 _15263_ ( .A1(_07236_ ), .A2(_07237_ ), .A3(_06723_ ), .ZN(_07238_ ) );
NAND3_X1 _15264_ ( .A1(_07234_ ), .A2(_07238_ ), .A3(_06625_ ), .ZN(_07239_ ) );
OR3_X1 _15265_ ( .A1(_07017_ ), .A2(_07018_ ), .A3(_05028_ ), .ZN(_07240_ ) );
NAND3_X1 _15266_ ( .A1(_07013_ ), .A2(_07014_ ), .A3(_06849_ ), .ZN(_07241_ ) );
NAND2_X1 _15267_ ( .A1(_07240_ ), .A2(_07241_ ), .ZN(_07242_ ) );
OAI211_X1 _15268_ ( .A(_06627_ ), .B(_07239_ ), .C1(_07242_ ), .C2(_06794_ ), .ZN(_07243_ ) );
NAND4_X1 _15269_ ( .A1(_07020_ ), .A2(_05015_ ), .A3(_06794_ ), .A4(_06872_ ), .ZN(_07244_ ) );
AND2_X1 _15270_ ( .A1(_07243_ ), .A2(_07244_ ), .ZN(_07245_ ) );
AOI21_X1 _15271_ ( .A(_06993_ ), .B1(_07233_ ), .B2(_07245_ ), .ZN(_07246_ ) );
NOR3_X1 _15272_ ( .A1(_07185_ ), .A2(_04962_ ), .A3(_06596_ ), .ZN(_07247_ ) );
NOR3_X1 _15273_ ( .A1(_07187_ ), .A2(_06934_ ), .A3(_07247_ ), .ZN(_07248_ ) );
OR2_X1 _15274_ ( .A1(_07245_ ), .A2(_07207_ ), .ZN(_07249_ ) );
BUF_X2 _15275_ ( .A(_07217_ ), .Z(_07250_ ) );
AND3_X1 _15276_ ( .A1(_07039_ ), .A2(_06849_ ), .A3(_07041_ ), .ZN(_07251_ ) );
AOI211_X1 _15277_ ( .A(_06625_ ), .B(_07251_ ), .C1(_06693_ ), .C2(_07046_ ), .ZN(_07252_ ) );
AND3_X1 _15278_ ( .A1(_07029_ ), .A2(_07030_ ), .A3(_06849_ ), .ZN(_07253_ ) );
NOR3_X1 _15279_ ( .A1(_07034_ ), .A2(_07035_ ), .A3(_06849_ ), .ZN(_07254_ ) );
NOR3_X1 _15280_ ( .A1(_07253_ ), .A2(_07254_ ), .A3(_06762_ ), .ZN(_07255_ ) );
OAI21_X1 _15281_ ( .A(_07250_ ), .B1(_07252_ ), .B2(_07255_ ), .ZN(_07256_ ) );
NAND2_X1 _15282_ ( .A1(_04962_ ), .A2(_06913_ ), .ZN(_07257_ ) );
NAND3_X1 _15283_ ( .A1(_05058_ ), .A2(_02526_ ), .A3(_06983_ ), .ZN(_07258_ ) );
AND4_X1 _15284_ ( .A1(_07249_ ), .A2(_07256_ ), .A3(_07257_ ), .A4(_07258_ ), .ZN(_07259_ ) );
OAI21_X1 _15285_ ( .A(_06955_ ), .B1(_05058_ ), .B2(_02526_ ), .ZN(_07260_ ) );
NAND2_X1 _15286_ ( .A1(_07259_ ), .A2(_07260_ ), .ZN(_07261_ ) );
OR3_X1 _15287_ ( .A1(_07246_ ), .A2(_07248_ ), .A3(_07261_ ), .ZN(_07262_ ) );
AOI21_X1 _15288_ ( .A(_07228_ ), .B1(_07262_ ), .B2(_06816_ ), .ZN(_07263_ ) );
NAND2_X1 _15289_ ( .A1(_05523_ ), .A2(_05280_ ), .ZN(_07264_ ) );
NAND2_X1 _15290_ ( .A1(_07264_ ), .A2(_06249_ ), .ZN(_07265_ ) );
OAI21_X1 _15291_ ( .A(_07223_ ), .B1(_07263_ ), .B2(_07265_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
AND4_X1 _15292_ ( .A1(\mycsreg.CSReg[0][13] ), .A2(_05331_ ), .A3(_05444_ ), .A4(_05394_ ), .ZN(_07266_ ) );
AND4_X1 _15293_ ( .A1(\mtvec [13] ), .A2(_05392_ ), .A3(_05444_ ), .A4(_05394_ ), .ZN(_07267_ ) );
NOR4_X1 _15294_ ( .A1(_05529_ ), .A2(_05538_ ), .A3(_07266_ ), .A4(_07267_ ), .ZN(_07268_ ) );
NAND3_X1 _15295_ ( .A1(_05315_ ), .A2(_05319_ ), .A3(_07268_ ), .ZN(_07269_ ) );
OAI211_X1 _15296_ ( .A(_07269_ ), .B(_06279_ ), .C1(\EX_LS_result_csreg_mem [13] ), .C2(_05315_ ), .ZN(_07270_ ) );
AND2_X1 _15297_ ( .A1(_07173_ ), .A2(_05143_ ), .ZN(_07271_ ) );
OR2_X1 _15298_ ( .A1(_07271_ ), .A2(_07171_ ), .ZN(_07272_ ) );
AND3_X1 _15299_ ( .A1(_07272_ ), .A2(_05145_ ), .A3(_07172_ ), .ZN(_07273_ ) );
AOI21_X1 _15300_ ( .A(_07172_ ), .B1(_07272_ ), .B2(_05145_ ), .ZN(_07274_ ) );
OR3_X1 _15301_ ( .A1(_07273_ ), .A2(_07274_ ), .A3(_07000_ ), .ZN(_07275_ ) );
AOI22_X1 _15302_ ( .A1(_05553_ ), .A2(_06824_ ), .B1(\ID_EX_imm [13] ), .B2(_06923_ ), .ZN(_07276_ ) );
AOI21_X1 _15303_ ( .A(_06542_ ), .B1(_07275_ ), .B2(_07276_ ), .ZN(_07277_ ) );
OR2_X1 _15304_ ( .A1(_07277_ ), .A2(_06932_ ), .ZN(_07278_ ) );
INV_X1 _15305_ ( .A(_07193_ ), .ZN(_07279_ ) );
AND2_X1 _15306_ ( .A1(_06985_ ), .A2(_06688_ ), .ZN(_07280_ ) );
INV_X1 _15307_ ( .A(_07280_ ), .ZN(_07281_ ) );
OAI211_X1 _15308_ ( .A(_06666_ ), .B(_07231_ ), .C1(_06675_ ), .C2(_06684_ ), .ZN(_07282_ ) );
AOI21_X1 _15309_ ( .A(_07279_ ), .B1(_07281_ ), .B2(_07282_ ), .ZN(_07283_ ) );
OAI21_X1 _15310_ ( .A(_06719_ ), .B1(_06749_ ), .B2(_06745_ ), .ZN(_07284_ ) );
OAI21_X1 _15311_ ( .A(_06683_ ), .B1(_06742_ ), .B2(_06772_ ), .ZN(_07285_ ) );
NAND3_X1 _15312_ ( .A1(_07284_ ), .A2(_06760_ ), .A3(_07285_ ), .ZN(_07286_ ) );
NAND3_X1 _15313_ ( .A1(_07091_ ), .A2(_07092_ ), .A3(_06790_ ), .ZN(_07287_ ) );
NAND3_X1 _15314_ ( .A1(_07286_ ), .A2(_07287_ ), .A3(_06795_ ), .ZN(_07288_ ) );
OAI211_X1 _15315_ ( .A(_06730_ ), .B(_07288_ ), .C1(_06726_ ), .C2(_07095_ ), .ZN(_07289_ ) );
NAND3_X1 _15316_ ( .A1(_06702_ ), .A2(_06792_ ), .A3(_07110_ ), .ZN(_07290_ ) );
NAND2_X1 _15317_ ( .A1(_07289_ ), .A2(_07290_ ), .ZN(_07291_ ) );
OAI21_X1 _15318_ ( .A(_06620_ ), .B1(_07283_ ), .B2(_07291_ ), .ZN(_07292_ ) );
NAND2_X1 _15319_ ( .A1(_07291_ ), .A2(_06907_ ), .ZN(_07293_ ) );
OR3_X1 _15320_ ( .A1(_06774_ ), .A2(_06766_ ), .A3(_06781_ ), .ZN(_07294_ ) );
NAND2_X1 _15321_ ( .A1(_06791_ ), .A2(_06800_ ), .ZN(_07295_ ) );
OAI21_X1 _15322_ ( .A(_07294_ ), .B1(_06796_ ), .B2(_07295_ ), .ZN(_07296_ ) );
NAND2_X1 _15323_ ( .A1(_07296_ ), .A2(_07250_ ), .ZN(_07297_ ) );
AOI22_X1 _15324_ ( .A1(_04973_ ), .A2(_07050_ ), .B1(_06593_ ), .B2(_07051_ ), .ZN(_07298_ ) );
AND4_X1 _15325_ ( .A1(_07292_ ), .A2(_07293_ ), .A3(_07297_ ), .A4(_07298_ ), .ZN(_07299_ ) );
AOI21_X1 _15326_ ( .A(_04979_ ), .B1(_07184_ ), .B2(_06587_ ), .ZN(_07300_ ) );
OR2_X1 _15327_ ( .A1(_07300_ ), .A2(_06594_ ), .ZN(_07301_ ) );
AOI21_X1 _15328_ ( .A(_06935_ ), .B1(_07301_ ), .B2(_04973_ ), .ZN(_07302_ ) );
OAI21_X1 _15329_ ( .A(_07302_ ), .B1(_04973_ ), .B2(_07301_ ), .ZN(_07303_ ) );
OAI21_X1 _15330_ ( .A(_06955_ ), .B1(_06631_ ), .B2(_02552_ ), .ZN(_07304_ ) );
NAND3_X1 _15331_ ( .A1(_07299_ ), .A2(_07303_ ), .A3(_07304_ ), .ZN(_07305_ ) );
AOI21_X1 _15332_ ( .A(_07278_ ), .B1(_07305_ ), .B2(_06816_ ), .ZN(_07306_ ) );
NAND2_X1 _15333_ ( .A1(_05556_ ), .A2(_05280_ ), .ZN(_07307_ ) );
NAND2_X1 _15334_ ( .A1(_07307_ ), .A2(_06249_ ), .ZN(_07308_ ) );
OAI21_X1 _15335_ ( .A(_07270_ ), .B1(_07306_ ), .B2(_07308_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
OR2_X1 _15336_ ( .A1(_05574_ ), .A2(_06921_ ), .ZN(_07309_ ) );
NAND3_X1 _15337_ ( .A1(_07173_ ), .A2(_07171_ ), .A3(_05143_ ), .ZN(_07310_ ) );
NAND3_X1 _15338_ ( .A1(_07272_ ), .A2(_06820_ ), .A3(_07310_ ), .ZN(_07311_ ) );
AOI22_X1 _15339_ ( .A1(_05563_ ), .A2(_06824_ ), .B1(\ID_EX_imm [12] ), .B2(_06923_ ), .ZN(_07312_ ) );
AOI21_X1 _15340_ ( .A(_06542_ ), .B1(_07311_ ), .B2(_07312_ ), .ZN(_07313_ ) );
OR2_X1 _15341_ ( .A1(_07313_ ), .A2(_05279_ ), .ZN(_07314_ ) );
NOR3_X1 _15342_ ( .A1(_06622_ ), .A2(_06763_ ), .A3(_07108_ ), .ZN(_07315_ ) );
INV_X1 _15343_ ( .A(_07315_ ), .ZN(_07316_ ) );
NAND4_X1 _15344_ ( .A1(_07084_ ), .A2(_06669_ ), .A3(_06667_ ), .A4(_07316_ ), .ZN(_07317_ ) );
OAI21_X1 _15345_ ( .A(_06750_ ), .B1(_07235_ ), .B2(_06890_ ), .ZN(_07318_ ) );
NOR2_X1 _15346_ ( .A1(_06679_ ), .A2(_02552_ ), .ZN(_07319_ ) );
OAI21_X1 _15347_ ( .A(_06746_ ), .B1(_07319_ ), .B2(_06879_ ), .ZN(_07320_ ) );
AOI21_X1 _15348_ ( .A(_06673_ ), .B1(_07318_ ), .B2(_07320_ ), .ZN(_07321_ ) );
AOI21_X1 _15349_ ( .A(_06723_ ), .B1(_07139_ ), .B2(_07140_ ), .ZN(_07322_ ) );
OAI21_X1 _15350_ ( .A(_06727_ ), .B1(_07321_ ), .B2(_07322_ ), .ZN(_07323_ ) );
OAI211_X1 _15351_ ( .A(_07323_ ), .B(_06729_ ), .C1(_06851_ ), .C2(_07038_ ), .ZN(_07324_ ) );
NAND3_X1 _15352_ ( .A1(_06858_ ), .A2(_05015_ ), .A3(_06795_ ), .ZN(_07325_ ) );
AND2_X1 _15353_ ( .A1(_07324_ ), .A2(_07325_ ), .ZN(_07326_ ) );
AOI21_X1 _15354_ ( .A(_06993_ ), .B1(_07317_ ), .B2(_07326_ ), .ZN(_07327_ ) );
AND3_X1 _15355_ ( .A1(_07184_ ), .A2(_04979_ ), .A3(_06587_ ), .ZN(_07328_ ) );
NOR3_X1 _15356_ ( .A1(_07328_ ), .A2(_07300_ ), .A3(_06934_ ), .ZN(_07329_ ) );
OR2_X1 _15357_ ( .A1(_07326_ ), .A2(_07208_ ), .ZN(_07330_ ) );
NOR2_X1 _15358_ ( .A1(_06873_ ), .A2(_07095_ ), .ZN(_07331_ ) );
AOI21_X1 _15359_ ( .A(_06763_ ), .B1(_06881_ ), .B2(_06888_ ), .ZN(_07332_ ) );
OAI21_X1 _15360_ ( .A(_07250_ ), .B1(_07331_ ), .B2(_07332_ ), .ZN(_07333_ ) );
NAND2_X1 _15361_ ( .A1(_04978_ ), .A2(_06913_ ), .ZN(_07334_ ) );
NAND3_X1 _15362_ ( .A1(_05073_ ), .A2(_02574_ ), .A3(_06983_ ), .ZN(_07335_ ) );
OAI21_X1 _15363_ ( .A(_04870_ ), .B1(_05073_ ), .B2(_02574_ ), .ZN(_07336_ ) );
AND3_X1 _15364_ ( .A1(_07334_ ), .A2(_07335_ ), .A3(_07336_ ), .ZN(_07337_ ) );
NAND3_X1 _15365_ ( .A1(_07330_ ), .A2(_07333_ ), .A3(_07337_ ), .ZN(_07338_ ) );
OR3_X1 _15366_ ( .A1(_07327_ ), .A2(_07329_ ), .A3(_07338_ ), .ZN(_07339_ ) );
BUF_X4 _15367_ ( .A(_06815_ ), .Z(_07340_ ) );
AOI21_X1 _15368_ ( .A(_07314_ ), .B1(_07339_ ), .B2(_07340_ ), .ZN(_07341_ ) );
OAI21_X1 _15369_ ( .A(_07061_ ), .B1(_05562_ ), .B2(_07062_ ), .ZN(_07342_ ) );
OAI21_X1 _15370_ ( .A(_07309_ ), .B1(_07341_ ), .B2(_07342_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
AOI22_X1 _15371_ ( .A1(_04044_ ), .A2(_06824_ ), .B1(\ID_EX_imm [30] ), .B2(_06923_ ), .ZN(_07343_ ) );
INV_X1 _15372_ ( .A(_04152_ ), .ZN(_07344_ ) );
NAND4_X1 _15373_ ( .A1(_05171_ ), .A2(_04226_ ), .A3(_04249_ ), .A4(_04271_ ), .ZN(_07345_ ) );
AND2_X1 _15374_ ( .A1(_07345_ ), .A2(_05181_ ), .ZN(_07346_ ) );
OR4_X1 _15375_ ( .A1(_07344_ ), .A2(_07346_ ), .A3(_04175_ ), .A4(_04174_ ), .ZN(_07347_ ) );
OAI21_X1 _15376_ ( .A(_07347_ ), .B1(_04174_ ), .B2(_05185_ ), .ZN(_07348_ ) );
AOI21_X1 _15377_ ( .A(_07000_ ), .B1(_07348_ ), .B2(_04103_ ), .ZN(_07349_ ) );
OAI21_X1 _15378_ ( .A(_07349_ ), .B1(_04103_ ), .B2(_07348_ ), .ZN(_07350_ ) );
AOI21_X1 _15379_ ( .A(_06542_ ), .B1(_07343_ ), .B2(_07350_ ), .ZN(_07351_ ) );
OR2_X1 _15380_ ( .A1(_07351_ ), .A2(_06932_ ), .ZN(_07352_ ) );
AND2_X1 _15381_ ( .A1(_05088_ ), .A2(_05092_ ), .ZN(_07353_ ) );
INV_X1 _15382_ ( .A(_07353_ ), .ZN(_07354_ ) );
INV_X2 _15383_ ( .A(_06910_ ), .ZN(_07355_ ) );
NOR3_X1 _15384_ ( .A1(_06545_ ), .A2(_04924_ ), .A3(_04923_ ), .ZN(_07356_ ) );
NAND4_X1 _15385_ ( .A1(_07355_ ), .A2(_04906_ ), .A3(_04913_ ), .A4(_07356_ ), .ZN(_07357_ ) );
AOI21_X1 _15386_ ( .A(_04924_ ), .B1(_04956_ ), .B2(_06614_ ), .ZN(_07358_ ) );
OR3_X1 _15387_ ( .A1(_07358_ ), .A2(_04907_ ), .A3(_04914_ ), .ZN(_07359_ ) );
OR2_X1 _15388_ ( .A1(_04905_ ), .A2(_02900_ ), .ZN(_07360_ ) );
NAND3_X1 _15389_ ( .A1(_02900_ ), .A2(_04904_ ), .A3(_04903_ ), .ZN(_07361_ ) );
NOR2_X1 _15390_ ( .A1(_04911_ ), .A2(_06501_ ), .ZN(_07362_ ) );
NAND3_X1 _15391_ ( .A1(_07360_ ), .A2(_07361_ ), .A3(_07362_ ), .ZN(_07363_ ) );
AND3_X1 _15392_ ( .A1(_07359_ ), .A2(_07360_ ), .A3(_07363_ ), .ZN(_07364_ ) );
AND2_X2 _15393_ ( .A1(_07357_ ), .A2(_07364_ ), .ZN(_07365_ ) );
INV_X1 _15394_ ( .A(_07365_ ), .ZN(_07366_ ) );
NAND3_X2 _15395_ ( .A1(_07366_ ), .A2(_05097_ ), .A3(_05102_ ), .ZN(_07367_ ) );
NOR2_X1 _15396_ ( .A1(_06470_ ), .A2(_05101_ ), .ZN(_07368_ ) );
NOR2_X1 _15397_ ( .A1(_05173_ ), .A2(_05096_ ), .ZN(_07369_ ) );
AOI21_X1 _15398_ ( .A(_07368_ ), .B1(_05102_ ), .B2(_07369_ ), .ZN(_07370_ ) );
AOI21_X2 _15399_ ( .A(_07354_ ), .B1(_07367_ ), .B2(_07370_ ), .ZN(_07371_ ) );
NOR2_X1 _15400_ ( .A1(_06837_ ), .A2(_05087_ ), .ZN(_07372_ ) );
AND3_X1 _15401_ ( .A1(_05087_ ), .A2(_02247_ ), .A3(_02246_ ), .ZN(_07373_ ) );
INV_X1 _15402_ ( .A(_07373_ ), .ZN(_07374_ ) );
INV_X1 _15403_ ( .A(_02965_ ), .ZN(_07375_ ) );
NOR2_X1 _15404_ ( .A1(_07375_ ), .A2(_05091_ ), .ZN(_07376_ ) );
AOI21_X1 _15405_ ( .A(_07372_ ), .B1(_07374_ ), .B2(_07376_ ), .ZN(_07377_ ) );
INV_X1 _15406_ ( .A(_07377_ ), .ZN(_07378_ ) );
OAI211_X2 _15407_ ( .A(_04895_ ), .B(_04900_ ), .C1(_07371_ ), .C2(_07378_ ), .ZN(_07379_ ) );
INV_X1 _15408_ ( .A(_04877_ ), .ZN(_07380_ ) );
AND2_X1 _15409_ ( .A1(_04893_ ), .A2(_02199_ ), .ZN(_07381_ ) );
AND2_X1 _15410_ ( .A1(_04899_ ), .A2(_02226_ ), .ZN(_07382_ ) );
AOI21_X1 _15411_ ( .A(_07381_ ), .B1(_07382_ ), .B2(_04895_ ), .ZN(_07383_ ) );
AND3_X1 _15412_ ( .A1(_07379_ ), .A2(_07380_ ), .A3(_07383_ ), .ZN(_07384_ ) );
AOI21_X1 _15413_ ( .A(_07380_ ), .B1(_07379_ ), .B2(_07383_ ), .ZN(_07385_ ) );
OR3_X2 _15414_ ( .A1(_07384_ ), .A2(_07385_ ), .A3(_06934_ ), .ZN(_07386_ ) );
OAI21_X1 _15415_ ( .A(_06683_ ), .B1(_06833_ ), .B2(_06839_ ), .ZN(_07387_ ) );
OAI21_X1 _15416_ ( .A(_06700_ ), .B1(_06846_ ), .B2(_06834_ ), .ZN(_07388_ ) );
AND3_X1 _15417_ ( .A1(_07387_ ), .A2(_07388_ ), .A3(_06703_ ), .ZN(_07389_ ) );
AND2_X1 _15418_ ( .A1(_06852_ ), .A2(_06838_ ), .ZN(_07390_ ) );
AOI21_X1 _15419_ ( .A(_06855_ ), .B1(_04894_ ), .B2(_06694_ ), .ZN(_07391_ ) );
MUX2_X1 _15420_ ( .A(_07390_ ), .B(_07391_ ), .S(_06715_ ), .Z(_07392_ ) );
AOI211_X1 _15421_ ( .A(_06762_ ), .B(_07389_ ), .C1(_07392_ ), .C2(_06760_ ), .ZN(_07393_ ) );
OAI21_X1 _15422_ ( .A(_06715_ ), .B1(_06843_ ), .B2(_06847_ ), .ZN(_07394_ ) );
OAI21_X1 _15423_ ( .A(_06719_ ), .B1(_06900_ ), .B2(_06844_ ), .ZN(_07395_ ) );
NAND2_X1 _15424_ ( .A1(_07394_ ), .A2(_07395_ ), .ZN(_07396_ ) );
NAND2_X1 _15425_ ( .A1(_07396_ ), .A2(_06872_ ), .ZN(_07397_ ) );
NAND3_X1 _15426_ ( .A1(_07026_ ), .A2(_06693_ ), .A3(_07027_ ), .ZN(_07398_ ) );
AOI21_X1 _15427_ ( .A(_06794_ ), .B1(_07397_ ), .B2(_07398_ ), .ZN(_07399_ ) );
OAI21_X1 _15428_ ( .A(_06734_ ), .B1(_07393_ ), .B2(_07399_ ), .ZN(_07400_ ) );
OR3_X1 _15429_ ( .A1(_07252_ ), .A2(_06627_ ), .A3(_07255_ ), .ZN(_07401_ ) );
AND3_X1 _15430_ ( .A1(_07400_ ), .A2(_07401_ ), .A3(_06739_ ), .ZN(_07402_ ) );
AND3_X1 _15431_ ( .A1(_06856_ ), .A2(_06849_ ), .A3(_06683_ ), .ZN(_07403_ ) );
NAND2_X1 _15432_ ( .A1(_07403_ ), .A2(_06727_ ), .ZN(_07404_ ) );
NOR2_X1 _15433_ ( .A1(_07404_ ), .A2(_05015_ ), .ZN(_07405_ ) );
AOI21_X1 _15434_ ( .A(_07405_ ), .B1(_07232_ ), .B2(_06670_ ), .ZN(_07406_ ) );
AOI21_X1 _15435_ ( .A(_06992_ ), .B1(_07406_ ), .B2(_07194_ ), .ZN(_07407_ ) );
AOI211_X1 _15436_ ( .A(_07402_ ), .B(_07407_ ), .C1(_06907_ ), .C2(_07405_ ), .ZN(_07408_ ) );
NAND2_X1 _15437_ ( .A1(_04877_ ), .A2(_06913_ ), .ZN(_07409_ ) );
OAI21_X1 _15438_ ( .A(_04870_ ), .B1(_05187_ ), .B2(_04876_ ), .ZN(_07410_ ) );
NAND3_X1 _15439_ ( .A1(_05187_ ), .A2(_04876_ ), .A3(_07051_ ), .ZN(_07411_ ) );
AND3_X1 _15440_ ( .A1(_07409_ ), .A2(_07410_ ), .A3(_07411_ ), .ZN(_07412_ ) );
AND2_X1 _15441_ ( .A1(_07408_ ), .A2(_07412_ ), .ZN(_07413_ ) );
AOI21_X1 _15442_ ( .A(_06814_ ), .B1(_07386_ ), .B2(_07413_ ), .ZN(_07414_ ) );
OAI221_X1 _15443_ ( .A(_06374_ ), .B1(_05343_ ), .B2(_03926_ ), .C1(_07352_ ), .C2(_07414_ ), .ZN(_07415_ ) );
NAND2_X1 _15444_ ( .A1(_05277_ ), .A2(_06372_ ), .ZN(_07416_ ) );
NAND2_X1 _15445_ ( .A1(_07415_ ), .A2(_07416_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
OR2_X1 _15446_ ( .A1(_05588_ ), .A2(_06921_ ), .ZN(_07417_ ) );
AND3_X1 _15447_ ( .A1(_05135_ ), .A2(_04550_ ), .A3(_04574_ ), .ZN(_07418_ ) );
OAI21_X1 _15448_ ( .A(_04504_ ), .B1(_07418_ ), .B2(_05142_ ), .ZN(_07419_ ) );
NAND2_X1 _15449_ ( .A1(_02647_ ), .A2(_04503_ ), .ZN(_07420_ ) );
AND2_X1 _15450_ ( .A1(_07419_ ), .A2(_07420_ ), .ZN(_07421_ ) );
XNOR2_X1 _15451_ ( .A(_07421_ ), .B(_04527_ ), .ZN(_07422_ ) );
NAND2_X1 _15452_ ( .A1(_07422_ ), .A2(_06537_ ), .ZN(_07423_ ) );
BUF_X4 _15453_ ( .A(_06525_ ), .Z(_07424_ ) );
AOI22_X1 _15454_ ( .A1(_05594_ ), .A2(_06823_ ), .B1(\ID_EX_imm [11] ), .B2(_07424_ ), .ZN(_07425_ ) );
AOI21_X1 _15455_ ( .A(_06542_ ), .B1(_07423_ ), .B2(_07425_ ), .ZN(_07426_ ) );
OR2_X1 _15456_ ( .A1(_07426_ ), .A2(_05279_ ), .ZN(_07427_ ) );
OAI211_X1 _15457_ ( .A(_06985_ ), .B(_07193_ ), .C1(_06689_ ), .C2(_06986_ ), .ZN(_07428_ ) );
AND3_X1 _15458_ ( .A1(_06952_ ), .A2(_06792_ ), .A3(_07095_ ), .ZN(_07429_ ) );
OAI21_X1 _15459_ ( .A(_06766_ ), .B1(_06943_ ), .B2(_06946_ ), .ZN(_07430_ ) );
NAND3_X1 _15460_ ( .A1(_07196_ ), .A2(_07197_ ), .A3(_06790_ ), .ZN(_07431_ ) );
OAI21_X1 _15461_ ( .A(_06747_ ), .B1(_06771_ ), .B2(_06769_ ), .ZN(_07432_ ) );
OAI21_X1 _15462_ ( .A(_06751_ ), .B1(_06742_ ), .B2(_06772_ ), .ZN(_07433_ ) );
NAND3_X1 _15463_ ( .A1(_07432_ ), .A2(_07433_ ), .A3(_06760_ ), .ZN(_07434_ ) );
NAND3_X1 _15464_ ( .A1(_07431_ ), .A2(_07434_ ), .A3(_06795_ ), .ZN(_07435_ ) );
AND3_X1 _15465_ ( .A1(_07430_ ), .A2(_06734_ ), .A3(_07435_ ), .ZN(_07436_ ) );
NOR2_X1 _15466_ ( .A1(_07429_ ), .A2(_07436_ ), .ZN(_07437_ ) );
AOI21_X1 _15467_ ( .A(_06993_ ), .B1(_07428_ ), .B2(_07437_ ), .ZN(_07438_ ) );
NOR2_X1 _15468_ ( .A1(_07437_ ), .A2(_07208_ ), .ZN(_07439_ ) );
INV_X1 _15469_ ( .A(_07217_ ), .ZN(_07440_ ) );
OR3_X1 _15470_ ( .A1(_06960_ ), .A2(_06795_ ), .A3(_07047_ ), .ZN(_07441_ ) );
NAND3_X1 _15471_ ( .A1(_06975_ ), .A2(_06979_ ), .A3(_06796_ ), .ZN(_07442_ ) );
AOI21_X1 _15472_ ( .A(_07440_ ), .B1(_07441_ ), .B2(_07442_ ), .ZN(_07443_ ) );
NAND3_X1 _15473_ ( .A1(_05069_ ), .A2(_02670_ ), .A3(_07051_ ), .ZN(_07444_ ) );
OAI21_X1 _15474_ ( .A(_07444_ ), .B1(_04985_ ), .B2(_05195_ ), .ZN(_07445_ ) );
NOR4_X1 _15475_ ( .A1(_07438_ ), .A2(_07439_ ), .A3(_07443_ ), .A4(_07445_ ), .ZN(_07446_ ) );
INV_X1 _15476_ ( .A(_06581_ ), .ZN(_07447_ ) );
OAI21_X1 _15477_ ( .A(_04989_ ), .B1(_06573_ ), .B2(_07447_ ), .ZN(_07448_ ) );
INV_X1 _15478_ ( .A(_06585_ ), .ZN(_07449_ ) );
AND3_X1 _15479_ ( .A1(_07448_ ), .A2(_04985_ ), .A3(_07449_ ), .ZN(_07450_ ) );
AOI21_X1 _15480_ ( .A(_04985_ ), .B1(_07448_ ), .B2(_07449_ ), .ZN(_07451_ ) );
OR3_X1 _15481_ ( .A1(_07450_ ), .A2(_07451_ ), .A3(_06935_ ), .ZN(_07452_ ) );
OAI21_X1 _15482_ ( .A(_06955_ ), .B1(_05069_ ), .B2(_02670_ ), .ZN(_07453_ ) );
NAND3_X1 _15483_ ( .A1(_07446_ ), .A2(_07452_ ), .A3(_07453_ ), .ZN(_07454_ ) );
AOI21_X1 _15484_ ( .A(_07427_ ), .B1(_07454_ ), .B2(_07340_ ), .ZN(_07455_ ) );
NAND2_X1 _15485_ ( .A1(_05597_ ), .A2(_05280_ ), .ZN(_07456_ ) );
NAND2_X1 _15486_ ( .A1(_07456_ ), .A2(_06249_ ), .ZN(_07457_ ) );
OAI21_X1 _15487_ ( .A(_07417_ ), .B1(_07455_ ), .B2(_07457_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OR2_X1 _15488_ ( .A1(_06352_ ), .A2(_06921_ ), .ZN(_07458_ ) );
OR3_X1 _15489_ ( .A1(_07418_ ), .A2(_04504_ ), .A3(_05142_ ), .ZN(_07459_ ) );
NAND3_X1 _15490_ ( .A1(_07459_ ), .A2(_06820_ ), .A3(_07419_ ), .ZN(_07460_ ) );
AOI22_X1 _15491_ ( .A1(_05629_ ), .A2(_06823_ ), .B1(\ID_EX_imm [10] ), .B2(_07424_ ), .ZN(_07461_ ) );
AOI21_X1 _15492_ ( .A(_06541_ ), .B1(_07460_ ), .B2(_07461_ ), .ZN(_07462_ ) );
OR2_X1 _15493_ ( .A1(_07462_ ), .A2(_05279_ ), .ZN(_07463_ ) );
AND4_X1 _15494_ ( .A1(_06677_ ), .A2(_06655_ ), .A3(_06675_ ), .A4(_07007_ ), .ZN(_07464_ ) );
OAI21_X1 _15495_ ( .A(_07193_ ), .B1(_07280_ ), .B2(_07464_ ), .ZN(_07465_ ) );
NAND3_X1 _15496_ ( .A1(_07022_ ), .A2(_05015_ ), .A3(_07038_ ), .ZN(_07466_ ) );
NAND3_X1 _15497_ ( .A1(_07236_ ), .A2(_07237_ ), .A3(_06693_ ), .ZN(_07467_ ) );
OAI21_X1 _15498_ ( .A(_06715_ ), .B1(_06878_ ), .B2(_06876_ ), .ZN(_07468_ ) );
OAI21_X1 _15499_ ( .A(_06719_ ), .B1(_07319_ ), .B2(_06879_ ), .ZN(_07469_ ) );
NAND3_X1 _15500_ ( .A1(_07468_ ), .A2(_07469_ ), .A3(_06724_ ), .ZN(_07470_ ) );
NAND3_X1 _15501_ ( .A1(_07467_ ), .A2(_07470_ ), .A3(_06794_ ), .ZN(_07471_ ) );
OAI211_X1 _15502_ ( .A(_06729_ ), .B(_07471_ ), .C1(_07016_ ), .C2(_06727_ ), .ZN(_07472_ ) );
AND2_X1 _15503_ ( .A1(_07466_ ), .A2(_07472_ ), .ZN(_07473_ ) );
AOI21_X1 _15504_ ( .A(_06993_ ), .B1(_07465_ ), .B2(_07473_ ), .ZN(_07474_ ) );
AOI21_X1 _15505_ ( .A(_07056_ ), .B1(_04988_ ), .B2(_06584_ ), .ZN(_07475_ ) );
OR3_X1 _15506_ ( .A1(_06573_ ), .A2(_04989_ ), .A3(_07447_ ), .ZN(_07476_ ) );
NAND3_X1 _15507_ ( .A1(_07476_ ), .A2(_06616_ ), .A3(_07448_ ), .ZN(_07477_ ) );
OR2_X1 _15508_ ( .A1(_07473_ ), .A2(_07208_ ), .ZN(_07478_ ) );
OAI21_X1 _15509_ ( .A(_07095_ ), .B1(_07037_ ), .B2(_07042_ ), .ZN(_07479_ ) );
OR3_X1 _15510_ ( .A1(_07046_ ), .A2(_07038_ ), .A3(_07108_ ), .ZN(_07480_ ) );
NAND2_X1 _15511_ ( .A1(_07479_ ), .A2(_07480_ ), .ZN(_07481_ ) );
NAND2_X1 _15512_ ( .A1(_07481_ ), .A2(_07250_ ), .ZN(_07482_ ) );
AOI22_X1 _15513_ ( .A1(_04989_ ), .A2(_06913_ ), .B1(_06585_ ), .B2(_07051_ ), .ZN(_07483_ ) );
NAND4_X1 _15514_ ( .A1(_07477_ ), .A2(_07478_ ), .A3(_07482_ ), .A4(_07483_ ), .ZN(_07484_ ) );
OR3_X1 _15515_ ( .A1(_07474_ ), .A2(_07475_ ), .A3(_07484_ ), .ZN(_07485_ ) );
AOI21_X1 _15516_ ( .A(_07463_ ), .B1(_07485_ ), .B2(_07340_ ), .ZN(_07486_ ) );
OAI21_X1 _15517_ ( .A(_07061_ ), .B1(_05627_ ), .B2(_07062_ ), .ZN(_07487_ ) );
OAI21_X1 _15518_ ( .A(_07458_ ), .B1(_07486_ ), .B2(_07487_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
OR2_X1 _15519_ ( .A1(_05652_ ), .A2(_06921_ ), .ZN(_07488_ ) );
AOI22_X1 _15520_ ( .A1(_05656_ ), .A2(_06824_ ), .B1(\ID_EX_imm [9] ), .B2(_06923_ ), .ZN(_07489_ ) );
AND2_X1 _15521_ ( .A1(_02600_ ), .A2(_04549_ ), .ZN(_07490_ ) );
AOI21_X1 _15522_ ( .A(_07490_ ), .B1(_05135_ ), .B2(_04550_ ), .ZN(_07491_ ) );
XNOR2_X1 _15523_ ( .A(_07491_ ), .B(_04574_ ), .ZN(_07492_ ) );
NAND2_X1 _15524_ ( .A1(_07492_ ), .A2(_06537_ ), .ZN(_07493_ ) );
AND2_X1 _15525_ ( .A1(_07489_ ), .A2(_07493_ ), .ZN(_07494_ ) );
OAI21_X1 _15526_ ( .A(_06518_ ), .B1(_07494_ ), .B2(_06543_ ), .ZN(_07495_ ) );
AND2_X1 _15527_ ( .A1(_07084_ ), .A2(_06689_ ), .ZN(_07496_ ) );
AND4_X1 _15528_ ( .A1(_06677_ ), .A2(_07083_ ), .A3(_06986_ ), .A4(_06684_ ), .ZN(_07497_ ) );
OAI21_X1 _15529_ ( .A(_07193_ ), .B1(_07496_ ), .B2(_07497_ ), .ZN(_07498_ ) );
NAND4_X1 _15530_ ( .A1(_07087_ ), .A2(_05015_ ), .A3(_06727_ ), .A4(_07088_ ), .ZN(_07499_ ) );
AOI21_X1 _15531_ ( .A(_06723_ ), .B1(_07284_ ), .B2(_07285_ ), .ZN(_07500_ ) );
OAI21_X1 _15532_ ( .A(_06683_ ), .B1(_06768_ ), .B2(_06776_ ), .ZN(_07501_ ) );
OAI21_X1 _15533_ ( .A(_06719_ ), .B1(_06771_ ), .B2(_06769_ ), .ZN(_07502_ ) );
AOI21_X1 _15534_ ( .A(_06703_ ), .B1(_07501_ ), .B2(_07502_ ), .ZN(_07503_ ) );
OAI21_X1 _15535_ ( .A(_06794_ ), .B1(_07500_ ), .B2(_07503_ ), .ZN(_07504_ ) );
OAI211_X1 _15536_ ( .A(_07504_ ), .B(_06729_ ), .C1(_06727_ ), .C2(_07094_ ), .ZN(_07505_ ) );
AND2_X1 _15537_ ( .A1(_07499_ ), .A2(_07505_ ), .ZN(_07506_ ) );
AOI21_X1 _15538_ ( .A(_06993_ ), .B1(_07498_ ), .B2(_07506_ ), .ZN(_07507_ ) );
AOI21_X1 _15539_ ( .A(_07056_ ), .B1(_04994_ ), .B2(_05062_ ), .ZN(_07508_ ) );
INV_X1 _15540_ ( .A(_04999_ ), .ZN(_07509_ ) );
AOI21_X1 _15541_ ( .A(_07509_ ), .B1(_06563_ ), .B2(_06572_ ), .ZN(_07510_ ) );
OR3_X1 _15542_ ( .A1(_07510_ ), .A2(_04995_ ), .A3(_06580_ ), .ZN(_07511_ ) );
OAI21_X1 _15543_ ( .A(_04995_ ), .B1(_07510_ ), .B2(_06580_ ), .ZN(_07512_ ) );
NAND3_X1 _15544_ ( .A1(_07511_ ), .A2(_06616_ ), .A3(_07512_ ), .ZN(_07513_ ) );
OR2_X1 _15545_ ( .A1(_07506_ ), .A2(_07208_ ), .ZN(_07514_ ) );
NAND3_X1 _15546_ ( .A1(_07102_ ), .A2(_07095_ ), .A3(_07105_ ), .ZN(_07515_ ) );
NAND4_X1 _15547_ ( .A1(_06959_ ), .A2(_06767_ ), .A3(_07158_ ), .A4(_07113_ ), .ZN(_07516_ ) );
NAND2_X1 _15548_ ( .A1(_07515_ ), .A2(_07516_ ), .ZN(_07517_ ) );
NAND2_X1 _15549_ ( .A1(_07517_ ), .A2(_07250_ ), .ZN(_07518_ ) );
AOI22_X1 _15550_ ( .A1(_04995_ ), .A2(_06913_ ), .B1(_05064_ ), .B2(_07051_ ), .ZN(_07519_ ) );
NAND4_X1 _15551_ ( .A1(_07513_ ), .A2(_07514_ ), .A3(_07518_ ), .A4(_07519_ ), .ZN(_07520_ ) );
OR3_X1 _15552_ ( .A1(_07507_ ), .A2(_07508_ ), .A3(_07520_ ), .ZN(_07521_ ) );
AOI21_X1 _15553_ ( .A(_07495_ ), .B1(_07521_ ), .B2(_07340_ ), .ZN(_07522_ ) );
NAND2_X1 _15554_ ( .A1(_05658_ ), .A2(_05280_ ), .ZN(_07523_ ) );
NAND2_X1 _15555_ ( .A1(_07523_ ), .A2(_06249_ ), .ZN(_07524_ ) );
OAI21_X1 _15556_ ( .A(_07488_ ), .B1(_07522_ ), .B2(_07524_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
OR2_X1 _15557_ ( .A1(_05674_ ), .A2(_06921_ ), .ZN(_07525_ ) );
AOI21_X1 _15558_ ( .A(_07000_ ), .B1(_05135_ ), .B2(_04550_ ), .ZN(_07526_ ) );
OAI21_X1 _15559_ ( .A(_07526_ ), .B1(_04550_ ), .B2(_05135_ ), .ZN(_07527_ ) );
AOI22_X1 _15560_ ( .A1(_05676_ ), .A2(_06823_ ), .B1(\ID_EX_imm [8] ), .B2(_07424_ ), .ZN(_07528_ ) );
AOI21_X1 _15561_ ( .A(_06541_ ), .B1(_07527_ ), .B2(_07528_ ), .ZN(_07529_ ) );
OR2_X1 _15562_ ( .A1(_07529_ ), .A2(_05279_ ), .ZN(_07530_ ) );
OAI211_X1 _15563_ ( .A(_06985_ ), .B(_07193_ ), .C1(_07103_ ), .C2(_06623_ ), .ZN(_07531_ ) );
NAND3_X1 _15564_ ( .A1(_07144_ ), .A2(_06793_ ), .A3(_06796_ ), .ZN(_07532_ ) );
NOR3_X1 _15565_ ( .A1(_06878_ ), .A2(_06746_ ), .A3(_06876_ ), .ZN(_07533_ ) );
NOR3_X1 _15566_ ( .A1(_06875_ ), .A2(_06699_ ), .A3(_06886_ ), .ZN(_07534_ ) );
NOR3_X1 _15567_ ( .A1(_07533_ ), .A2(_07534_ ), .A3(_06673_ ), .ZN(_07535_ ) );
AOI21_X1 _15568_ ( .A(_06723_ ), .B1(_07318_ ), .B2(_07320_ ), .ZN(_07536_ ) );
OAI21_X1 _15569_ ( .A(_06795_ ), .B1(_07535_ ), .B2(_07536_ ), .ZN(_07537_ ) );
OAI211_X1 _15570_ ( .A(_07537_ ), .B(_06730_ ), .C1(_07110_ ), .C2(_07142_ ), .ZN(_07538_ ) );
AND2_X1 _15571_ ( .A1(_07532_ ), .A2(_07538_ ), .ZN(_07539_ ) );
AOI21_X1 _15572_ ( .A(_06993_ ), .B1(_07531_ ), .B2(_07539_ ), .ZN(_07540_ ) );
AOI21_X1 _15573_ ( .A(_07208_ ), .B1(_07532_ ), .B2(_07538_ ), .ZN(_07541_ ) );
NAND3_X1 _15574_ ( .A1(_07157_ ), .A2(_07159_ ), .A3(_06796_ ), .ZN(_07542_ ) );
OR2_X1 _15575_ ( .A1(_07150_ ), .A2(_07095_ ), .ZN(_07543_ ) );
AND3_X1 _15576_ ( .A1(_07542_ ), .A2(_07250_ ), .A3(_07543_ ), .ZN(_07544_ ) );
NOR3_X1 _15577_ ( .A1(_07540_ ), .A2(_07541_ ), .A3(_07544_ ), .ZN(_07545_ ) );
AND3_X1 _15578_ ( .A1(_06563_ ), .A2(_07509_ ), .A3(_06572_ ), .ZN(_07546_ ) );
OR3_X1 _15579_ ( .A1(_07546_ ), .A2(_07510_ ), .A3(_06935_ ), .ZN(_07547_ ) );
AND2_X1 _15580_ ( .A1(_04999_ ), .A2(_07050_ ), .ZN(_07548_ ) );
NOR3_X1 _15581_ ( .A1(_04998_ ), .A2(_06579_ ), .A3(_07099_ ), .ZN(_07549_ ) );
AOI21_X1 _15582_ ( .A(_07056_ ), .B1(_04998_ ), .B2(_06579_ ), .ZN(_07550_ ) );
NOR3_X1 _15583_ ( .A1(_07548_ ), .A2(_07549_ ), .A3(_07550_ ), .ZN(_07551_ ) );
NAND3_X1 _15584_ ( .A1(_07545_ ), .A2(_07547_ ), .A3(_07551_ ), .ZN(_07552_ ) );
AOI21_X1 _15585_ ( .A(_07530_ ), .B1(_07552_ ), .B2(_07340_ ), .ZN(_07553_ ) );
NAND2_X1 _15586_ ( .A1(_05678_ ), .A2(_05280_ ), .ZN(_07554_ ) );
NAND2_X1 _15587_ ( .A1(_07554_ ), .A2(_06249_ ), .ZN(_07555_ ) );
OAI21_X1 _15588_ ( .A(_07525_ ), .B1(_07553_ ), .B2(_07555_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
NAND3_X1 _15589_ ( .A1(_05689_ ), .A2(_05690_ ), .A3(_06341_ ), .ZN(_07556_ ) );
OAI21_X1 _15590_ ( .A(_04838_ ), .B1(_05129_ ), .B2(_05133_ ), .ZN(_07557_ ) );
OAI21_X1 _15591_ ( .A(_07557_ ), .B1(_02870_ ), .B2(_04837_ ), .ZN(_07558_ ) );
AND2_X1 _15592_ ( .A1(_07558_ ), .A2(_04815_ ), .ZN(_07559_ ) );
OAI21_X1 _15593_ ( .A(_06536_ ), .B1(_07558_ ), .B2(_04815_ ), .ZN(_07560_ ) );
OR2_X1 _15594_ ( .A1(_07559_ ), .A2(_07560_ ), .ZN(_07561_ ) );
AOI22_X1 _15595_ ( .A1(_05694_ ), .A2(_06823_ ), .B1(\ID_EX_imm [7] ), .B2(_07424_ ), .ZN(_07562_ ) );
AOI21_X1 _15596_ ( .A(_06541_ ), .B1(_07561_ ), .B2(_07562_ ), .ZN(_07563_ ) );
OR2_X1 _15597_ ( .A1(_07563_ ), .A2(_05279_ ), .ZN(_07564_ ) );
NAND4_X1 _15598_ ( .A1(_06655_ ), .A2(_06689_ ), .A3(_06677_ ), .A4(_07193_ ), .ZN(_07565_ ) );
AND3_X1 _15599_ ( .A1(_06622_ ), .A2(_03005_ ), .A3(_06724_ ), .ZN(_07566_ ) );
MUX2_X1 _15600_ ( .A(_07566_ ), .B(_07202_ ), .S(_06794_ ), .Z(_07567_ ) );
OR2_X1 _15601_ ( .A1(_07567_ ), .A2(_06734_ ), .ZN(_07568_ ) );
AND3_X1 _15602_ ( .A1(_07432_ ), .A2(_07433_ ), .A3(_06790_ ), .ZN(_07569_ ) );
OAI21_X1 _15603_ ( .A(_06746_ ), .B1(_06775_ ), .B2(_06779_ ), .ZN(_07570_ ) );
OAI21_X1 _15604_ ( .A(_06700_ ), .B1(_06768_ ), .B2(_06776_ ), .ZN(_07571_ ) );
NAND2_X1 _15605_ ( .A1(_07570_ ), .A2(_07571_ ), .ZN(_07572_ ) );
INV_X1 _15606_ ( .A(_07572_ ), .ZN(_07573_ ) );
AOI211_X1 _15607_ ( .A(_06766_ ), .B(_07569_ ), .C1(_07573_ ), .C2(_07158_ ), .ZN(_07574_ ) );
NAND3_X1 _15608_ ( .A1(_07196_ ), .A2(_07197_ ), .A3(_06760_ ), .ZN(_07575_ ) );
AND3_X1 _15609_ ( .A1(_07195_ ), .A2(_06766_ ), .A3(_07575_ ), .ZN(_07576_ ) );
OAI21_X1 _15610_ ( .A(_06730_ ), .B1(_07574_ ), .B2(_07576_ ), .ZN(_07577_ ) );
NAND2_X1 _15611_ ( .A1(_07568_ ), .A2(_07577_ ), .ZN(_07578_ ) );
AOI21_X1 _15612_ ( .A(_06993_ ), .B1(_07565_ ), .B2(_07578_ ), .ZN(_07579_ ) );
AOI21_X1 _15613_ ( .A(_07056_ ), .B1(_05003_ ), .B2(_06370_ ), .ZN(_07580_ ) );
NAND3_X1 _15614_ ( .A1(_06558_ ), .A2(_06560_ ), .A3(_06562_ ), .ZN(_07581_ ) );
INV_X1 _15615_ ( .A(_06571_ ), .ZN(_07582_ ) );
AOI21_X1 _15616_ ( .A(_05010_ ), .B1(_07581_ ), .B2(_07582_ ), .ZN(_07583_ ) );
OR3_X1 _15617_ ( .A1(_07583_ ), .A2(_05004_ ), .A3(_06565_ ), .ZN(_07584_ ) );
OAI21_X1 _15618_ ( .A(_05004_ ), .B1(_07583_ ), .B2(_06565_ ), .ZN(_07585_ ) );
NAND3_X1 _15619_ ( .A1(_07584_ ), .A2(_06616_ ), .A3(_07585_ ), .ZN(_07586_ ) );
NAND3_X1 _15620_ ( .A1(_07568_ ), .A2(_06737_ ), .A3(_07577_ ), .ZN(_07587_ ) );
NOR3_X1 _15621_ ( .A1(_07211_ ), .A2(_06762_ ), .A3(_07440_ ), .ZN(_07588_ ) );
AOI221_X4 _15622_ ( .A(_07588_ ), .B1(_06564_ ), .B2(_06983_ ), .C1(_05004_ ), .C2(_05194_ ), .ZN(_07589_ ) );
NAND3_X1 _15623_ ( .A1(_07586_ ), .A2(_07587_ ), .A3(_07589_ ), .ZN(_07590_ ) );
OR3_X1 _15624_ ( .A1(_07579_ ), .A2(_07580_ ), .A3(_07590_ ), .ZN(_07591_ ) );
AOI21_X1 _15625_ ( .A(_07564_ ), .B1(_07591_ ), .B2(_07340_ ), .ZN(_07592_ ) );
NAND2_X1 _15626_ ( .A1(_05696_ ), .A2(_05280_ ), .ZN(_07593_ ) );
NAND2_X1 _15627_ ( .A1(_07593_ ), .A2(_06249_ ), .ZN(_07594_ ) );
OAI21_X1 _15628_ ( .A(_07556_ ), .B1(_07592_ ), .B2(_07594_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
NOR2_X1 _15629_ ( .A1(_05710_ ), .A2(_05206_ ), .ZN(_07595_ ) );
AND2_X1 _15630_ ( .A1(_07006_ ), .A2(_06872_ ), .ZN(_07596_ ) );
NOR4_X1 _15631_ ( .A1(_07230_ ), .A2(_07231_ ), .A3(_07279_ ), .A4(_07596_ ), .ZN(_07597_ ) );
MUX2_X1 _15632_ ( .A(_07403_ ), .B(_07242_ ), .S(_06625_ ), .Z(_07598_ ) );
NAND2_X1 _15633_ ( .A1(_07598_ ), .A2(_06792_ ), .ZN(_07599_ ) );
NAND3_X1 _15634_ ( .A1(_07234_ ), .A2(_07238_ ), .A3(_06766_ ), .ZN(_07600_ ) );
NOR3_X1 _15635_ ( .A1(_06885_ ), .A2(_06751_ ), .A3(_06883_ ), .ZN(_07601_ ) );
NOR3_X1 _15636_ ( .A1(_06875_ ), .A2(_06886_ ), .A3(_06747_ ), .ZN(_07602_ ) );
OAI21_X1 _15637_ ( .A(_06741_ ), .B1(_07601_ ), .B2(_07602_ ), .ZN(_07603_ ) );
NAND3_X1 _15638_ ( .A1(_07468_ ), .A2(_07469_ ), .A3(_07108_ ), .ZN(_07604_ ) );
NAND3_X1 _15639_ ( .A1(_07603_ ), .A2(_06795_ ), .A3(_07604_ ), .ZN(_07605_ ) );
NAND3_X1 _15640_ ( .A1(_07600_ ), .A2(_06734_ ), .A3(_07605_ ), .ZN(_07606_ ) );
NAND2_X1 _15641_ ( .A1(_07599_ ), .A2(_07606_ ), .ZN(_07607_ ) );
OAI21_X1 _15642_ ( .A(_06620_ ), .B1(_07597_ ), .B2(_07607_ ), .ZN(_07608_ ) );
AND3_X1 _15643_ ( .A1(_07581_ ), .A2(_05010_ ), .A3(_07582_ ), .ZN(_07609_ ) );
OR3_X1 _15644_ ( .A1(_07609_ ), .A2(_07583_ ), .A3(_06934_ ), .ZN(_07610_ ) );
NAND2_X1 _15645_ ( .A1(_07607_ ), .A2(_06737_ ), .ZN(_07611_ ) );
AND2_X1 _15646_ ( .A1(_07046_ ), .A2(_06673_ ), .ZN(_07612_ ) );
NOR3_X1 _15647_ ( .A1(_07612_ ), .A2(_07251_ ), .A3(_06762_ ), .ZN(_07613_ ) );
AND2_X1 _15648_ ( .A1(_07613_ ), .A2(_07217_ ), .ZN(_07614_ ) );
AOI221_X4 _15649_ ( .A(_07614_ ), .B1(_06565_ ), .B2(_06983_ ), .C1(_05009_ ), .C2(_05194_ ), .ZN(_07615_ ) );
NAND4_X1 _15650_ ( .A1(_07608_ ), .A2(_07610_ ), .A3(_07611_ ), .A4(_07615_ ), .ZN(_07616_ ) );
AOI21_X1 _15651_ ( .A(_07056_ ), .B1(_05008_ ), .B2(_02870_ ), .ZN(_07617_ ) );
OAI21_X1 _15652_ ( .A(_06815_ ), .B1(_07616_ ), .B2(_07617_ ), .ZN(_07618_ ) );
OR3_X1 _15653_ ( .A1(_05129_ ), .A2(_04838_ ), .A3(_05133_ ), .ZN(_07619_ ) );
NAND3_X1 _15654_ ( .A1(_07619_ ), .A2(_06820_ ), .A3(_07557_ ), .ZN(_07620_ ) );
AOI22_X1 _15655_ ( .A1(_05707_ ), .A2(_06823_ ), .B1(\ID_EX_imm [6] ), .B2(_07424_ ), .ZN(_07621_ ) );
AOI21_X1 _15656_ ( .A(_06541_ ), .B1(_07620_ ), .B2(_07621_ ), .ZN(_07622_ ) );
NOR2_X1 _15657_ ( .A1(_07622_ ), .A2(_05279_ ), .ZN(_07623_ ) );
AOI21_X1 _15658_ ( .A(_07595_ ), .B1(_07618_ ), .B2(_07623_ ), .ZN(_07624_ ) );
MUX2_X1 _15659_ ( .A(_05721_ ), .B(_07624_ ), .S(_06228_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _15660_ ( .A1(_05735_ ), .A2(_05737_ ), .ZN(_07625_ ) );
NAND2_X1 _15661_ ( .A1(_07625_ ), .A2(_06372_ ), .ZN(_07626_ ) );
AOI22_X1 _15662_ ( .A1(_05727_ ), .A2(_06823_ ), .B1(\ID_EX_imm [5] ), .B2(_07424_ ), .ZN(_07627_ ) );
AND2_X1 _15663_ ( .A1(_02864_ ), .A2(_04717_ ), .ZN(_07628_ ) );
AOI21_X1 _15664_ ( .A(_07628_ ), .B1(_05128_ ), .B2(_04719_ ), .ZN(_07629_ ) );
XOR2_X1 _15665_ ( .A(_07629_ ), .B(_04861_ ), .Z(_07630_ ) );
OAI21_X1 _15666_ ( .A(_07627_ ), .B1(_07630_ ), .B2(_07000_ ), .ZN(_07631_ ) );
AOI21_X1 _15667_ ( .A(_03885_ ), .B1(_07631_ ), .B2(_06540_ ), .ZN(_07632_ ) );
OAI21_X1 _15668_ ( .A(_06985_ ), .B1(_06986_ ), .B2(_06684_ ), .ZN(_07633_ ) );
NOR3_X1 _15669_ ( .A1(_07633_ ), .A2(_07231_ ), .A3(_07279_ ), .ZN(_07634_ ) );
NAND2_X1 _15670_ ( .A1(_06728_ ), .A2(_06792_ ), .ZN(_07635_ ) );
NAND3_X1 _15671_ ( .A1(_07286_ ), .A2(_07287_ ), .A3(_06766_ ), .ZN(_07636_ ) );
AND3_X1 _15672_ ( .A1(_07501_ ), .A2(_07502_ ), .A3(_06790_ ), .ZN(_07637_ ) );
OAI21_X1 _15673_ ( .A(_06747_ ), .B1(_06784_ ), .B2(_06778_ ), .ZN(_07638_ ) );
BUF_X4 _15674_ ( .A(_06719_ ), .Z(_07639_ ) );
OAI21_X1 _15675_ ( .A(_07639_ ), .B1(_06775_ ), .B2(_06779_ ), .ZN(_07640_ ) );
NAND2_X1 _15676_ ( .A1(_07638_ ), .A2(_07640_ ), .ZN(_07641_ ) );
OAI21_X1 _15677_ ( .A(_07038_ ), .B1(_07641_ ), .B2(_07108_ ), .ZN(_07642_ ) );
OAI211_X1 _15678_ ( .A(_07636_ ), .B(_06734_ ), .C1(_07637_ ), .C2(_07642_ ), .ZN(_07643_ ) );
NAND2_X1 _15679_ ( .A1(_07635_ ), .A2(_07643_ ), .ZN(_07644_ ) );
OAI21_X1 _15680_ ( .A(_06621_ ), .B1(_07634_ ), .B2(_07644_ ), .ZN(_07645_ ) );
NAND3_X1 _15681_ ( .A1(_06558_ ), .A2(_06560_ ), .A3(_05052_ ), .ZN(_07646_ ) );
NAND2_X1 _15682_ ( .A1(_07646_ ), .A2(_06570_ ), .ZN(_07647_ ) );
XNOR2_X1 _15683_ ( .A(_07647_ ), .B(_05019_ ), .ZN(_07648_ ) );
OR2_X1 _15684_ ( .A1(_07648_ ), .A2(_06934_ ), .ZN(_07649_ ) );
AOI21_X1 _15685_ ( .A(_07208_ ), .B1(_07635_ ), .B2(_07643_ ), .ZN(_07650_ ) );
NOR3_X1 _15686_ ( .A1(_06567_ ), .A2(_06566_ ), .A3(_05195_ ), .ZN(_07651_ ) );
OAI22_X1 _15687_ ( .A1(_06568_ ), .A2(_07099_ ), .B1(_06566_ ), .B2(_04871_ ), .ZN(_07652_ ) );
NOR3_X1 _15688_ ( .A1(_07295_ ), .A2(_06767_ ), .A3(_07440_ ), .ZN(_07653_ ) );
NOR4_X1 _15689_ ( .A1(_07650_ ), .A2(_07651_ ), .A3(_07652_ ), .A4(_07653_ ), .ZN(_07654_ ) );
AND3_X1 _15690_ ( .A1(_07645_ ), .A2(_07649_ ), .A3(_07654_ ), .ZN(_07655_ ) );
OAI21_X1 _15691_ ( .A(_07632_ ), .B1(_07655_ ), .B2(_06814_ ), .ZN(_07656_ ) );
OAI21_X1 _15692_ ( .A(_07656_ ), .B1(_05208_ ), .B2(_05725_ ), .ZN(_07657_ ) );
OAI21_X1 _15693_ ( .A(_07626_ ), .B1(_07657_ ), .B2(_06245_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
AND2_X1 _15694_ ( .A1(_05758_ ), .A2(_03885_ ), .ZN(_07658_ ) );
NAND3_X1 _15695_ ( .A1(_06830_ ), .A2(_06689_ ), .A3(_07193_ ), .ZN(_07659_ ) );
OR2_X1 _15696_ ( .A1(_06859_ ), .A2(_06729_ ), .ZN(_07660_ ) );
NOR3_X1 _15697_ ( .A1(_07533_ ), .A2(_07534_ ), .A3(_06723_ ), .ZN(_07661_ ) );
NOR3_X1 _15698_ ( .A1(_06885_ ), .A2(_06746_ ), .A3(_06883_ ), .ZN(_07662_ ) );
NOR3_X1 _15699_ ( .A1(_06882_ ), .A2(_06750_ ), .A3(_06869_ ), .ZN(_07663_ ) );
NOR2_X1 _15700_ ( .A1(_07662_ ), .A2(_07663_ ), .ZN(_07664_ ) );
AOI211_X1 _15701_ ( .A(_06762_ ), .B(_07661_ ), .C1(_06872_ ), .C2(_07664_ ), .ZN(_07665_ ) );
NOR3_X1 _15702_ ( .A1(_07321_ ), .A2(_07322_ ), .A3(_06625_ ), .ZN(_07666_ ) );
OR3_X1 _15703_ ( .A1(_07665_ ), .A2(_05015_ ), .A3(_07666_ ), .ZN(_07667_ ) );
NAND2_X1 _15704_ ( .A1(_07660_ ), .A2(_07667_ ), .ZN(_07668_ ) );
AOI21_X1 _15705_ ( .A(_06992_ ), .B1(_07659_ ), .B2(_07668_ ), .ZN(_07669_ ) );
NOR3_X1 _15706_ ( .A1(_06873_ ), .A2(_07103_ ), .A3(_07440_ ), .ZN(_07670_ ) );
NAND2_X1 _15707_ ( .A1(_05052_ ), .A2(_06913_ ), .ZN(_07671_ ) );
NAND3_X1 _15708_ ( .A1(_06792_ ), .A2(_02864_ ), .A3(_06983_ ), .ZN(_07672_ ) );
NAND2_X1 _15709_ ( .A1(_07671_ ), .A2(_07672_ ), .ZN(_07673_ ) );
OR3_X1 _15710_ ( .A1(_07669_ ), .A2(_07670_ ), .A3(_07673_ ), .ZN(_07674_ ) );
AOI21_X1 _15711_ ( .A(_05052_ ), .B1(_06558_ ), .B2(_06560_ ), .ZN(_07675_ ) );
NOR2_X1 _15712_ ( .A1(_07675_ ), .A2(_06934_ ), .ZN(_07676_ ) );
NAND2_X1 _15713_ ( .A1(_07676_ ), .A2(_07646_ ), .ZN(_07677_ ) );
OAI21_X1 _15714_ ( .A(_06955_ ), .B1(_06793_ ), .B2(_02864_ ), .ZN(_07678_ ) );
OAI211_X1 _15715_ ( .A(_07677_ ), .B(_07678_ ), .C1(_07668_ ), .C2(_07208_ ), .ZN(_07679_ ) );
OAI21_X1 _15716_ ( .A(_06815_ ), .B1(_07674_ ), .B2(_07679_ ), .ZN(_07680_ ) );
AOI21_X1 _15717_ ( .A(_07000_ ), .B1(_05128_ ), .B2(_04719_ ), .ZN(_07681_ ) );
OAI21_X1 _15718_ ( .A(_07681_ ), .B1(_04719_ ), .B2(_05128_ ), .ZN(_07682_ ) );
AOI22_X1 _15719_ ( .A1(_05756_ ), .A2(_06823_ ), .B1(\ID_EX_imm [4] ), .B2(_07424_ ), .ZN(_07683_ ) );
AOI21_X1 _15720_ ( .A(_06541_ ), .B1(_07682_ ), .B2(_07683_ ), .ZN(_07684_ ) );
NOR2_X1 _15721_ ( .A1(_07684_ ), .A2(_05279_ ), .ZN(_07685_ ) );
AOI21_X1 _15722_ ( .A(_07658_ ), .B1(_07680_ ), .B2(_07685_ ), .ZN(_07686_ ) );
MUX2_X1 _15723_ ( .A(_05754_ ), .B(_07686_ ), .S(_06228_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
INV_X1 _15724_ ( .A(_06401_ ), .ZN(_07687_ ) );
AND2_X1 _15725_ ( .A1(_05123_ ), .A2(_05125_ ), .ZN(_07688_ ) );
XNOR2_X1 _15726_ ( .A(_07688_ ), .B(_04696_ ), .ZN(_07689_ ) );
NAND2_X1 _15727_ ( .A1(_07689_ ), .A2(_06537_ ), .ZN(_07690_ ) );
AOI22_X1 _15728_ ( .A1(_05774_ ), .A2(_06823_ ), .B1(\ID_EX_imm [3] ), .B2(_07424_ ), .ZN(_07691_ ) );
AOI21_X1 _15729_ ( .A(_06541_ ), .B1(_07690_ ), .B2(_07691_ ), .ZN(_07692_ ) );
OR2_X1 _15730_ ( .A1(_07692_ ), .A2(_05279_ ), .ZN(_07693_ ) );
NAND4_X1 _15731_ ( .A1(_06985_ ), .A2(_06689_ ), .A3(_06986_ ), .A4(_07193_ ), .ZN(_07694_ ) );
NOR2_X1 _15732_ ( .A1(_06785_ ), .A2(_06788_ ), .ZN(_07695_ ) );
NOR2_X1 _15733_ ( .A1(_06784_ ), .A2(_06778_ ), .ZN(_07696_ ) );
MUX2_X1 _15734_ ( .A(_07695_ ), .B(_07696_ ), .S(_06700_ ), .Z(_07697_ ) );
MUX2_X1 _15735_ ( .A(_07573_ ), .B(_07697_ ), .S(_06724_ ), .Z(_07698_ ) );
AND2_X1 _15736_ ( .A1(_07698_ ), .A2(_07038_ ), .ZN(_07699_ ) );
AOI21_X1 _15737_ ( .A(_07038_ ), .B1(_07431_ ), .B2(_07434_ ), .ZN(_07700_ ) );
OR3_X1 _15738_ ( .A1(_07699_ ), .A2(_06792_ ), .A3(_07700_ ), .ZN(_07701_ ) );
OR2_X1 _15739_ ( .A1(_06953_ ), .A2(_06730_ ), .ZN(_07702_ ) );
NAND2_X1 _15740_ ( .A1(_07701_ ), .A2(_07702_ ), .ZN(_07703_ ) );
AOI21_X1 _15741_ ( .A(_06993_ ), .B1(_07694_ ), .B2(_07703_ ), .ZN(_07704_ ) );
AND3_X1 _15742_ ( .A1(_07701_ ), .A2(_06907_ ), .A3(_07702_ ), .ZN(_07705_ ) );
AND3_X1 _15743_ ( .A1(_06961_ ), .A2(_06794_ ), .A3(_07217_ ), .ZN(_07706_ ) );
AOI221_X4 _15744_ ( .A(_07706_ ), .B1(_06548_ ), .B2(_06983_ ), .C1(_05034_ ), .C2(_05194_ ), .ZN(_07707_ ) );
INV_X1 _15745_ ( .A(_06555_ ), .ZN(_07708_ ) );
INV_X1 _15746_ ( .A(_05041_ ), .ZN(_07709_ ) );
AOI21_X1 _15747_ ( .A(_06557_ ), .B1(_07708_ ), .B2(_07709_ ), .ZN(_07710_ ) );
INV_X1 _15748_ ( .A(_07710_ ), .ZN(_07711_ ) );
AOI21_X1 _15749_ ( .A(_05034_ ), .B1(_07711_ ), .B2(_06551_ ), .ZN(_07712_ ) );
NOR4_X1 _15750_ ( .A1(_07710_ ), .A2(_06548_ ), .A3(_06559_ ), .A4(_06550_ ), .ZN(_07713_ ) );
OAI21_X1 _15751_ ( .A(_06616_ ), .B1(_07712_ ), .B2(_07713_ ), .ZN(_07714_ ) );
OAI211_X1 _15752_ ( .A(_07707_ ), .B(_07714_ ), .C1(_06559_ ), .C2(_07056_ ), .ZN(_07715_ ) );
OR3_X1 _15753_ ( .A1(_07704_ ), .A2(_07705_ ), .A3(_07715_ ), .ZN(_07716_ ) );
AOI21_X1 _15754_ ( .A(_07693_ ), .B1(_07716_ ), .B2(_07340_ ), .ZN(_07717_ ) );
OAI21_X1 _15755_ ( .A(_07061_ ), .B1(_05208_ ), .B2(_05772_ ), .ZN(_07718_ ) );
OAI21_X1 _15756_ ( .A(_07687_ ), .B1(_07717_ ), .B2(_07718_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
INV_X1 _15757_ ( .A(_06412_ ), .ZN(_07719_ ) );
OR3_X1 _15758_ ( .A1(_04791_ ), .A2(_05122_ ), .A3(_04742_ ), .ZN(_07720_ ) );
NAND3_X1 _15759_ ( .A1(_07720_ ), .A2(_05123_ ), .A3(_06820_ ), .ZN(_07721_ ) );
AOI22_X1 _15760_ ( .A1(_05781_ ), .A2(_06823_ ), .B1(\ID_EX_imm [2] ), .B2(_07424_ ), .ZN(_07722_ ) );
AOI21_X1 _15761_ ( .A(_06541_ ), .B1(_07721_ ), .B2(_07722_ ), .ZN(_07723_ ) );
OR2_X1 _15762_ ( .A1(_07723_ ), .A2(_05279_ ), .ZN(_07724_ ) );
NAND3_X1 _15763_ ( .A1(_07084_ ), .A2(_06986_ ), .A3(_07007_ ), .ZN(_07725_ ) );
NOR3_X1 _15764_ ( .A1(_07725_ ), .A2(_07231_ ), .A3(_07279_ ), .ZN(_07726_ ) );
NAND2_X1 _15765_ ( .A1(_07023_ ), .A2(_06793_ ), .ZN(_07727_ ) );
OAI21_X1 _15766_ ( .A(_07047_ ), .B1(_07601_ ), .B2(_07602_ ), .ZN(_07728_ ) );
OAI21_X1 _15767_ ( .A(_07639_ ), .B1(_06882_ ), .B2(_06869_ ), .ZN(_07729_ ) );
NOR2_X1 _15768_ ( .A1(_06868_ ), .A2(_06866_ ), .ZN(_07730_ ) );
OAI211_X1 _15769_ ( .A(_07729_ ), .B(_07158_ ), .C1(_07730_ ), .C2(_07639_ ), .ZN(_07731_ ) );
AOI21_X1 _15770_ ( .A(_07103_ ), .B1(_07728_ ), .B2(_07731_ ), .ZN(_07732_ ) );
AOI21_X1 _15771_ ( .A(_06796_ ), .B1(_07467_ ), .B2(_07470_ ), .ZN(_07733_ ) );
OAI21_X1 _15772_ ( .A(_06731_ ), .B1(_07732_ ), .B2(_07733_ ), .ZN(_07734_ ) );
NAND2_X1 _15773_ ( .A1(_07727_ ), .A2(_07734_ ), .ZN(_07735_ ) );
OAI21_X1 _15774_ ( .A(_06621_ ), .B1(_07726_ ), .B2(_07735_ ), .ZN(_07736_ ) );
NAND2_X1 _15775_ ( .A1(_07735_ ), .A2(_06907_ ), .ZN(_07737_ ) );
AOI21_X1 _15776_ ( .A(_06934_ ), .B1(_06556_ ), .B2(_06557_ ), .ZN(_07738_ ) );
AND2_X1 _15777_ ( .A1(_07711_ ), .A2(_07738_ ), .ZN(_07739_ ) );
NOR4_X1 _15778_ ( .A1(_07046_ ), .A2(_06792_ ), .A3(_06767_ ), .A4(_07047_ ), .ZN(_07740_ ) );
AND2_X1 _15779_ ( .A1(_07740_ ), .A2(_06739_ ), .ZN(_07741_ ) );
AOI21_X1 _15780_ ( .A(_04871_ ), .B1(_07158_ ), .B2(_05047_ ), .ZN(_07742_ ) );
OAI22_X1 _15781_ ( .A1(_06557_ ), .A2(_05195_ ), .B1(_06551_ ), .B2(_07099_ ), .ZN(_07743_ ) );
NOR4_X1 _15782_ ( .A1(_07739_ ), .A2(_07741_ ), .A3(_07742_ ), .A4(_07743_ ), .ZN(_07744_ ) );
NAND3_X1 _15783_ ( .A1(_07736_ ), .A2(_07737_ ), .A3(_07744_ ), .ZN(_07745_ ) );
AOI21_X1 _15784_ ( .A(_07724_ ), .B1(_07745_ ), .B2(_07340_ ), .ZN(_07746_ ) );
OAI21_X1 _15785_ ( .A(_07061_ ), .B1(_05208_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07747_ ) );
OAI21_X1 _15786_ ( .A(_07719_ ), .B1(_07746_ ), .B2(_07747_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
NAND3_X1 _15787_ ( .A1(_05334_ ), .A2(_05339_ ), .A3(_06341_ ), .ZN(_07748_ ) );
OAI22_X1 _15788_ ( .A1(_05300_ ), .A2(_06523_ ), .B1(_02200_ ), .B2(_06527_ ), .ZN(_07749_ ) );
NOR2_X1 _15789_ ( .A1(_07346_ ), .A2(_07344_ ), .ZN(_07750_ ) );
AND2_X1 _15790_ ( .A1(_05184_ ), .A2(_02226_ ), .ZN(_07751_ ) );
OR3_X1 _15791_ ( .A1(_07750_ ), .A2(_07751_ ), .A3(_04176_ ), .ZN(_07752_ ) );
OAI21_X1 _15792_ ( .A(_04176_ ), .B1(_07750_ ), .B2(_07751_ ), .ZN(_07753_ ) );
AND3_X1 _15793_ ( .A1(_07752_ ), .A2(_06820_ ), .A3(_07753_ ), .ZN(_07754_ ) );
OAI21_X1 _15794_ ( .A(_06540_ ), .B1(_07749_ ), .B2(_07754_ ), .ZN(_07755_ ) );
NAND2_X1 _15795_ ( .A1(_07755_ ), .A2(_05343_ ), .ZN(_07756_ ) );
OAI21_X1 _15796_ ( .A(_04900_ ), .B1(_07371_ ), .B2(_07378_ ), .ZN(_07757_ ) );
INV_X1 _15797_ ( .A(_07757_ ), .ZN(_07758_ ) );
OAI21_X1 _15798_ ( .A(_04895_ ), .B1(_07758_ ), .B2(_07382_ ), .ZN(_07759_ ) );
OAI211_X1 _15799_ ( .A(_07757_ ), .B(_04896_ ), .C1(_02976_ ), .C2(_05116_ ), .ZN(_07760_ ) );
NAND3_X1 _15800_ ( .A1(_07759_ ), .A2(_06617_ ), .A3(_07760_ ), .ZN(_07761_ ) );
NAND2_X1 _15801_ ( .A1(_04895_ ), .A2(_07050_ ), .ZN(_07762_ ) );
NAND3_X1 _15802_ ( .A1(_04893_ ), .A2(_02199_ ), .A3(_07051_ ), .ZN(_07763_ ) );
OAI21_X1 _15803_ ( .A(_06955_ ), .B1(_04893_ ), .B2(_02199_ ), .ZN(_07764_ ) );
AND3_X1 _15804_ ( .A1(_07762_ ), .A2(_07763_ ), .A3(_07764_ ), .ZN(_07765_ ) );
NAND2_X1 _15805_ ( .A1(_06702_ ), .A2(_07038_ ), .ZN(_07766_ ) );
NOR2_X1 _15806_ ( .A1(_07766_ ), .A2(_05015_ ), .ZN(_07767_ ) );
OAI21_X1 _15807_ ( .A(_07282_ ), .B1(_07231_ ), .B2(_07230_ ), .ZN(_07768_ ) );
AOI21_X1 _15808_ ( .A(_07767_ ), .B1(_07768_ ), .B2(_06670_ ), .ZN(_07769_ ) );
AND2_X1 _15809_ ( .A1(_07084_ ), .A2(_06667_ ), .ZN(_07770_ ) );
AND2_X1 _15810_ ( .A1(_07770_ ), .A2(_06669_ ), .ZN(_07771_ ) );
INV_X1 _15811_ ( .A(_07771_ ), .ZN(_07772_ ) );
AOI21_X1 _15812_ ( .A(_06992_ ), .B1(_07769_ ), .B2(_07772_ ), .ZN(_07773_ ) );
AOI21_X1 _15813_ ( .A(_07773_ ), .B1(_06907_ ), .B2(_07767_ ), .ZN(_07774_ ) );
OAI21_X1 _15814_ ( .A(_06763_ ), .B1(_06754_ ), .B2(_06761_ ), .ZN(_07775_ ) );
NOR2_X1 _15815_ ( .A1(_06711_ ), .A2(_06708_ ), .ZN(_07776_ ) );
NAND2_X1 _15816_ ( .A1(_07776_ ), .A2(_07639_ ), .ZN(_07777_ ) );
OAI211_X1 _15817_ ( .A(_06696_ ), .B(_07113_ ), .C1(_02226_ ), .C2(_06680_ ), .ZN(_07778_ ) );
NAND3_X1 _15818_ ( .A1(_07777_ ), .A2(_06741_ ), .A3(_07778_ ), .ZN(_07779_ ) );
OR3_X1 _15819_ ( .A1(_06716_ ), .A2(_06747_ ), .A3(_06721_ ), .ZN(_07780_ ) );
OR3_X1 _15820_ ( .A1(_06720_ ), .A2(_06751_ ), .A3(_06712_ ), .ZN(_07781_ ) );
NAND2_X1 _15821_ ( .A1(_07780_ ), .A2(_07781_ ), .ZN(_07782_ ) );
OAI211_X1 _15822_ ( .A(_07779_ ), .B(_06795_ ), .C1(_07158_ ), .C2(_07782_ ), .ZN(_07783_ ) );
NAND3_X1 _15823_ ( .A1(_07775_ ), .A2(_07783_ ), .A3(_06730_ ), .ZN(_07784_ ) );
AND2_X1 _15824_ ( .A1(_07784_ ), .A2(_06739_ ), .ZN(_07785_ ) );
OAI21_X1 _15825_ ( .A(_07785_ ), .B1(_06731_ ), .B2(_07296_ ), .ZN(_07786_ ) );
AND2_X1 _15826_ ( .A1(_07774_ ), .A2(_07786_ ), .ZN(_07787_ ) );
NAND3_X1 _15827_ ( .A1(_07761_ ), .A2(_07765_ ), .A3(_07787_ ), .ZN(_07788_ ) );
AOI21_X1 _15828_ ( .A(_07756_ ), .B1(_07788_ ), .B2(_07340_ ), .ZN(_07789_ ) );
OAI21_X1 _15829_ ( .A(_07061_ ), .B1(_05295_ ), .B2(_07062_ ), .ZN(_07790_ ) );
OAI21_X1 _15830_ ( .A(_07748_ ), .B1(_07789_ ), .B2(_07790_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
OR2_X1 _15831_ ( .A1(_06429_ ), .A2(_06252_ ), .ZN(_07791_ ) );
NOR2_X1 _15832_ ( .A1(_04788_ ), .A2(_04790_ ), .ZN(_07792_ ) );
NOR3_X1 _15833_ ( .A1(_04791_ ), .A2(_07792_ ), .A3(_07000_ ), .ZN(_07793_ ) );
OAI22_X1 _15834_ ( .A1(_05798_ ), .A2(_06523_ ), .B1(_02718_ ), .B2(_06527_ ), .ZN(_07794_ ) );
OAI21_X1 _15835_ ( .A(_06540_ ), .B1(_07793_ ), .B2(_07794_ ), .ZN(_07795_ ) );
NAND2_X1 _15836_ ( .A1(_07795_ ), .A2(_05343_ ), .ZN(_07796_ ) );
NAND3_X1 _15837_ ( .A1(_06985_ ), .A2(_06986_ ), .A3(_06684_ ), .ZN(_07797_ ) );
NOR3_X1 _15838_ ( .A1(_07797_ ), .A2(_07231_ ), .A3(_07279_ ), .ZN(_07798_ ) );
NAND2_X1 _15839_ ( .A1(_07123_ ), .A2(_06793_ ), .ZN(_07799_ ) );
NAND3_X1 _15840_ ( .A1(_07638_ ), .A2(_07047_ ), .A3(_07640_ ), .ZN(_07800_ ) );
NOR3_X1 _15841_ ( .A1(_06787_ ), .A2(_07639_ ), .A3(_06798_ ), .ZN(_07801_ ) );
AOI21_X1 _15842_ ( .A(_07801_ ), .B1(_07639_ ), .B2(_07695_ ), .ZN(_07802_ ) );
OAI211_X1 _15843_ ( .A(_07110_ ), .B(_07800_ ), .C1(_07802_ ), .C2(_07047_ ), .ZN(_07803_ ) );
OAI21_X1 _15844_ ( .A(_07103_ ), .B1(_07500_ ), .B2(_07503_ ), .ZN(_07804_ ) );
NAND3_X1 _15845_ ( .A1(_07803_ ), .A2(_06735_ ), .A3(_07804_ ), .ZN(_07805_ ) );
NAND2_X1 _15846_ ( .A1(_07799_ ), .A2(_07805_ ), .ZN(_07806_ ) );
OAI21_X1 _15847_ ( .A(_06621_ ), .B1(_07798_ ), .B2(_07806_ ), .ZN(_07807_ ) );
XNOR2_X1 _15848_ ( .A(_07113_ ), .B(_02717_ ), .ZN(_07808_ ) );
INV_X1 _15849_ ( .A(_07808_ ), .ZN(_07809_ ) );
AOI21_X1 _15850_ ( .A(_06935_ ), .B1(_07809_ ), .B2(_06554_ ), .ZN(_07810_ ) );
NAND2_X1 _15851_ ( .A1(_07810_ ), .A2(_07708_ ), .ZN(_07811_ ) );
AOI21_X1 _15852_ ( .A(_07208_ ), .B1(_07799_ ), .B2(_07805_ ), .ZN(_07812_ ) );
AND3_X1 _15853_ ( .A1(_07114_ ), .A2(_06796_ ), .A3(_07250_ ), .ZN(_07813_ ) );
NOR3_X1 _15854_ ( .A1(_07113_ ), .A2(_05038_ ), .A3(_07099_ ), .ZN(_07814_ ) );
OAI22_X1 _15855_ ( .A1(_07809_ ), .A2(_05195_ ), .B1(_05039_ ), .B2(_04871_ ), .ZN(_07815_ ) );
NOR4_X1 _15856_ ( .A1(_07812_ ), .A2(_07813_ ), .A3(_07814_ ), .A4(_07815_ ), .ZN(_07816_ ) );
NAND3_X1 _15857_ ( .A1(_07807_ ), .A2(_07811_ ), .A3(_07816_ ), .ZN(_07817_ ) );
AOI21_X1 _15858_ ( .A(_07796_ ), .B1(_07817_ ), .B2(_07340_ ), .ZN(_07818_ ) );
OAI21_X1 _15859_ ( .A(_07061_ ), .B1(_05208_ ), .B2(\ID_EX_pc [1] ), .ZN(_07819_ ) );
OAI21_X1 _15860_ ( .A(_07791_ ), .B1(_07818_ ), .B2(_07819_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
OR2_X1 _15861_ ( .A1(_06435_ ), .A2(_06252_ ), .ZN(_07820_ ) );
INV_X1 _15862_ ( .A(_05115_ ), .ZN(_07821_ ) );
AOI221_X4 _15863_ ( .A(_04873_ ), .B1(_03005_ ), .B2(_04885_ ), .C1(_04890_ ), .C2(_05118_ ), .ZN(_07822_ ) );
AND3_X1 _15864_ ( .A1(_05112_ ), .A2(_07821_ ), .A3(_07822_ ), .ZN(_07823_ ) );
NAND4_X1 _15865_ ( .A1(_06655_ ), .A2(_05018_ ), .A3(_06628_ ), .A4(_06677_ ), .ZN(_07824_ ) );
OR2_X1 _15866_ ( .A1(_07145_ ), .A2(_06729_ ), .ZN(_07825_ ) );
OR3_X1 _15867_ ( .A1(_07535_ ), .A2(_06625_ ), .A3(_07536_ ), .ZN(_07826_ ) );
AND2_X1 _15868_ ( .A1(_06679_ ), .A2(_06552_ ), .ZN(_07827_ ) );
NOR3_X1 _15869_ ( .A1(_07827_ ), .A2(_06865_ ), .A3(_06750_ ), .ZN(_07828_ ) );
AOI21_X1 _15870_ ( .A(_07828_ ), .B1(_06751_ ), .B2(_07730_ ), .ZN(_07829_ ) );
MUX2_X1 _15871_ ( .A(_07664_ ), .B(_07829_ ), .S(_06724_ ), .Z(_07830_ ) );
OAI211_X1 _15872_ ( .A(_06729_ ), .B(_07826_ ), .C1(_07830_ ), .C2(_06762_ ), .ZN(_07831_ ) );
NAND2_X1 _15873_ ( .A1(_07825_ ), .A2(_07831_ ), .ZN(_07832_ ) );
AOI21_X1 _15874_ ( .A(_06992_ ), .B1(_07824_ ), .B2(_07832_ ), .ZN(_07833_ ) );
AND3_X1 _15875_ ( .A1(_07825_ ), .A2(_06736_ ), .A3(_07831_ ), .ZN(_07834_ ) );
AND3_X1 _15876_ ( .A1(_07150_ ), .A2(_06795_ ), .A3(_07217_ ), .ZN(_07835_ ) );
NOR4_X1 _15877_ ( .A1(_07823_ ), .A2(_07833_ ), .A3(_07834_ ), .A4(_07835_ ), .ZN(_07836_ ) );
OAI21_X1 _15878_ ( .A(_06617_ ), .B1(_06797_ ), .B2(_06862_ ), .ZN(_07837_ ) );
OAI21_X1 _15879_ ( .A(_06913_ ), .B1(_06797_ ), .B2(_06862_ ), .ZN(_07838_ ) );
NAND3_X1 _15880_ ( .A1(_06694_ ), .A2(_04743_ ), .A3(_06983_ ), .ZN(_07839_ ) );
OAI21_X1 _15881_ ( .A(_04870_ ), .B1(_06694_ ), .B2(_04743_ ), .ZN(_07840_ ) );
AND3_X1 _15882_ ( .A1(_07838_ ), .A2(_07839_ ), .A3(_07840_ ), .ZN(_07841_ ) );
AND3_X1 _15883_ ( .A1(_07836_ ), .A2(_07837_ ), .A3(_07841_ ), .ZN(_07842_ ) );
OAI21_X1 _15884_ ( .A(_05343_ ), .B1(_07842_ ), .B2(_06814_ ), .ZN(_07843_ ) );
AOI21_X1 _15885_ ( .A(_06809_ ), .B1(_04790_ ), .B2(_04765_ ), .ZN(_07844_ ) );
AOI221_X4 _15886_ ( .A(_07844_ ), .B1(\ID_EX_imm [0] ), .B2(_07424_ ), .C1(_05120_ ), .C2(_06812_ ), .ZN(_07845_ ) );
NAND3_X1 _15887_ ( .A1(_05830_ ), .A2(_06520_ ), .A3(_06519_ ), .ZN(_07846_ ) );
AOI21_X1 _15888_ ( .A(_06543_ ), .B1(_07845_ ), .B2(_07846_ ), .ZN(_07847_ ) );
OAI22_X1 _15889_ ( .A1(_07843_ ), .A2(_07847_ ), .B1(\ID_EX_pc [0] ), .B2(_05343_ ), .ZN(_07848_ ) );
OAI21_X1 _15890_ ( .A(_07820_ ), .B1(_07848_ ), .B2(_06372_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
NAND3_X1 _15891_ ( .A1(_05617_ ), .A2(_05620_ ), .A3(_06341_ ), .ZN(_07849_ ) );
OAI22_X1 _15892_ ( .A1(_05610_ ), .A2(_06523_ ), .B1(_06445_ ), .B2(_06527_ ), .ZN(_07850_ ) );
OAI21_X1 _15893_ ( .A(_06820_ ), .B1(_07346_ ), .B2(_07344_ ), .ZN(_07851_ ) );
AOI21_X1 _15894_ ( .A(_07851_ ), .B1(_07344_ ), .B2(_07346_ ), .ZN(_07852_ ) );
OAI21_X1 _15895_ ( .A(_06540_ ), .B1(_07850_ ), .B2(_07852_ ), .ZN(_07853_ ) );
NAND2_X1 _15896_ ( .A1(_07853_ ), .A2(_06518_ ), .ZN(_07854_ ) );
AND2_X1 _15897_ ( .A1(_07367_ ), .A2(_07370_ ), .ZN(_07855_ ) );
OAI211_X1 _15898_ ( .A(_04901_ ), .B(_07377_ ), .C1(_07855_ ), .C2(_07354_ ), .ZN(_07856_ ) );
NAND3_X1 _15899_ ( .A1(_07856_ ), .A2(_06617_ ), .A3(_07757_ ), .ZN(_07857_ ) );
NAND2_X1 _15900_ ( .A1(_04900_ ), .A2(_07050_ ), .ZN(_07858_ ) );
OAI21_X1 _15901_ ( .A(_06955_ ), .B1(_04899_ ), .B2(_02226_ ), .ZN(_07859_ ) );
NAND3_X1 _15902_ ( .A1(_04899_ ), .A2(_02226_ ), .A3(_07051_ ), .ZN(_07860_ ) );
AND3_X1 _15903_ ( .A1(_07858_ ), .A2(_07859_ ), .A3(_07860_ ), .ZN(_07861_ ) );
NOR2_X1 _15904_ ( .A1(_06833_ ), .A2(_06839_ ), .ZN(_07862_ ) );
MUX2_X1 _15905_ ( .A(_07862_ ), .B(_07390_ ), .S(_07113_ ), .Z(_07863_ ) );
NOR2_X1 _15906_ ( .A1(_07863_ ), .A2(_07108_ ), .ZN(_07864_ ) );
OAI21_X1 _15907_ ( .A(_07113_ ), .B1(_06846_ ), .B2(_06834_ ), .ZN(_07865_ ) );
OAI21_X1 _15908_ ( .A(_07639_ ), .B1(_06843_ ), .B2(_06847_ ), .ZN(_07866_ ) );
AOI21_X1 _15909_ ( .A(_06741_ ), .B1(_07865_ ), .B2(_07866_ ), .ZN(_07867_ ) );
OAI21_X1 _15910_ ( .A(_07095_ ), .B1(_07864_ ), .B2(_07867_ ), .ZN(_07868_ ) );
OAI211_X1 _15911_ ( .A(_07868_ ), .B(_06765_ ), .C1(_06796_ ), .C2(_06903_ ), .ZN(_07869_ ) );
OAI21_X1 _15912_ ( .A(_06793_ ), .B1(_07331_ ), .B2(_07332_ ), .ZN(_07870_ ) );
AOI21_X1 _15913_ ( .A(_06740_ ), .B1(_07869_ ), .B2(_07870_ ), .ZN(_07871_ ) );
NOR3_X1 _15914_ ( .A1(_06857_ ), .A2(_06767_ ), .A3(_07047_ ), .ZN(_07872_ ) );
AND3_X1 _15915_ ( .A1(_07872_ ), .A2(_06765_ ), .A3(_06737_ ), .ZN(_07873_ ) );
NAND2_X1 _15916_ ( .A1(_07872_ ), .A2(_06735_ ), .ZN(_07874_ ) );
NAND4_X1 _15917_ ( .A1(_07083_ ), .A2(_06677_ ), .A3(_06670_ ), .A4(_07316_ ), .ZN(_07875_ ) );
INV_X1 _15918_ ( .A(_07770_ ), .ZN(_07876_ ) );
OAI211_X1 _15919_ ( .A(_07874_ ), .B(_07875_ ), .C1(_07876_ ), .C2(_06691_ ), .ZN(_07877_ ) );
AOI211_X1 _15920_ ( .A(_07871_ ), .B(_07873_ ), .C1(_07877_ ), .C2(_06621_ ), .ZN(_07878_ ) );
NAND3_X1 _15921_ ( .A1(_07857_ ), .A2(_07861_ ), .A3(_07878_ ), .ZN(_07879_ ) );
AOI21_X1 _15922_ ( .A(_07854_ ), .B1(_07879_ ), .B2(_06815_ ), .ZN(_07880_ ) );
OAI21_X1 _15923_ ( .A(_07061_ ), .B1(_05608_ ), .B2(_07062_ ), .ZN(_07881_ ) );
OAI21_X1 _15924_ ( .A(_07849_ ), .B1(_07880_ ), .B2(_07881_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
OAI211_X1 _15925_ ( .A(_06452_ ), .B(_06279_ ), .C1(\EX_LS_result_csreg_mem [27] ), .C2(_05315_ ), .ZN(_07882_ ) );
OAI22_X1 _15926_ ( .A1(_05817_ ), .A2(_06523_ ), .B1(_02249_ ), .B2(_06527_ ), .ZN(_07883_ ) );
AND3_X1 _15927_ ( .A1(_05171_ ), .A2(_04249_ ), .A3(_04271_ ), .ZN(_07884_ ) );
OR3_X1 _15928_ ( .A1(_07884_ ), .A2(_05177_ ), .A3(_05175_ ), .ZN(_07885_ ) );
AND2_X1 _15929_ ( .A1(_07885_ ), .A2(_04225_ ), .ZN(_07886_ ) );
AOI21_X1 _15930_ ( .A(_07886_ ), .B1(_02965_ ), .B2(_05179_ ), .ZN(_07887_ ) );
XNOR2_X1 _15931_ ( .A(_07887_ ), .B(_04203_ ), .ZN(_07888_ ) );
AOI21_X1 _15932_ ( .A(_07883_ ), .B1(_07888_ ), .B2(_06537_ ), .ZN(_07889_ ) );
OAI21_X1 _15933_ ( .A(_06518_ ), .B1(_07889_ ), .B2(_06543_ ), .ZN(_07890_ ) );
INV_X1 _15934_ ( .A(_05092_ ), .ZN(_07891_ ) );
AOI21_X1 _15935_ ( .A(_07891_ ), .B1(_07367_ ), .B2(_07370_ ), .ZN(_07892_ ) );
OR3_X1 _15936_ ( .A1(_07892_ ), .A2(_05088_ ), .A3(_07376_ ), .ZN(_07893_ ) );
OAI21_X1 _15937_ ( .A(_05088_ ), .B1(_07892_ ), .B2(_07376_ ), .ZN(_07894_ ) );
NAND3_X1 _15938_ ( .A1(_07893_ ), .A2(_06617_ ), .A3(_07894_ ), .ZN(_07895_ ) );
AOI211_X1 _15939_ ( .A(_06765_ ), .B(_06740_ ), .C1(_07441_ ), .C2(_07442_ ), .ZN(_07896_ ) );
OAI21_X1 _15940_ ( .A(_06747_ ), .B1(_06716_ ), .B2(_06721_ ), .ZN(_07897_ ) );
OAI21_X1 _15941_ ( .A(_07639_ ), .B1(_06755_ ), .B2(_06717_ ), .ZN(_07898_ ) );
AND3_X1 _15942_ ( .A1(_07897_ ), .A2(_07898_ ), .A3(_07108_ ), .ZN(_07899_ ) );
OAI21_X1 _15943_ ( .A(_07113_ ), .B1(_06711_ ), .B2(_06708_ ), .ZN(_07900_ ) );
OAI21_X1 _15944_ ( .A(_07639_ ), .B1(_06720_ ), .B2(_06712_ ), .ZN(_07901_ ) );
AND2_X1 _15945_ ( .A1(_07900_ ), .A2(_07901_ ), .ZN(_07902_ ) );
AOI211_X1 _15946_ ( .A(_06767_ ), .B(_07899_ ), .C1(_07158_ ), .C2(_07902_ ), .ZN(_07903_ ) );
AOI211_X1 _15947_ ( .A(_07440_ ), .B(_07903_ ), .C1(_07103_ ), .C2(_06972_ ), .ZN(_07904_ ) );
AOI211_X1 _15948_ ( .A(_07896_ ), .B(_07904_ ), .C1(_07374_ ), .C2(_06955_ ), .ZN(_07905_ ) );
AND2_X1 _15949_ ( .A1(_06952_ ), .A2(_07095_ ), .ZN(_07906_ ) );
AOI21_X1 _15950_ ( .A(_06990_ ), .B1(_06735_ ), .B2(_07906_ ), .ZN(_07907_ ) );
OAI211_X1 _15951_ ( .A(_07084_ ), .B(_06670_ ), .C1(_06689_ ), .C2(_06986_ ), .ZN(_07908_ ) );
AOI21_X1 _15952_ ( .A(_06992_ ), .B1(_07907_ ), .B2(_07908_ ), .ZN(_07909_ ) );
AND3_X1 _15953_ ( .A1(_07906_ ), .A2(_06735_ ), .A3(_06737_ ), .ZN(_07910_ ) );
NOR3_X1 _15954_ ( .A1(_07372_ ), .A2(_07373_ ), .A3(_05195_ ), .ZN(_07911_ ) );
NOR3_X1 _15955_ ( .A1(_06837_ ), .A2(_05087_ ), .A3(_07099_ ), .ZN(_07912_ ) );
NOR4_X1 _15956_ ( .A1(_07909_ ), .A2(_07910_ ), .A3(_07911_ ), .A4(_07912_ ), .ZN(_07913_ ) );
NAND3_X1 _15957_ ( .A1(_07895_ ), .A2(_07905_ ), .A3(_07913_ ), .ZN(_07914_ ) );
AOI21_X1 _15958_ ( .A(_07890_ ), .B1(_07914_ ), .B2(_06815_ ), .ZN(_07915_ ) );
OAI21_X1 _15959_ ( .A(_06237_ ), .B1(_05812_ ), .B2(_07062_ ), .ZN(_07916_ ) );
OAI21_X1 _15960_ ( .A(_07882_ ), .B1(_07915_ ), .B2(_07916_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
OR2_X1 _15961_ ( .A1(_06465_ ), .A2(_06252_ ), .ZN(_07917_ ) );
OAI22_X1 _15962_ ( .A1(_05849_ ), .A2(_06523_ ), .B1(_02966_ ), .B2(_06527_ ), .ZN(_07918_ ) );
NOR2_X1 _15963_ ( .A1(_07885_ ), .A2(_04225_ ), .ZN(_07919_ ) );
NOR3_X1 _15964_ ( .A1(_07886_ ), .A2(_07919_ ), .A3(_07000_ ), .ZN(_07920_ ) );
OAI21_X1 _15965_ ( .A(_06540_ ), .B1(_07918_ ), .B2(_07920_ ), .ZN(_07921_ ) );
NAND2_X1 _15966_ ( .A1(_07921_ ), .A2(_06518_ ), .ZN(_07922_ ) );
OAI21_X1 _15967_ ( .A(_06617_ ), .B1(_07855_ ), .B2(_07891_ ), .ZN(_07923_ ) );
AOI21_X1 _15968_ ( .A(_07923_ ), .B1(_07891_ ), .B2(_07855_ ), .ZN(_07924_ ) );
NOR2_X1 _15969_ ( .A1(_07021_ ), .A2(_06766_ ), .ZN(_07925_ ) );
AOI21_X1 _15970_ ( .A(_06990_ ), .B1(_06735_ ), .B2(_07925_ ), .ZN(_07926_ ) );
OAI21_X1 _15971_ ( .A(_06670_ ), .B1(_07280_ ), .B2(_07464_ ), .ZN(_07927_ ) );
AOI21_X1 _15972_ ( .A(_06993_ ), .B1(_07926_ ), .B2(_07927_ ), .ZN(_07928_ ) );
NAND2_X1 _15973_ ( .A1(_05092_ ), .A2(_06913_ ), .ZN(_07929_ ) );
NAND3_X1 _15974_ ( .A1(_07925_ ), .A2(_06734_ ), .A3(_06737_ ), .ZN(_07930_ ) );
NAND2_X1 _15975_ ( .A1(_07376_ ), .A2(_06983_ ), .ZN(_07931_ ) );
AOI21_X1 _15976_ ( .A(_02965_ ), .B1(_05089_ ), .B2(_05090_ ), .ZN(_07932_ ) );
OR2_X1 _15977_ ( .A1(_07932_ ), .A2(_04871_ ), .ZN(_07933_ ) );
AND4_X1 _15978_ ( .A1(_07929_ ), .A2(_07930_ ), .A3(_07931_ ), .A4(_07933_ ), .ZN(_07934_ ) );
NOR2_X1 _15979_ ( .A1(_06734_ ), .A2(_06740_ ), .ZN(_07935_ ) );
NAND2_X1 _15980_ ( .A1(_07481_ ), .A2(_07935_ ), .ZN(_07936_ ) );
OR2_X1 _15981_ ( .A1(_07032_ ), .A2(_07095_ ), .ZN(_07937_ ) );
NAND3_X1 _15982_ ( .A1(_07387_ ), .A2(_07388_ ), .A3(_07158_ ), .ZN(_07938_ ) );
OAI211_X1 _15983_ ( .A(_07938_ ), .B(_06796_ ), .C1(_07396_ ), .C2(_07158_ ), .ZN(_07939_ ) );
NAND3_X1 _15984_ ( .A1(_07937_ ), .A2(_07250_ ), .A3(_07939_ ), .ZN(_07940_ ) );
NAND3_X1 _15985_ ( .A1(_07934_ ), .A2(_07936_ ), .A3(_07940_ ), .ZN(_07941_ ) );
OR3_X1 _15986_ ( .A1(_07924_ ), .A2(_07928_ ), .A3(_07941_ ), .ZN(_07942_ ) );
AOI21_X1 _15987_ ( .A(_07922_ ), .B1(_07942_ ), .B2(_06815_ ), .ZN(_07943_ ) );
NAND2_X1 _15988_ ( .A1(_05846_ ), .A2(_06932_ ), .ZN(_07944_ ) );
NAND2_X1 _15989_ ( .A1(_07944_ ), .A2(_06249_ ), .ZN(_07945_ ) );
OAI21_X1 _15990_ ( .A(_07917_ ), .B1(_07943_ ), .B2(_07945_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
NAND3_X1 _15991_ ( .A1(_06474_ ), .A2(_06475_ ), .A3(_06341_ ), .ZN(_07946_ ) );
OAI22_X1 _15992_ ( .A1(_05871_ ), .A2(_06523_ ), .B1(_02968_ ), .B2(_06527_ ), .ZN(_07947_ ) );
AOI21_X1 _15993_ ( .A(_05174_ ), .B1(_05171_ ), .B2(_04271_ ), .ZN(_07948_ ) );
XNOR2_X1 _15994_ ( .A(_07948_ ), .B(_04249_ ), .ZN(_07949_ ) );
AOI21_X1 _15995_ ( .A(_07947_ ), .B1(_07949_ ), .B2(_06537_ ), .ZN(_07950_ ) );
OAI21_X1 _15996_ ( .A(_06518_ ), .B1(_07950_ ), .B2(_06543_ ), .ZN(_07951_ ) );
AOI21_X1 _15997_ ( .A(_05098_ ), .B1(_07357_ ), .B2(_07364_ ), .ZN(_07952_ ) );
OR3_X1 _15998_ ( .A1(_07952_ ), .A2(_07369_ ), .A3(_05103_ ), .ZN(_07953_ ) );
OAI21_X1 _15999_ ( .A(_05103_ ), .B1(_07952_ ), .B2(_07369_ ), .ZN(_07954_ ) );
AOI21_X1 _16000_ ( .A(_06935_ ), .B1(_07953_ ), .B2(_07954_ ), .ZN(_07955_ ) );
NAND2_X1 _16001_ ( .A1(_07517_ ), .A2(_07935_ ), .ZN(_07956_ ) );
NAND2_X1 _16002_ ( .A1(_07782_ ), .A2(_07158_ ), .ZN(_07957_ ) );
NAND3_X1 _16003_ ( .A1(_06756_ ), .A2(_06759_ ), .A3(_07047_ ), .ZN(_07958_ ) );
AOI21_X1 _16004_ ( .A(_06767_ ), .B1(_07957_ ), .B2(_07958_ ), .ZN(_07959_ ) );
AND3_X1 _16005_ ( .A1(_07107_ ), .A2(_07109_ ), .A3(_06763_ ), .ZN(_07960_ ) );
OAI21_X1 _16006_ ( .A(_07250_ ), .B1(_07959_ ), .B2(_07960_ ), .ZN(_00304_ ) );
AOI21_X1 _16007_ ( .A(_02940_ ), .B1(_05099_ ), .B2(_05100_ ), .ZN(_00305_ ) );
OAI211_X1 _16008_ ( .A(_07956_ ), .B(_00304_ ), .C1(_00305_ ), .C2(_07056_ ), .ZN(_00306_ ) );
NAND4_X1 _16009_ ( .A1(_06985_ ), .A2(_07231_ ), .A3(_06986_ ), .A4(_06684_ ), .ZN(_00307_ ) );
AOI21_X1 _16010_ ( .A(_06671_ ), .B1(_07281_ ), .B2(_00307_ ), .ZN(_00308_ ) );
AND3_X1 _16011_ ( .A1(_07087_ ), .A2(_06625_ ), .A3(_07088_ ), .ZN(_00309_ ) );
AND2_X1 _16012_ ( .A1(_00309_ ), .A2(_06729_ ), .ZN(_00310_ ) );
OR2_X1 _16013_ ( .A1(_06990_ ), .A2(_00310_ ), .ZN(_00311_ ) );
OAI21_X1 _16014_ ( .A(_06620_ ), .B1(_00308_ ), .B2(_00311_ ), .ZN(_00312_ ) );
NAND3_X1 _16015_ ( .A1(_00309_ ), .A2(_06735_ ), .A3(_06737_ ), .ZN(_00313_ ) );
AOI22_X1 _16016_ ( .A1(_05102_ ), .A2(_06913_ ), .B1(_07368_ ), .B2(_07051_ ), .ZN(_00314_ ) );
NAND3_X1 _16017_ ( .A1(_00312_ ), .A2(_00313_ ), .A3(_00314_ ), .ZN(_00315_ ) );
OR3_X1 _16018_ ( .A1(_07955_ ), .A2(_00306_ ), .A3(_00315_ ), .ZN(_00316_ ) );
AOI21_X1 _16019_ ( .A(_07951_ ), .B1(_00316_ ), .B2(_06815_ ), .ZN(_00317_ ) );
OAI21_X1 _16020_ ( .A(_06237_ ), .B1(_05867_ ), .B2(_07062_ ), .ZN(_00318_ ) );
OAI21_X1 _16021_ ( .A(_07946_ ), .B1(_00317_ ), .B2(_00318_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _16022_ ( .A1(_06488_ ), .A2(_06372_ ), .ZN(_00319_ ) );
OAI22_X1 _16023_ ( .A1(_05890_ ), .A2(_06523_ ), .B1(_02272_ ), .B2(_06527_ ), .ZN(_00320_ ) );
OR2_X1 _16024_ ( .A1(_05171_ ), .A2(_04271_ ), .ZN(_00321_ ) );
AOI21_X1 _16025_ ( .A(_07000_ ), .B1(_05171_ ), .B2(_04271_ ), .ZN(_00322_ ) );
AOI21_X1 _16026_ ( .A(_00320_ ), .B1(_00321_ ), .B2(_00322_ ), .ZN(_00323_ ) );
OAI21_X1 _16027_ ( .A(_06518_ ), .B1(_00323_ ), .B2(_06543_ ), .ZN(_00324_ ) );
NOR2_X1 _16028_ ( .A1(_07952_ ), .A2(_06935_ ), .ZN(_00325_ ) );
OAI21_X1 _16029_ ( .A(_00325_ ), .B1(_05097_ ), .B2(_07366_ ), .ZN(_00326_ ) );
NAND2_X1 _16030_ ( .A1(_07144_ ), .A2(_07110_ ), .ZN(_00327_ ) );
OAI211_X1 _16031_ ( .A(_06655_ ), .B(_06677_ ), .C1(_07103_ ), .C2(_06623_ ), .ZN(_00328_ ) );
OAI221_X1 _16032_ ( .A(_07194_ ), .B1(_06793_ ), .B2(_00327_ ), .C1(_06671_ ), .C2(_00328_ ), .ZN(_00329_ ) );
NAND2_X1 _16033_ ( .A1(_00329_ ), .A2(_06621_ ), .ZN(_00330_ ) );
AOI21_X1 _16034_ ( .A(_02271_ ), .B1(_05094_ ), .B2(_05095_ ), .ZN(_00331_ ) );
OR2_X1 _16035_ ( .A1(_00331_ ), .A2(_04871_ ), .ZN(_00332_ ) );
NOR3_X1 _16036_ ( .A1(_00327_ ), .A2(_06793_ ), .A3(_07208_ ), .ZN(_00333_ ) );
NAND2_X1 _16037_ ( .A1(_07155_ ), .A2(_06767_ ), .ZN(_00334_ ) );
AOI21_X1 _16038_ ( .A(_07108_ ), .B1(_07865_ ), .B2(_07866_ ), .ZN(_00335_ ) );
AOI21_X1 _16039_ ( .A(_06741_ ), .B1(_06899_ ), .B2(_06901_ ), .ZN(_00336_ ) );
OAI21_X1 _16040_ ( .A(_06795_ ), .B1(_00335_ ), .B2(_00336_ ), .ZN(_00337_ ) );
AND3_X1 _16041_ ( .A1(_00334_ ), .A2(_07250_ ), .A3(_00337_ ), .ZN(_00338_ ) );
NOR2_X1 _16042_ ( .A1(_00333_ ), .A2(_00338_ ), .ZN(_00339_ ) );
AOI22_X1 _16043_ ( .A1(_05097_ ), .A2(_07050_ ), .B1(_07369_ ), .B2(_07051_ ), .ZN(_00340_ ) );
NAND3_X1 _16044_ ( .A1(_07542_ ), .A2(_07543_ ), .A3(_07935_ ), .ZN(_00341_ ) );
AND4_X1 _16045_ ( .A1(_00332_ ), .A2(_00339_ ), .A3(_00340_ ), .A4(_00341_ ), .ZN(_00342_ ) );
NAND3_X1 _16046_ ( .A1(_00326_ ), .A2(_00330_ ), .A3(_00342_ ), .ZN(_00343_ ) );
AOI21_X1 _16047_ ( .A(_00324_ ), .B1(_00343_ ), .B2(_06815_ ), .ZN(_00344_ ) );
OAI21_X1 _16048_ ( .A(_06237_ ), .B1(_05887_ ), .B2(_07062_ ), .ZN(_00345_ ) );
OAI21_X1 _16049_ ( .A(_00319_ ), .B1(_00344_ ), .B2(_00345_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
INV_X1 _16050_ ( .A(_06497_ ), .ZN(_00346_ ) );
OAI22_X1 _16051_ ( .A1(_05912_ ), .A2(_06522_ ), .B1(_02308_ ), .B2(_06527_ ), .ZN(_00347_ ) );
OAI21_X1 _16052_ ( .A(_05166_ ), .B1(_06533_ ), .B2(_04479_ ), .ZN(_00348_ ) );
AOI21_X1 _16053_ ( .A(_05162_ ), .B1(_00348_ ), .B2(_04430_ ), .ZN(_00349_ ) );
XNOR2_X1 _16054_ ( .A(_00349_ ), .B(_04407_ ), .ZN(_00350_ ) );
AOI21_X1 _16055_ ( .A(_00347_ ), .B1(_00350_ ), .B2(_06537_ ), .ZN(_00351_ ) );
OAI21_X1 _16056_ ( .A(_06518_ ), .B1(_00351_ ), .B2(_06543_ ), .ZN(_00352_ ) );
NAND2_X1 _16057_ ( .A1(_07355_ ), .A2(_07356_ ), .ZN(_00353_ ) );
AOI21_X1 _16058_ ( .A(_04914_ ), .B1(_00353_ ), .B2(_07358_ ), .ZN(_00354_ ) );
OAI21_X1 _16059_ ( .A(_04906_ ), .B1(_00354_ ), .B2(_07362_ ), .ZN(_00355_ ) );
NAND2_X1 _16060_ ( .A1(_00355_ ), .A2(_06617_ ), .ZN(_00356_ ) );
NOR3_X1 _16061_ ( .A1(_00354_ ), .A2(_04906_ ), .A3(_07362_ ), .ZN(_00357_ ) );
OR2_X1 _16062_ ( .A1(_00356_ ), .A2(_00357_ ), .ZN(_00358_ ) );
NAND3_X1 _16063_ ( .A1(_07360_ ), .A2(_07361_ ), .A3(_07050_ ), .ZN(_00359_ ) );
NAND2_X1 _16064_ ( .A1(_07361_ ), .A2(_06955_ ), .ZN(_00360_ ) );
OR3_X1 _16065_ ( .A1(_04905_ ), .A2(_02900_ ), .A3(_07099_ ), .ZN(_00361_ ) );
AND3_X1 _16066_ ( .A1(_00359_ ), .A2(_00360_ ), .A3(_00361_ ), .ZN(_00362_ ) );
AOI21_X1 _16067_ ( .A(_06668_ ), .B1(_06765_ ), .B2(_07231_ ), .ZN(_00363_ ) );
AND2_X1 _16068_ ( .A1(_07567_ ), .A2(_06730_ ), .ZN(_00364_ ) );
OAI21_X1 _16069_ ( .A(_06621_ ), .B1(_00363_ ), .B2(_00364_ ), .ZN(_00365_ ) );
NAND2_X1 _16070_ ( .A1(_06966_ ), .A2(_07108_ ), .ZN(_00366_ ) );
NAND2_X1 _16071_ ( .A1(_07897_ ), .A2(_07898_ ), .ZN(_00367_ ) );
NAND2_X1 _16072_ ( .A1(_00367_ ), .A2(_06741_ ), .ZN(_00368_ ) );
AOI21_X1 _16073_ ( .A(_06763_ ), .B1(_00366_ ), .B2(_00368_ ), .ZN(_00369_ ) );
AOI211_X1 _16074_ ( .A(_06792_ ), .B(_00369_ ), .C1(_07103_ ), .C2(_07215_ ), .ZN(_00370_ ) );
NOR3_X1 _16075_ ( .A1(_07211_ ), .A2(_06765_ ), .A3(_07103_ ), .ZN(_00371_ ) );
OAI21_X1 _16076_ ( .A(_06739_ ), .B1(_00370_ ), .B2(_00371_ ), .ZN(_00372_ ) );
NAND3_X1 _16077_ ( .A1(_07567_ ), .A2(_06731_ ), .A3(_06907_ ), .ZN(_00373_ ) );
AND3_X1 _16078_ ( .A1(_00365_ ), .A2(_00372_ ), .A3(_00373_ ), .ZN(_00374_ ) );
NAND3_X1 _16079_ ( .A1(_00358_ ), .A2(_00362_ ), .A3(_00374_ ), .ZN(_00375_ ) );
AOI21_X1 _16080_ ( .A(_00352_ ), .B1(_06816_ ), .B2(_00375_ ), .ZN(_00376_ ) );
OAI21_X1 _16081_ ( .A(_06237_ ), .B1(_05905_ ), .B2(_05343_ ), .ZN(_00377_ ) );
OAI21_X1 _16082_ ( .A(_00346_ ), .B1(_00376_ ), .B2(_00377_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _16083_ ( .A1(_05940_ ), .A2(_06372_ ), .ZN(_00378_ ) );
OAI22_X1 _16084_ ( .A1(_05929_ ), .A2(_06522_ ), .B1(_02334_ ), .B2(_06526_ ), .ZN(_00379_ ) );
OR2_X1 _16085_ ( .A1(_00348_ ), .A2(_04430_ ), .ZN(_00380_ ) );
AOI21_X1 _16086_ ( .A(_07000_ ), .B1(_00348_ ), .B2(_04430_ ), .ZN(_00381_ ) );
AOI21_X1 _16087_ ( .A(_00379_ ), .B1(_00380_ ), .B2(_00381_ ), .ZN(_00382_ ) );
OAI21_X1 _16088_ ( .A(_06518_ ), .B1(_00382_ ), .B2(_06543_ ), .ZN(_00383_ ) );
AND3_X1 _16089_ ( .A1(_00353_ ), .A2(_04914_ ), .A3(_07358_ ), .ZN(_00384_ ) );
OR3_X1 _16090_ ( .A1(_00384_ ), .A2(_00354_ ), .A3(_06935_ ), .ZN(_00385_ ) );
OAI21_X1 _16091_ ( .A(_06739_ ), .B1(_07613_ ), .B2(_06731_ ), .ZN(_00386_ ) );
NOR3_X1 _16092_ ( .A1(_07253_ ), .A2(_07254_ ), .A3(_06796_ ), .ZN(_00387_ ) );
AND3_X1 _16093_ ( .A1(_07397_ ), .A2(_07398_ ), .A3(_07110_ ), .ZN(_00388_ ) );
NOR3_X1 _16094_ ( .A1(_00387_ ), .A2(_00388_ ), .A3(_06793_ ), .ZN(_00389_ ) );
OR2_X1 _16095_ ( .A1(_00386_ ), .A2(_00389_ ), .ZN(_00390_ ) );
NOR4_X1 _16096_ ( .A1(_07230_ ), .A2(_07231_ ), .A3(_06671_ ), .A4(_07596_ ), .ZN(_00391_ ) );
AND2_X1 _16097_ ( .A1(_07598_ ), .A2(_06729_ ), .ZN(_00392_ ) );
OR3_X1 _16098_ ( .A1(_00391_ ), .A2(_06990_ ), .A3(_00392_ ), .ZN(_00393_ ) );
NAND2_X1 _16099_ ( .A1(_00393_ ), .A2(_06621_ ), .ZN(_00394_ ) );
NAND3_X1 _16100_ ( .A1(_07598_ ), .A2(_06731_ ), .A3(_06907_ ), .ZN(_00395_ ) );
OR3_X1 _16101_ ( .A1(_04911_ ), .A2(_06501_ ), .A3(_07099_ ), .ZN(_00396_ ) );
AOI21_X1 _16102_ ( .A(_04871_ ), .B1(_04911_ ), .B2(_06501_ ), .ZN(_00397_ ) );
AOI21_X1 _16103_ ( .A(_00397_ ), .B1(_04913_ ), .B2(_07050_ ), .ZN(_00398_ ) );
AND4_X1 _16104_ ( .A1(_00394_ ), .A2(_00395_ ), .A3(_00396_ ), .A4(_00398_ ), .ZN(_00399_ ) );
NAND3_X1 _16105_ ( .A1(_00385_ ), .A2(_00390_ ), .A3(_00399_ ), .ZN(_00400_ ) );
AOI21_X1 _16106_ ( .A(_00383_ ), .B1(_00400_ ), .B2(_06815_ ), .ZN(_00401_ ) );
NAND2_X1 _16107_ ( .A1(_05927_ ), .A2(_06932_ ), .ZN(_00402_ ) );
NAND2_X1 _16108_ ( .A1(_00402_ ), .A2(_06374_ ), .ZN(_00403_ ) );
OAI21_X1 _16109_ ( .A(_00378_ ), .B1(_00401_ ), .B2(_00403_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NOR3_X1 _16110_ ( .A1(_05981_ ), .A2(_05982_ ), .A3(_06252_ ), .ZN(_00404_ ) );
INV_X1 _16111_ ( .A(_00404_ ), .ZN(_00405_ ) );
NOR2_X1 _16112_ ( .A1(_02172_ ), .A2(_04101_ ), .ZN(_00406_ ) );
AOI21_X1 _16113_ ( .A(_00406_ ), .B1(_07348_ ), .B2(_04103_ ), .ZN(_00407_ ) );
XNOR2_X1 _16114_ ( .A(_00407_ ), .B(_04128_ ), .ZN(_00408_ ) );
AOI22_X1 _16115_ ( .A1(_00408_ ), .A2(_06537_ ), .B1(\ID_EX_imm [31] ), .B2(_06923_ ), .ZN(_00409_ ) );
OR2_X1 _16116_ ( .A1(_05974_ ), .A2(_06523_ ), .ZN(_00410_ ) );
AOI21_X1 _16117_ ( .A(_06543_ ), .B1(_00409_ ), .B2(_00410_ ), .ZN(_00411_ ) );
AND2_X1 _16118_ ( .A1(_05187_ ), .A2(_04876_ ), .ZN(_00412_ ) );
OR3_X2 _16119_ ( .A1(_07385_ ), .A2(_04889_ ), .A3(_00412_ ), .ZN(_00413_ ) );
OAI21_X1 _16120_ ( .A(_04889_ ), .B1(_07385_ ), .B2(_00412_ ), .ZN(_00414_ ) );
NAND3_X1 _16121_ ( .A1(_00413_ ), .A2(_06617_ ), .A3(_00414_ ), .ZN(_00415_ ) );
NAND2_X1 _16122_ ( .A1(_06628_ ), .A2(_03005_ ), .ZN(_00416_ ) );
AOI21_X1 _16123_ ( .A(_06992_ ), .B1(_06668_ ), .B2(_00416_ ), .ZN(_00417_ ) );
OAI211_X1 _16124_ ( .A(_06695_ ), .B(_07113_ ), .C1(_03005_ ), .C2(_06694_ ), .ZN(_00418_ ) );
OAI211_X1 _16125_ ( .A(_06696_ ), .B(_07639_ ), .C1(_02226_ ), .C2(_06680_ ), .ZN(_00419_ ) );
AOI21_X1 _16126_ ( .A(_07108_ ), .B1(_00418_ ), .B2(_00419_ ), .ZN(_00420_ ) );
AOI211_X1 _16127_ ( .A(_06767_ ), .B(_00420_ ), .C1(_07047_ ), .C2(_07902_ ), .ZN(_00421_ ) );
AOI21_X1 _16128_ ( .A(_07110_ ), .B1(_00366_ ), .B2(_00368_ ), .ZN(_00422_ ) );
NOR3_X1 _16129_ ( .A1(_00421_ ), .A2(_07440_ ), .A3(_00422_ ), .ZN(_00423_ ) );
AND3_X1 _16130_ ( .A1(_07212_ ), .A2(_07216_ ), .A3(_07935_ ), .ZN(_00424_ ) );
AND3_X1 _16131_ ( .A1(_06628_ ), .A2(_03005_ ), .A3(_06736_ ), .ZN(_00425_ ) );
AOI221_X4 _16132_ ( .A(_00425_ ), .B1(_04886_ ), .B2(_04870_ ), .C1(_04889_ ), .C2(_05194_ ), .ZN(_00426_ ) );
OR2_X1 _16133_ ( .A1(_04887_ ), .A2(_06804_ ), .ZN(_00427_ ) );
NAND2_X1 _16134_ ( .A1(_00426_ ), .A2(_00427_ ), .ZN(_00428_ ) );
NOR4_X1 _16135_ ( .A1(_00417_ ), .A2(_00423_ ), .A3(_00424_ ), .A4(_00428_ ), .ZN(_00429_ ) );
AOI21_X1 _16136_ ( .A(_06814_ ), .B1(_00415_ ), .B2(_00429_ ), .ZN(_00430_ ) );
NOR3_X1 _16137_ ( .A1(_00411_ ), .A2(_00430_ ), .A3(_05280_ ), .ZN(_00431_ ) );
NAND2_X1 _16138_ ( .A1(_05968_ ), .A2(_06932_ ), .ZN(_00432_ ) );
NAND2_X1 _16139_ ( .A1(_00432_ ), .A2(_06374_ ), .ZN(_00433_ ) );
OAI21_X1 _16140_ ( .A(_00405_ ), .B1(_00431_ ), .B2(_00433_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
AND3_X1 _16141_ ( .A1(\myexu.state_$_ANDNOT__B_Y ), .A2(_03902_ ), .A3(_03904_ ), .ZN(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ) );
AND2_X1 _16142_ ( .A1(_06206_ ), .A2(_02093_ ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16143_ ( .A(IDU_ready_IFU ), .ZN(_00434_ ) );
NAND2_X1 _16144_ ( .A1(_00434_ ), .A2(IDU_valid_EXU ), .ZN(_00435_ ) );
OAI21_X1 _16145_ ( .A(_00435_ ), .B1(_03323_ ), .B2(_03219_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16146_ ( .A1(_03296_ ), .A2(_03219_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16147_ ( .A1(_03296_ ), .A2(_03219_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16148_ ( .A(_03216_ ), .ZN(_00436_ ) );
NOR4_X1 _16149_ ( .A1(_03296_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03091_ ), .A4(_00436_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16150_ ( .A1(_03618_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03091_ ), .A4(_03215_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16151_ ( .A(_03834_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16152_ ( .A(_00435_ ), .B1(_00436_ ), .B2(_00434_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16153_ ( .A(\myidu.state [2] ), .ZN(_00437_ ) );
OAI22_X1 _16154_ ( .A1(_03323_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B1(_00437_ ), .B2(loaduse_clear ), .ZN(_00438_ ) );
AOI221_X4 _16155_ ( .A(_00438_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .C1(IDU_ready_IFU ), .C2(_00436_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16156_ ( .A(_03291_ ), .ZN(_00439_ ) );
OAI21_X1 _16157_ ( .A(_03345_ ), .B1(_00439_ ), .B2(_03083_ ), .ZN(_00440_ ) );
OAI21_X1 _16158_ ( .A(_03355_ ), .B1(_03232_ ), .B2(_03273_ ), .ZN(_00441_ ) );
NAND4_X1 _16159_ ( .A1(_03217_ ), .A2(_00440_ ), .A3(_03151_ ), .A4(_00441_ ), .ZN(_00442_ ) );
NAND3_X1 _16160_ ( .A1(_03151_ ), .A2(IDU_valid_EXU ), .A3(_06009_ ), .ZN(_00443_ ) );
NAND2_X1 _16161_ ( .A1(_00208_ ), .A2(loaduse_clear ), .ZN(_00444_ ) );
NAND3_X1 _16162_ ( .A1(_00442_ ), .A2(_00443_ ), .A3(_00444_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16163_ ( .A(_03151_ ), .B(_03883_ ), .C1(_03216_ ), .C2(_00434_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
AOI21_X1 _16164_ ( .A(_03078_ ), .B1(_03346_ ), .B2(_03353_ ), .ZN(_00445_ ) );
OAI211_X1 _16165_ ( .A(_03216_ ), .B(_00445_ ), .C1(_03232_ ), .C2(_03273_ ), .ZN(_00446_ ) );
OR2_X1 _16166_ ( .A1(_00446_ ), .A2(_00434_ ), .ZN(_00447_ ) );
OR3_X1 _16167_ ( .A1(_03078_ ), .A2(_00437_ ), .A3(loaduse_clear ), .ZN(_00448_ ) );
AND3_X1 _16168_ ( .A1(_03341_ ), .A2(_03077_ ), .A3(_03344_ ), .ZN(_00449_ ) );
NAND4_X1 _16169_ ( .A1(_03334_ ), .A2(IDU_ready_IFU ), .A3(_03216_ ), .A4(_00449_ ), .ZN(_00450_ ) );
NAND3_X1 _16170_ ( .A1(_00447_ ), .A2(_00448_ ), .A3(_00450_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16171_ ( .A1(_03213_ ), .A2(IDU_ready_IFU ), .ZN(_00451_ ) );
NOR2_X1 _16172_ ( .A1(_03213_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00452_ ) );
NOR2_X1 _16173_ ( .A1(\myifu.state [0] ), .A2(\myifu.state [1] ), .ZN(_00453_ ) );
NOR4_X1 _16174_ ( .A1(_00451_ ), .A2(_00452_ ), .A3(reset ), .A4(_00453_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
CLKBUF_X2 _16175_ ( .A(_06082_ ), .Z(_00454_ ) );
OR3_X1 _16176_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00455_ ) );
OAI21_X1 _16177_ ( .A(_00455_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06084_ ), .ZN(_00456_ ) );
MUX2_X1 _16178_ ( .A(\io_master_rdata [31] ), .B(_00456_ ), .S(_02072_ ), .Z(_00457_ ) );
AND2_X1 _16179_ ( .A1(_00457_ ), .A2(\io_master_arburst [0] ), .ZN(\myifu.data_in [31] ) );
BUF_X4 _16180_ ( .A(_06050_ ), .Z(_00458_ ) );
CLKBUF_X2 _16181_ ( .A(_06082_ ), .Z(_00459_ ) );
OR3_X1 _16182_ ( .A1(_02024_ ), .A2(_01530_ ), .A3(_00459_ ), .ZN(_00460_ ) );
OAI211_X1 _16183_ ( .A(_02072_ ), .B(_00460_ ), .C1(_01649_ ), .C2(_06084_ ), .ZN(_00461_ ) );
OAI21_X1 _16184_ ( .A(\io_master_rdata [30] ), .B1(_01986_ ), .B2(_02022_ ), .ZN(_00462_ ) );
AOI21_X1 _16185_ ( .A(_00458_ ), .B1(_00461_ ), .B2(_00462_ ), .ZN(\myifu.data_in [30] ) );
MUX2_X1 _16186_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\io_master_araddr [2] ), .Z(_00463_ ) );
OR3_X1 _16187_ ( .A1(_01986_ ), .A2(_02022_ ), .A3(_00463_ ), .ZN(_00464_ ) );
OAI21_X1 _16188_ ( .A(\io_master_rdata [21] ), .B1(_01986_ ), .B2(_02022_ ), .ZN(_00465_ ) );
AOI21_X1 _16189_ ( .A(_06049_ ), .B1(_00464_ ), .B2(_00465_ ), .ZN(\myifu.data_in [21] ) );
AND2_X4 _16190_ ( .A1(_03824_ ), .A2(_03827_ ), .ZN(_00466_ ) );
BUF_X16 _16191_ ( .A(_00466_ ), .Z(_00467_ ) );
OR3_X1 _16192_ ( .A1(_01953_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06082_ ), .ZN(_00468_ ) );
OAI211_X1 _16193_ ( .A(_00467_ ), .B(_00468_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06083_ ), .ZN(_00469_ ) );
BUF_X8 _16194_ ( .A(_00466_ ), .Z(_00470_ ) );
OAI21_X2 _16195_ ( .A(_00469_ ), .B1(\io_master_rdata [20] ), .B2(_00470_ ), .ZN(_00471_ ) );
BUF_X4 _16196_ ( .A(_06050_ ), .Z(_00472_ ) );
NOR2_X1 _16197_ ( .A1(_00471_ ), .A2(_00472_ ), .ZN(\myifu.data_in [20] ) );
OR3_X1 _16198_ ( .A1(_01953_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00473_ ) );
OAI211_X1 _16199_ ( .A(_00467_ ), .B(_00473_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06083_ ), .ZN(_00474_ ) );
OAI21_X2 _16200_ ( .A(_00474_ ), .B1(\io_master_rdata [19] ), .B2(_00470_ ), .ZN(_00475_ ) );
NOR2_X1 _16201_ ( .A1(_00475_ ), .A2(_00472_ ), .ZN(\myifu.data_in [19] ) );
OR3_X1 _16202_ ( .A1(_01953_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06082_ ), .ZN(_00476_ ) );
OAI211_X1 _16203_ ( .A(_00467_ ), .B(_00476_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06083_ ), .ZN(_00477_ ) );
OAI21_X2 _16204_ ( .A(_00477_ ), .B1(\io_master_rdata [18] ), .B2(_00470_ ), .ZN(_00478_ ) );
NOR2_X1 _16205_ ( .A1(_00478_ ), .A2(_00472_ ), .ZN(\myifu.data_in [18] ) );
OR3_X1 _16206_ ( .A1(_01953_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00479_ ) );
OAI211_X1 _16207_ ( .A(_00467_ ), .B(_00479_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06083_ ), .ZN(_00480_ ) );
OAI21_X2 _16208_ ( .A(_00480_ ), .B1(\io_master_rdata [17] ), .B2(_00470_ ), .ZN(_00481_ ) );
NOR2_X1 _16209_ ( .A1(_00481_ ), .A2(_00472_ ), .ZN(\myifu.data_in [17] ) );
BUF_X16 _16210_ ( .A(_00467_ ), .Z(_00482_ ) );
BUF_X8 _16211_ ( .A(_00482_ ), .Z(_00483_ ) );
OR2_X1 _16212_ ( .A1(_00483_ ), .A2(\io_master_rdata [16] ), .ZN(_00484_ ) );
BUF_X2 _16213_ ( .A(_00483_ ), .Z(_00485_ ) );
CLKBUF_X2 _16214_ ( .A(_00459_ ), .Z(_00486_ ) );
OR3_X1 _16215_ ( .A1(_02026_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00487_ ) );
OAI211_X1 _16216_ ( .A(_00485_ ), .B(_00487_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00488_ ) );
AND3_X1 _16217_ ( .A1(_00484_ ), .A2(_00488_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16218_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00489_ ) );
OAI211_X1 _16219_ ( .A(_00482_ ), .B(_00489_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06084_ ), .ZN(_00490_ ) );
OAI21_X1 _16220_ ( .A(_00490_ ), .B1(_00482_ ), .B2(\io_master_rdata [15] ), .ZN(_00491_ ) );
NOR2_X1 _16221_ ( .A1(_00491_ ), .A2(_00472_ ), .ZN(\myifu.data_in [15] ) );
BUF_X8 _16222_ ( .A(_00482_ ), .Z(_00492_ ) );
OR2_X1 _16223_ ( .A1(_00492_ ), .A2(\io_master_rdata [14] ), .ZN(_00493_ ) );
OR3_X1 _16224_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00494_ ) );
OAI211_X1 _16225_ ( .A(_00483_ ), .B(_00494_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00495_ ) );
AND3_X1 _16226_ ( .A1(_00493_ ), .A2(_00495_ ), .A3(_02027_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16227_ ( .A1(_00485_ ), .A2(\io_master_rdata [13] ), .ZN(_00496_ ) );
OR3_X1 _16228_ ( .A1(_02026_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00497_ ) );
OAI211_X1 _16229_ ( .A(_00485_ ), .B(_00497_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00498_ ) );
AND3_X1 _16230_ ( .A1(_00496_ ), .A2(_00498_ ), .A3(_02027_ ), .ZN(\myifu.data_in [13] ) );
OR3_X1 _16231_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00499_ ) );
OAI211_X1 _16232_ ( .A(_00483_ ), .B(_00499_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00500_ ) );
OAI21_X1 _16233_ ( .A(_00500_ ), .B1(_00483_ ), .B2(\io_master_rdata [12] ), .ZN(_00501_ ) );
NOR2_X1 _16234_ ( .A1(_00501_ ), .A2(_00472_ ), .ZN(\myifu.data_in [12] ) );
OR2_X1 _16235_ ( .A1(_00483_ ), .A2(\io_master_rdata [29] ), .ZN(_00502_ ) );
OR3_X1 _16236_ ( .A1(_02026_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00503_ ) );
OAI211_X1 _16237_ ( .A(_00485_ ), .B(_00503_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00504_ ) );
AND3_X1 _16238_ ( .A1(_00502_ ), .A2(_00504_ ), .A3(_02027_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16239_ ( .A1(_00492_ ), .A2(\io_master_rdata [11] ), .ZN(_00505_ ) );
OR3_X1 _16240_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00506_ ) );
OAI211_X1 _16241_ ( .A(_00483_ ), .B(_00506_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00507_ ) );
AND3_X1 _16242_ ( .A1(_00505_ ), .A2(_00507_ ), .A3(_02027_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16243_ ( .A1(_00492_ ), .A2(\io_master_rdata [10] ), .ZN(_00508_ ) );
OR3_X1 _16244_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00509_ ) );
OAI211_X1 _16245_ ( .A(_00483_ ), .B(_00509_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00510_ ) );
AND3_X1 _16246_ ( .A1(_00508_ ), .A2(_00510_ ), .A3(_02027_ ), .ZN(\myifu.data_in [10] ) );
OR3_X1 _16247_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00511_ ) );
OAI211_X1 _16248_ ( .A(_00483_ ), .B(_00511_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00512_ ) );
OAI21_X1 _16249_ ( .A(_00512_ ), .B1(_00483_ ), .B2(\io_master_rdata [9] ), .ZN(_00513_ ) );
NOR2_X1 _16250_ ( .A1(_00513_ ), .A2(_00472_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16251_ ( .A1(_00485_ ), .A2(\io_master_rdata [8] ), .ZN(_00514_ ) );
OR3_X1 _16252_ ( .A1(_02026_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00515_ ) );
OAI211_X1 _16253_ ( .A(_00485_ ), .B(_00515_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00516_ ) );
AND3_X1 _16254_ ( .A1(_00514_ ), .A2(_00516_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [8] ) );
OR2_X1 _16255_ ( .A1(_00492_ ), .A2(\io_master_rdata [7] ), .ZN(_00517_ ) );
OR3_X1 _16256_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00518_ ) );
OAI211_X1 _16257_ ( .A(_00492_ ), .B(_00518_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00519_ ) );
AND3_X1 _16258_ ( .A1(_00517_ ), .A2(_00519_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16259_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00520_ ) );
OAI211_X4 _16260_ ( .A(_00470_ ), .B(_00520_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06084_ ), .ZN(_00521_ ) );
OAI21_X4 _16261_ ( .A(_00521_ ), .B1(\io_master_rdata [6] ), .B2(_00482_ ), .ZN(_00522_ ) );
NOR2_X1 _16262_ ( .A1(_00522_ ), .A2(_00472_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16263_ ( .A1(_02026_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00523_ ) );
OAI211_X1 _16264_ ( .A(_00485_ ), .B(_00523_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00524_ ) );
OAI21_X1 _16265_ ( .A(_00524_ ), .B1(\io_master_rdata [5] ), .B2(_00485_ ), .ZN(_00525_ ) );
NOR2_X1 _16266_ ( .A1(_00525_ ), .A2(_00472_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16267_ ( .A1(_01953_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00526_ ) );
OAI211_X2 _16268_ ( .A(_00467_ ), .B(_00526_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06084_ ), .ZN(_00527_ ) );
OAI21_X2 _16269_ ( .A(_00527_ ), .B1(\io_master_rdata [4] ), .B2(_00470_ ), .ZN(_00528_ ) );
NOR2_X1 _16270_ ( .A1(_00528_ ), .A2(_00472_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16271_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00529_ ) );
OAI211_X2 _16272_ ( .A(_00467_ ), .B(_00529_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06084_ ), .ZN(_00530_ ) );
OAI21_X2 _16273_ ( .A(_00530_ ), .B1(\io_master_rdata [3] ), .B2(_00470_ ), .ZN(_00531_ ) );
NOR2_X1 _16274_ ( .A1(_00531_ ), .A2(_00458_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16275_ ( .A1(_01953_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00532_ ) );
OAI211_X1 _16276_ ( .A(_00467_ ), .B(_00532_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06083_ ), .ZN(_00533_ ) );
OAI21_X2 _16277_ ( .A(_00533_ ), .B1(\io_master_rdata [2] ), .B2(_00470_ ), .ZN(_00534_ ) );
NOR2_X1 _16278_ ( .A1(_00534_ ), .A2(_00458_ ), .ZN(\myifu.data_in [2] ) );
OR3_X1 _16279_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00535_ ) );
OAI211_X1 _16280_ ( .A(_00482_ ), .B(_00535_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00536_ ) );
OAI21_X2 _16281_ ( .A(_00536_ ), .B1(_00492_ ), .B2(\io_master_rdata [28] ), .ZN(_00537_ ) );
NOR2_X1 _16282_ ( .A1(_00537_ ), .A2(_00458_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16283_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00538_ ) );
OAI211_X2 _16284_ ( .A(_00467_ ), .B(_00538_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06084_ ), .ZN(_00539_ ) );
OAI21_X2 _16285_ ( .A(_00539_ ), .B1(\io_master_rdata [1] ), .B2(_00470_ ), .ZN(_00540_ ) );
NOR2_X1 _16286_ ( .A1(_00540_ ), .A2(_00458_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16287_ ( .A1(_02026_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00486_ ), .ZN(_00541_ ) );
OAI211_X1 _16288_ ( .A(_00485_ ), .B(_00541_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00542_ ) );
OAI21_X1 _16289_ ( .A(_00542_ ), .B1(\io_master_rdata [0] ), .B2(_00485_ ), .ZN(_00543_ ) );
NOR2_X1 _16290_ ( .A1(_00543_ ), .A2(_00458_ ), .ZN(\myifu.data_in [0] ) );
OR3_X1 _16291_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00544_ ) );
OAI211_X1 _16292_ ( .A(_00482_ ), .B(_00544_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06084_ ), .ZN(_00545_ ) );
OAI21_X2 _16293_ ( .A(_00545_ ), .B1(_00492_ ), .B2(\io_master_rdata [27] ), .ZN(_00546_ ) );
NOR2_X1 _16294_ ( .A1(_00546_ ), .A2(_00458_ ), .ZN(\myifu.data_in [27] ) );
OR3_X1 _16295_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00547_ ) );
OAI211_X1 _16296_ ( .A(_00482_ ), .B(_00547_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00548_ ) );
OAI21_X2 _16297_ ( .A(_00548_ ), .B1(_00492_ ), .B2(\io_master_rdata [26] ), .ZN(_00549_ ) );
NOR2_X1 _16298_ ( .A1(_00549_ ), .A2(_00458_ ), .ZN(\myifu.data_in [26] ) );
OR3_X1 _16299_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00550_ ) );
OAI211_X1 _16300_ ( .A(_00482_ ), .B(_00550_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00551_ ) );
OAI21_X2 _16301_ ( .A(_00551_ ), .B1(\io_master_rdata [25] ), .B2(_00492_ ), .ZN(_00552_ ) );
NOR2_X1 _16302_ ( .A1(_00552_ ), .A2(_00458_ ), .ZN(\myifu.data_in [25] ) );
OR3_X1 _16303_ ( .A1(_02026_ ), .A2(_01735_ ), .A3(_00486_ ), .ZN(_00553_ ) );
OAI211_X1 _16304_ ( .A(_02072_ ), .B(_00553_ ), .C1(_01669_ ), .C2(\io_master_araddr [2] ), .ZN(_00554_ ) );
OAI21_X1 _16305_ ( .A(\io_master_rdata [24] ), .B1(_01986_ ), .B2(_02022_ ), .ZN(_00555_ ) );
AOI21_X1 _16306_ ( .A(_06051_ ), .B1(_00554_ ), .B2(_00555_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16307_ ( .A1(_02025_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00459_ ), .ZN(_00556_ ) );
OAI211_X1 _16308_ ( .A(_00482_ ), .B(_00556_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06085_ ), .ZN(_00557_ ) );
OAI21_X1 _16309_ ( .A(_00557_ ), .B1(_00492_ ), .B2(\io_master_rdata [23] ), .ZN(_00558_ ) );
NOR2_X1 _16310_ ( .A1(_00558_ ), .A2(_00458_ ), .ZN(\myifu.data_in [23] ) );
OR2_X2 _16311_ ( .A1(_00467_ ), .A2(\io_master_rdata [22] ), .ZN(_00559_ ) );
OR3_X1 _16312_ ( .A1(_02024_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00454_ ), .ZN(_00560_ ) );
OAI211_X2 _16313_ ( .A(_00470_ ), .B(_00560_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06084_ ), .ZN(_00561_ ) );
AND3_X1 _16314_ ( .A1(_00559_ ), .A2(_00561_ ), .A3(_02027_ ), .ZN(\myifu.data_in [22] ) );
OR2_X1 _16315_ ( .A1(_00242_ ), .A2(_02063_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
OAI21_X1 _16316_ ( .A(_02062_ ), .B1(_06005_ ), .B2(_06007_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
OAI21_X1 _16317_ ( .A(_02062_ ), .B1(_06008_ ), .B2(_06007_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16318_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .ZN(_00562_ ) );
OAI21_X1 _16319_ ( .A(_02062_ ), .B1(_00562_ ), .B2(_06007_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
AOI221_X4 _16320_ ( .A(_03488_ ), .B1(\IF_ID_inst [16] ), .B2(_03083_ ), .C1(_03232_ ), .C2(\IF_ID_inst [8] ), .ZN(_00563_ ) );
AND4_X1 _16321_ ( .A1(_03074_ ), .A2(_03306_ ), .A3(_03380_ ), .A4(_03381_ ), .ZN(_00564_ ) );
AND4_X1 _16322_ ( .A1(_03261_ ), .A2(_03376_ ), .A3(_03312_ ), .A4(_00564_ ), .ZN(_00565_ ) );
AND2_X1 _16323_ ( .A1(_03231_ ), .A2(_03396_ ), .ZN(_00566_ ) );
AND2_X1 _16324_ ( .A1(_00565_ ), .A2(_00566_ ), .ZN(_00567_ ) );
INV_X1 _16325_ ( .A(_00567_ ), .ZN(_00568_ ) );
OAI21_X1 _16326_ ( .A(_00563_ ), .B1(_00568_ ), .B2(_03081_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
AND3_X1 _16327_ ( .A1(_03159_ ), .A2(\IF_ID_inst [31] ), .A3(_03123_ ), .ZN(_00569_ ) );
INV_X1 _16328_ ( .A(_00569_ ), .ZN(_00570_ ) );
OAI221_X1 _16329_ ( .A(_00570_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03291_ ), .C1(_00566_ ), .C2(_03076_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
NOR2_X1 _16330_ ( .A1(_03291_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00571_ ) );
INV_X1 _16331_ ( .A(_00571_ ), .ZN(_00572_ ) );
OR2_X1 _16332_ ( .A1(_03231_ ), .A2(_03076_ ), .ZN(_00573_ ) );
AND2_X1 _16333_ ( .A1(_00572_ ), .A2(_00573_ ), .ZN(_00574_ ) );
BUF_X4 _16334_ ( .A(_00574_ ), .Z(_00575_ ) );
BUF_X4 _16335_ ( .A(_00570_ ), .Z(_00576_ ) );
BUF_X4 _16336_ ( .A(_03396_ ), .Z(_00577_ ) );
OAI211_X1 _16337_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03080_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16338_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03081_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16339_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03084_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
OAI21_X1 _16340_ ( .A(\IF_ID_inst [19] ), .B1(_03161_ ), .B2(_03166_ ), .ZN(_00578_ ) );
BUF_X2 _16341_ ( .A(_03231_ ), .Z(_00579_ ) );
BUF_X2 _16342_ ( .A(_03291_ ), .Z(_00580_ ) );
OAI221_X1 _16343_ ( .A(_00578_ ), .B1(_00579_ ), .B2(_03076_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI21_X1 _16344_ ( .A(\IF_ID_inst [18] ), .B1(_03161_ ), .B2(_03166_ ), .ZN(_00581_ ) );
OAI221_X1 _16345_ ( .A(_00581_ ), .B1(_00579_ ), .B2(_03076_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI21_X1 _16346_ ( .A(\IF_ID_inst [17] ), .B1(_03161_ ), .B2(_03166_ ), .ZN(_00582_ ) );
OAI221_X1 _16347_ ( .A(_00582_ ), .B1(_00579_ ), .B2(_03076_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI21_X1 _16348_ ( .A(\IF_ID_inst [16] ), .B1(_03161_ ), .B2(_03166_ ), .ZN(_00583_ ) );
OAI221_X1 _16349_ ( .A(_00583_ ), .B1(_00579_ ), .B2(_03076_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
INV_X1 _16350_ ( .A(\IF_ID_inst [15] ), .ZN(_00584_ ) );
NOR2_X1 _16351_ ( .A1(_03161_ ), .A2(_03166_ ), .ZN(_00585_ ) );
OAI221_X1 _16352_ ( .A(_00573_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03291_ ), .C1(_00584_ ), .C2(_00585_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16353_ ( .A(_00573_ ), .B1(_03131_ ), .B2(_00585_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00580_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16354_ ( .A(_00573_ ), .B1(_03139_ ), .B2(_00585_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_03291_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16355_ ( .A(_00573_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03291_ ), .C1(_03142_ ), .C2(_00585_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16356_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03085_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
OR2_X1 _16357_ ( .A1(_03223_ ), .A2(_03100_ ), .ZN(_00586_ ) );
OR2_X1 _16358_ ( .A1(_03366_ ), .A2(_03076_ ), .ZN(_00587_ ) );
NAND4_X1 _16359_ ( .A1(_00572_ ), .A2(_03438_ ), .A3(_00586_ ), .A4(_00587_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16360_ ( .A(_03452_ ), .ZN(_00588_ ) );
OAI221_X1 _16361_ ( .A(_00588_ ), .B1(_00579_ ), .B2(_03080_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
OAI221_X1 _16362_ ( .A(_03448_ ), .B1(_00579_ ), .B2(_03085_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16363_ ( .A(_03522_ ), .ZN(_00589_ ) );
OAI221_X1 _16364_ ( .A(_00589_ ), .B1(_00579_ ), .B2(_03086_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
INV_X1 _16365_ ( .A(_03515_ ), .ZN(_00590_ ) );
OAI221_X1 _16366_ ( .A(_00590_ ), .B1(_00579_ ), .B2(_03087_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16367_ ( .A(_03475_ ), .ZN(_00591_ ) );
OAI221_X1 _16368_ ( .A(_00591_ ), .B1(_00579_ ), .B2(_03088_ ), .C1(_00580_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
OR2_X1 _16369_ ( .A1(_00579_ ), .A2(_03089_ ), .ZN(_00592_ ) );
OAI221_X1 _16370_ ( .A(_00592_ ), .B1(_03089_ ), .B2(_03311_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .C2(_03291_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16371_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03086_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16372_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03087_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16373_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03088_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16374_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03089_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16375_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03090_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16376_ ( .A(_00575_ ), .B(_00576_ ), .C1(_03092_ ), .C2(_00577_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16377_ ( .A(_00574_ ), .B(_00570_ ), .C1(_03093_ ), .C2(_03396_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
AOI221_X4 _16378_ ( .A(_03506_ ), .B1(\IF_ID_inst [19] ), .B2(_03083_ ), .C1(_03232_ ), .C2(\IF_ID_inst [11] ), .ZN(_00593_ ) );
OAI21_X1 _16379_ ( .A(_00593_ ), .B1(_00568_ ), .B2(_03090_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
AOI221_X4 _16380_ ( .A(_03497_ ), .B1(\IF_ID_inst [18] ), .B2(_03083_ ), .C1(_03232_ ), .C2(\IF_ID_inst [10] ), .ZN(_00594_ ) );
OAI21_X1 _16381_ ( .A(_00594_ ), .B1(_00568_ ), .B2(_03092_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
AOI22_X1 _16382_ ( .A1(_03232_ ), .A2(\IF_ID_inst [9] ), .B1(\IF_ID_inst [17] ), .B2(_03083_ ), .ZN(_00595_ ) );
AOI21_X1 _16383_ ( .A(_03161_ ), .B1(_00565_ ), .B2(_00566_ ), .ZN(_00596_ ) );
OAI21_X1 _16384_ ( .A(_00595_ ), .B1(_00596_ ), .B2(_03093_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16385_ ( .A1(_03366_ ), .A2(_03100_ ), .ZN(_00597_ ) );
OAI221_X1 _16386_ ( .A(_00597_ ), .B1(_00584_ ), .B2(_03075_ ), .C1(_00568_ ), .C2(_03084_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AND2_X2 _16387_ ( .A1(_03819_ ), .A2(_03830_ ), .ZN(_00598_ ) );
BUF_X4 _16388_ ( .A(_00598_ ), .Z(_00599_ ) );
AOI21_X1 _16389_ ( .A(\IF_ID_pc [1] ), .B1(_03832_ ), .B2(\IF_ID_pc [2] ), .ZN(_00600_ ) );
INV_X1 _16390_ ( .A(_00600_ ), .ZN(_00601_ ) );
OAI21_X1 _16391_ ( .A(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .B1(_03832_ ), .B2(\IF_ID_pc [2] ), .ZN(_00602_ ) );
NOR2_X1 _16392_ ( .A1(_00601_ ), .A2(_00602_ ), .ZN(_00603_ ) );
BUF_X4 _16393_ ( .A(_00603_ ), .Z(_00604_ ) );
NAND2_X1 _16394_ ( .A1(_00514_ ), .A2(_00516_ ), .ZN(_00605_ ) );
BUF_X4 _16395_ ( .A(_06049_ ), .Z(_00606_ ) );
OAI211_X1 _16396_ ( .A(_00599_ ), .B(_00604_ ), .C1(_00605_ ), .C2(_00606_ ), .ZN(_00607_ ) );
AND2_X1 _16397_ ( .A1(_00598_ ), .A2(_00603_ ), .ZN(_00608_ ) );
BUF_X4 _16398_ ( .A(_00608_ ), .Z(_00609_ ) );
BUF_X4 _16399_ ( .A(_00609_ ), .Z(_00610_ ) );
OAI211_X1 _16400_ ( .A(_00607_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_03489_ ), .ZN(_00611_ ) );
AND3_X1 _16401_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00612_ ) );
AND3_X1 _16402_ ( .A1(_03747_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00613_ ) );
AOI211_X1 _16403_ ( .A(_00612_ ), .B(_00613_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_06004_ ), .ZN(_00614_ ) );
NAND2_X1 _16404_ ( .A1(_06006_ ), .A2(\IF_ID_pc [2] ), .ZN(_00615_ ) );
BUF_X2 _16405_ ( .A(_00615_ ), .Z(_00616_ ) );
NAND2_X2 _16406_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00617_ ) );
BUF_X4 _16407_ ( .A(_00617_ ), .Z(_00618_ ) );
BUF_X4 _16408_ ( .A(_00618_ ), .Z(_00619_ ) );
NAND3_X1 _16409_ ( .A1(_03756_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00620_ ) );
NAND4_X1 _16410_ ( .A1(_00614_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00620_ ), .ZN(_00621_ ) );
NOR2_X1 _16411_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00622_ ) );
BUF_X4 _16412_ ( .A(_00622_ ), .Z(_00623_ ) );
BUF_X4 _16413_ ( .A(_00623_ ), .Z(_00624_ ) );
BUF_X4 _16414_ ( .A(_03746_ ), .Z(_00625_ ) );
BUF_X4 _16415_ ( .A(_00625_ ), .Z(_00626_ ) );
NAND3_X1 _16416_ ( .A1(_00626_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00627_ ) );
NAND3_X1 _16417_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00628_ ) );
AND2_X1 _16418_ ( .A1(_00627_ ), .A2(_00628_ ), .ZN(_00629_ ) );
NAND2_X1 _16419_ ( .A1(_00615_ ), .A2(_00617_ ), .ZN(_00630_ ) );
BUF_X2 _16420_ ( .A(_00630_ ), .Z(_00631_ ) );
BUF_X4 _16421_ ( .A(_03755_ ), .Z(_00632_ ) );
BUF_X4 _16422_ ( .A(_00632_ ), .Z(_00633_ ) );
NAND3_X1 _16423_ ( .A1(_00633_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00634_ ) );
BUF_X4 _16424_ ( .A(_03755_ ), .Z(_00635_ ) );
BUF_X4 _16425_ ( .A(_00635_ ), .Z(_00636_ ) );
NAND3_X1 _16426_ ( .A1(_03748_ ), .A2(_00636_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00637_ ) );
NAND4_X1 _16427_ ( .A1(_00629_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00637_ ), .ZN(_00638_ ) );
NAND3_X1 _16428_ ( .A1(_00621_ ), .A2(_00624_ ), .A3(_00638_ ), .ZN(_00639_ ) );
NAND2_X1 _16429_ ( .A1(_00611_ ), .A2(_00639_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16430_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00640_ ) );
CLKBUF_X2 _16431_ ( .A(_03746_ ), .Z(_00641_ ) );
AND3_X1 _16432_ ( .A1(_00641_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00642_ ) );
BUF_X4 _16433_ ( .A(_06003_ ), .Z(_00643_ ) );
AOI211_X1 _16434_ ( .A(_00640_ ), .B(_00642_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00643_ ), .ZN(_00644_ ) );
BUF_X4 _16435_ ( .A(_00615_ ), .Z(_00645_ ) );
BUF_X4 _16436_ ( .A(_00635_ ), .Z(_00646_ ) );
NAND3_X1 _16437_ ( .A1(_00646_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00647_ ) );
NAND4_X1 _16438_ ( .A1(_00644_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_00647_ ), .ZN(_00648_ ) );
BUF_X4 _16439_ ( .A(_00625_ ), .Z(_00649_ ) );
NAND3_X1 _16440_ ( .A1(_00649_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00650_ ) );
NAND3_X1 _16441_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00651_ ) );
AND2_X1 _16442_ ( .A1(_00650_ ), .A2(_00651_ ), .ZN(_00652_ ) );
BUF_X4 _16443_ ( .A(_00630_ ), .Z(_00653_ ) );
BUF_X4 _16444_ ( .A(_00653_ ), .Z(_00654_ ) );
BUF_X4 _16445_ ( .A(_00635_ ), .Z(_00655_ ) );
NAND3_X1 _16446_ ( .A1(_00655_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00656_ ) );
BUF_X4 _16447_ ( .A(_03747_ ), .Z(_00657_ ) );
NAND3_X1 _16448_ ( .A1(_00657_ ), .A2(_00632_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00658_ ) );
NAND4_X1 _16449_ ( .A1(_00652_ ), .A2(_00654_ ), .A3(_00656_ ), .A4(_00658_ ), .ZN(_00659_ ) );
NAND3_X1 _16450_ ( .A1(_00648_ ), .A2(_00623_ ), .A3(_00659_ ), .ZN(_00660_ ) );
OAI21_X1 _16451_ ( .A(\myifu.state [2] ), .B1(_00609_ ), .B2(_03251_ ), .ZN(_00661_ ) );
OAI21_X1 _16452_ ( .A(_02026_ ), .B1(_02072_ ), .B2(_03816_ ), .ZN(_00662_ ) );
AND3_X1 _16453_ ( .A1(_02068_ ), .A2(_01975_ ), .A3(_02071_ ), .ZN(_00663_ ) );
AND2_X1 _16454_ ( .A1(_03817_ ), .A2(\io_master_rid [0] ), .ZN(_00664_ ) );
AOI21_X1 _16455_ ( .A(_00664_ ), .B1(_02068_ ), .B2(_02071_ ), .ZN(_00665_ ) );
NOR3_X1 _16456_ ( .A1(_00662_ ), .A2(_00663_ ), .A3(_00665_ ), .ZN(_00666_ ) );
OAI21_X1 _16457_ ( .A(_02026_ ), .B1(_02072_ ), .B2(_03815_ ), .ZN(_00667_ ) );
NOR3_X1 _16458_ ( .A1(_00667_ ), .A2(_03829_ ), .A3(_03828_ ), .ZN(_00668_ ) );
NAND2_X1 _16459_ ( .A1(_00666_ ), .A2(_00668_ ), .ZN(_00669_ ) );
NOR4_X1 _16460_ ( .A1(\myifu.data_in [31] ), .A2(_00669_ ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_00670_ ) );
OAI21_X1 _16461_ ( .A(_00660_ ), .B1(_00661_ ), .B2(_00670_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
AND2_X1 _16462_ ( .A1(_00461_ ), .A2(_00462_ ), .ZN(_00671_ ) );
OAI211_X1 _16463_ ( .A(_00599_ ), .B(_00604_ ), .C1(_00671_ ), .C2(_06049_ ), .ZN(_00672_ ) );
OAI211_X1 _16464_ ( .A(_00672_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_03453_ ), .ZN(_00673_ ) );
AND3_X1 _16465_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00674_ ) );
AND3_X1 _16466_ ( .A1(_03747_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00675_ ) );
AOI211_X1 _16467_ ( .A(_00674_ ), .B(_00675_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_06004_ ), .ZN(_00676_ ) );
NAND3_X1 _16468_ ( .A1(_03756_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00677_ ) );
NAND4_X1 _16469_ ( .A1(_00676_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00677_ ), .ZN(_00678_ ) );
NAND3_X1 _16470_ ( .A1(_00626_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00679_ ) );
NAND3_X1 _16471_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00680_ ) );
AND2_X1 _16472_ ( .A1(_00679_ ), .A2(_00680_ ), .ZN(_00681_ ) );
NAND3_X1 _16473_ ( .A1(_00633_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00682_ ) );
NAND3_X1 _16474_ ( .A1(_03748_ ), .A2(_00636_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00683_ ) );
NAND4_X1 _16475_ ( .A1(_00681_ ), .A2(_00631_ ), .A3(_00682_ ), .A4(_00683_ ), .ZN(_00684_ ) );
NAND3_X1 _16476_ ( .A1(_00678_ ), .A2(_00624_ ), .A3(_00684_ ), .ZN(_00685_ ) );
NAND2_X1 _16477_ ( .A1(_00673_ ), .A2(_00685_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
AND3_X1 _16478_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00686_ ) );
AND3_X1 _16479_ ( .A1(_00625_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00687_ ) );
AOI211_X1 _16480_ ( .A(_00686_ ), .B(_00687_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_00643_ ), .ZN(_00688_ ) );
NAND3_X1 _16481_ ( .A1(_00646_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00689_ ) );
NAND4_X1 _16482_ ( .A1(_00688_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_00689_ ), .ZN(_00690_ ) );
NAND3_X1 _16483_ ( .A1(_00649_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00691_ ) );
NAND3_X1 _16484_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00692_ ) );
AND2_X1 _16485_ ( .A1(_00691_ ), .A2(_00692_ ), .ZN(_00693_ ) );
NAND3_X1 _16486_ ( .A1(_00655_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00694_ ) );
NAND3_X1 _16487_ ( .A1(_00657_ ), .A2(_00632_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00695_ ) );
NAND4_X1 _16488_ ( .A1(_00693_ ), .A2(_00653_ ), .A3(_00694_ ), .A4(_00695_ ), .ZN(_00696_ ) );
NAND3_X1 _16489_ ( .A1(_00690_ ), .A2(_00623_ ), .A3(_00696_ ), .ZN(_00697_ ) );
INV_X1 _16490_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00698_ ) );
OAI21_X1 _16491_ ( .A(\myifu.state [2] ), .B1(_00609_ ), .B2(_00698_ ), .ZN(_00699_ ) );
NOR4_X1 _16492_ ( .A1(_00669_ ), .A2(\myifu.data_in [21] ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_00700_ ) );
OAI21_X1 _16493_ ( .A(_00697_ ), .B1(_00699_ ), .B2(_00700_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
INV_X1 _16494_ ( .A(\myifu.state [2] ), .ZN(_00701_ ) );
INV_X1 _16495_ ( .A(_00608_ ), .ZN(_00702_ ) );
BUF_X4 _16496_ ( .A(_00702_ ), .Z(_00703_ ) );
AOI21_X1 _16497_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00704_ ) );
OAI211_X1 _16498_ ( .A(_00599_ ), .B(_00604_ ), .C1(_00471_ ), .C2(_06050_ ), .ZN(_00705_ ) );
NAND2_X1 _16499_ ( .A1(_00704_ ), .A2(_00705_ ), .ZN(_00706_ ) );
AND3_X1 _16500_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00707_ ) );
AND3_X1 _16501_ ( .A1(_03747_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00708_ ) );
AOI211_X1 _16502_ ( .A(_00707_ ), .B(_00708_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_06004_ ), .ZN(_00709_ ) );
NAND3_X1 _16503_ ( .A1(_03756_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00710_ ) );
NAND4_X1 _16504_ ( .A1(_00709_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00710_ ), .ZN(_00711_ ) );
NAND3_X1 _16505_ ( .A1(_00626_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00712_ ) );
NAND3_X1 _16506_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00713_ ) );
AND2_X1 _16507_ ( .A1(_00712_ ), .A2(_00713_ ), .ZN(_00714_ ) );
NAND3_X1 _16508_ ( .A1(_00633_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00715_ ) );
NAND3_X1 _16509_ ( .A1(_03748_ ), .A2(_00636_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00716_ ) );
NAND4_X1 _16510_ ( .A1(_00714_ ), .A2(_00631_ ), .A3(_00715_ ), .A4(_00716_ ), .ZN(_00717_ ) );
NAND3_X1 _16511_ ( .A1(_00711_ ), .A2(_00624_ ), .A3(_00717_ ), .ZN(_00718_ ) );
NAND2_X1 _16512_ ( .A1(_00706_ ), .A2(_00718_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
AOI21_X1 _16513_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00719_ ) );
OAI211_X1 _16514_ ( .A(_00599_ ), .B(_00604_ ), .C1(_00475_ ), .C2(_06050_ ), .ZN(_00720_ ) );
NAND2_X1 _16515_ ( .A1(_00719_ ), .A2(_00720_ ), .ZN(_00721_ ) );
AND3_X1 _16516_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00722_ ) );
CLKBUF_X2 _16517_ ( .A(_03746_ ), .Z(_00723_ ) );
AND3_X1 _16518_ ( .A1(_00723_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00724_ ) );
AOI211_X1 _16519_ ( .A(_00722_ ), .B(_00724_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_06004_ ), .ZN(_00725_ ) );
NAND3_X1 _16520_ ( .A1(_03756_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00726_ ) );
NAND4_X1 _16521_ ( .A1(_00725_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00726_ ), .ZN(_00727_ ) );
NAND3_X1 _16522_ ( .A1(_00626_ ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00728_ ) );
NAND3_X1 _16523_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00729_ ) );
AND2_X1 _16524_ ( .A1(_00728_ ), .A2(_00729_ ), .ZN(_00730_ ) );
BUF_X4 _16525_ ( .A(_00653_ ), .Z(_00731_ ) );
NAND3_X1 _16526_ ( .A1(_00633_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00732_ ) );
NAND3_X1 _16527_ ( .A1(_03748_ ), .A2(_00636_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00733_ ) );
NAND4_X1 _16528_ ( .A1(_00730_ ), .A2(_00731_ ), .A3(_00732_ ), .A4(_00733_ ), .ZN(_00734_ ) );
NAND3_X1 _16529_ ( .A1(_00727_ ), .A2(_00624_ ), .A3(_00734_ ), .ZN(_00735_ ) );
NAND2_X1 _16530_ ( .A1(_00721_ ), .A2(_00735_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
BUF_X4 _16531_ ( .A(_00598_ ), .Z(_00736_ ) );
BUF_X4 _16532_ ( .A(_00603_ ), .Z(_00737_ ) );
OAI211_X1 _16533_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00478_ ), .C2(_06049_ ), .ZN(_00738_ ) );
INV_X1 _16534_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00739_ ) );
OAI211_X1 _16535_ ( .A(_00738_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_00739_ ), .ZN(_00740_ ) );
AND3_X1 _16536_ ( .A1(fanout_net_10 ), .A2(fanout_net_6 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00741_ ) );
AND3_X1 _16537_ ( .A1(_00723_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00742_ ) );
AOI211_X1 _16538_ ( .A(_00741_ ), .B(_00742_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_06004_ ), .ZN(_00743_ ) );
NAND3_X1 _16539_ ( .A1(_03756_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00744_ ) );
NAND4_X1 _16540_ ( .A1(_00743_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00744_ ), .ZN(_00745_ ) );
NAND3_X1 _16541_ ( .A1(_00626_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00746_ ) );
NAND3_X1 _16542_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00747_ ) );
AND2_X1 _16543_ ( .A1(_00746_ ), .A2(_00747_ ), .ZN(_00748_ ) );
BUF_X4 _16544_ ( .A(_00635_ ), .Z(_00749_ ) );
NAND3_X1 _16545_ ( .A1(_00749_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00750_ ) );
NAND3_X1 _16546_ ( .A1(_03748_ ), .A2(_00636_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00751_ ) );
NAND4_X1 _16547_ ( .A1(_00748_ ), .A2(_00731_ ), .A3(_00750_ ), .A4(_00751_ ), .ZN(_00752_ ) );
NAND3_X1 _16548_ ( .A1(_00745_ ), .A2(_00624_ ), .A3(_00752_ ), .ZN(_00753_ ) );
NAND2_X1 _16549_ ( .A1(_00740_ ), .A2(_00753_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
OAI211_X1 _16550_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00481_ ), .C2(_06049_ ), .ZN(_00754_ ) );
INV_X1 _16551_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00755_ ) );
OAI211_X1 _16552_ ( .A(_00754_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_00755_ ), .ZN(_00756_ ) );
AND3_X1 _16553_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00757_ ) );
AND3_X1 _16554_ ( .A1(_00723_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00758_ ) );
AOI211_X1 _16555_ ( .A(_00757_ ), .B(_00758_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_06004_ ), .ZN(_00759_ ) );
NAND3_X1 _16556_ ( .A1(_03756_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00760_ ) );
NAND4_X1 _16557_ ( .A1(_00759_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00760_ ), .ZN(_00761_ ) );
NAND3_X1 _16558_ ( .A1(_00626_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00762_ ) );
NAND3_X1 _16559_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00763_ ) );
AND2_X1 _16560_ ( .A1(_00762_ ), .A2(_00763_ ), .ZN(_00764_ ) );
NAND3_X1 _16561_ ( .A1(_00749_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00765_ ) );
NAND3_X1 _16562_ ( .A1(_03748_ ), .A2(_00636_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00766_ ) );
NAND4_X1 _16563_ ( .A1(_00764_ ), .A2(_00731_ ), .A3(_00765_ ), .A4(_00766_ ), .ZN(_00767_ ) );
NAND3_X1 _16564_ ( .A1(_00761_ ), .A2(_00624_ ), .A3(_00767_ ), .ZN(_00768_ ) );
NAND2_X1 _16565_ ( .A1(_00756_ ), .A2(_00768_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NAND2_X1 _16566_ ( .A1(_00484_ ), .A2(_00488_ ), .ZN(_00769_ ) );
OAI211_X1 _16567_ ( .A(_00598_ ), .B(_00603_ ), .C1(_00769_ ), .C2(_01954_ ), .ZN(_00770_ ) );
NAND2_X1 _16568_ ( .A1(_00770_ ), .A2(\myifu.state [2] ), .ZN(_00771_ ) );
AOI21_X1 _16569_ ( .A(_00771_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00703_ ), .ZN(_00772_ ) );
AND3_X1 _16570_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00773_ ) );
AND3_X1 _16571_ ( .A1(_03746_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00774_ ) );
AOI211_X1 _16572_ ( .A(_00773_ ), .B(_00774_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_06003_ ), .ZN(_00775_ ) );
NAND3_X1 _16573_ ( .A1(_00635_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00776_ ) );
NAND4_X1 _16574_ ( .A1(_00775_ ), .A2(_00615_ ), .A3(_00617_ ), .A4(_00776_ ), .ZN(_00777_ ) );
NAND3_X1 _16575_ ( .A1(_00625_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00778_ ) );
NAND3_X1 _16576_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00779_ ) );
AND2_X1 _16577_ ( .A1(_00778_ ), .A2(_00779_ ), .ZN(_00780_ ) );
NAND3_X1 _16578_ ( .A1(_00635_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00781_ ) );
NAND3_X1 _16579_ ( .A1(_03747_ ), .A2(_03755_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00782_ ) );
NAND4_X1 _16580_ ( .A1(_00780_ ), .A2(_00653_ ), .A3(_00781_ ), .A4(_00782_ ), .ZN(_00783_ ) );
AND3_X1 _16581_ ( .A1(_00777_ ), .A2(_00622_ ), .A3(_00783_ ), .ZN(_00784_ ) );
OR2_X1 _16582_ ( .A1(_00772_ ), .A2(_00784_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
OAI211_X1 _16583_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00606_ ), .C2(_00491_ ), .ZN(_00785_ ) );
INV_X1 _16584_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00786_ ) );
OAI211_X1 _16585_ ( .A(_00785_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_00786_ ), .ZN(_00787_ ) );
AND3_X1 _16586_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00788_ ) );
AND3_X1 _16587_ ( .A1(_00723_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00789_ ) );
BUF_X4 _16588_ ( .A(_06003_ ), .Z(_00790_ ) );
AOI211_X1 _16589_ ( .A(_00788_ ), .B(_00789_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_00790_ ), .ZN(_00791_ ) );
BUF_X4 _16590_ ( .A(_00632_ ), .Z(_00792_ ) );
NAND3_X1 _16591_ ( .A1(_00792_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00793_ ) );
NAND4_X1 _16592_ ( .A1(_00791_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00793_ ), .ZN(_00794_ ) );
NAND3_X1 _16593_ ( .A1(_00626_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00795_ ) );
NAND3_X1 _16594_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00796_ ) );
AND2_X1 _16595_ ( .A1(_00795_ ), .A2(_00796_ ), .ZN(_00797_ ) );
NAND3_X1 _16596_ ( .A1(_00749_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00798_ ) );
BUF_X4 _16597_ ( .A(_03747_ ), .Z(_00799_ ) );
BUF_X4 _16598_ ( .A(_00635_ ), .Z(_00800_ ) );
NAND3_X1 _16599_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00801_ ) );
NAND4_X1 _16600_ ( .A1(_00797_ ), .A2(_00731_ ), .A3(_00798_ ), .A4(_00801_ ), .ZN(_00802_ ) );
NAND3_X1 _16601_ ( .A1(_00794_ ), .A2(_00624_ ), .A3(_00802_ ), .ZN(_00803_ ) );
NAND2_X1 _16602_ ( .A1(_00787_ ), .A2(_00803_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
AND3_X1 _16603_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00804_ ) );
AND3_X1 _16604_ ( .A1(_00625_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00805_ ) );
AOI211_X1 _16605_ ( .A(_00804_ ), .B(_00805_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_00643_ ), .ZN(_00806_ ) );
NAND3_X1 _16606_ ( .A1(_00636_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00807_ ) );
NAND4_X1 _16607_ ( .A1(_00806_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_00807_ ), .ZN(_00808_ ) );
NAND3_X1 _16608_ ( .A1(_00649_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00809_ ) );
NAND3_X1 _16609_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00810_ ) );
AND2_X1 _16610_ ( .A1(_00809_ ), .A2(_00810_ ), .ZN(_00811_ ) );
NAND3_X1 _16611_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00812_ ) );
NAND3_X1 _16612_ ( .A1(_00657_ ), .A2(_00632_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00813_ ) );
NAND4_X1 _16613_ ( .A1(_00811_ ), .A2(_00653_ ), .A3(_00812_ ), .A4(_00813_ ), .ZN(_00814_ ) );
NAND3_X1 _16614_ ( .A1(_00808_ ), .A2(_00623_ ), .A3(_00814_ ), .ZN(_00815_ ) );
INV_X1 _16615_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00816_ ) );
OAI21_X1 _16616_ ( .A(\myifu.state [2] ), .B1(_00609_ ), .B2(_00816_ ), .ZN(_00817_ ) );
NOR4_X1 _16617_ ( .A1(\myifu.data_in [14] ), .A2(_00669_ ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_00818_ ) );
OAI21_X1 _16618_ ( .A(_00815_ ), .B1(_00817_ ), .B2(_00818_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
AND3_X1 _16619_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00819_ ) );
AND3_X1 _16620_ ( .A1(_00625_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00820_ ) );
AOI211_X1 _16621_ ( .A(_00819_ ), .B(_00820_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_00643_ ), .ZN(_00821_ ) );
NAND3_X1 _16622_ ( .A1(_00636_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00822_ ) );
NAND4_X1 _16623_ ( .A1(_00821_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_00822_ ), .ZN(_00823_ ) );
NAND3_X1 _16624_ ( .A1(_00649_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00824_ ) );
NAND3_X1 _16625_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00825_ ) );
AND2_X1 _16626_ ( .A1(_00824_ ), .A2(_00825_ ), .ZN(_00826_ ) );
NAND3_X1 _16627_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_00827_ ) );
NAND3_X1 _16628_ ( .A1(_00657_ ), .A2(_00632_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_00828_ ) );
NAND4_X1 _16629_ ( .A1(_00826_ ), .A2(_00653_ ), .A3(_00827_ ), .A4(_00828_ ), .ZN(_00829_ ) );
NAND3_X1 _16630_ ( .A1(_00823_ ), .A2(_00623_ ), .A3(_00829_ ), .ZN(_00830_ ) );
INV_X1 _16631_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00831_ ) );
OAI21_X1 _16632_ ( .A(\myifu.state [2] ), .B1(_00609_ ), .B2(_00831_ ), .ZN(_00832_ ) );
NOR4_X1 _16633_ ( .A1(\myifu.data_in [13] ), .A2(_00669_ ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_00833_ ) );
OAI21_X1 _16634_ ( .A(_00830_ ), .B1(_00832_ ), .B2(_00833_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
OAI211_X1 _16635_ ( .A(_00598_ ), .B(_00603_ ), .C1(_06049_ ), .C2(_00501_ ), .ZN(_00834_ ) );
NAND2_X1 _16636_ ( .A1(_00834_ ), .A2(\myifu.state [2] ), .ZN(_00835_ ) );
AOI21_X1 _16637_ ( .A(_00835_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00702_ ), .ZN(_00836_ ) );
AND3_X1 _16638_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_00837_ ) );
AND3_X1 _16639_ ( .A1(_03746_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_00838_ ) );
AOI211_X1 _16640_ ( .A(_00837_ ), .B(_00838_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_06003_ ), .ZN(_00839_ ) );
NAND3_X1 _16641_ ( .A1(_00635_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_00840_ ) );
NAND4_X1 _16642_ ( .A1(_00839_ ), .A2(_00615_ ), .A3(_00617_ ), .A4(_00840_ ), .ZN(_00841_ ) );
NAND3_X1 _16643_ ( .A1(_00625_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_00842_ ) );
NAND3_X1 _16644_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_00843_ ) );
AND2_X1 _16645_ ( .A1(_00842_ ), .A2(_00843_ ), .ZN(_00844_ ) );
NAND3_X1 _16646_ ( .A1(_03755_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_00845_ ) );
NAND3_X1 _16647_ ( .A1(_03747_ ), .A2(_03755_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_00846_ ) );
NAND4_X1 _16648_ ( .A1(_00844_ ), .A2(_00653_ ), .A3(_00845_ ), .A4(_00846_ ), .ZN(_00847_ ) );
AND3_X1 _16649_ ( .A1(_00841_ ), .A2(_00622_ ), .A3(_00847_ ), .ZN(_00848_ ) );
OR2_X1 _16650_ ( .A1(_00836_ ), .A2(_00848_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
OR4_X1 _16651_ ( .A1(_00669_ ), .A2(\myifu.data_in [29] ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_00849_ ) );
AOI21_X1 _16652_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00850_ ) );
NAND2_X1 _16653_ ( .A1(_00849_ ), .A2(_00850_ ), .ZN(_00851_ ) );
AND3_X1 _16654_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_00852_ ) );
AND3_X1 _16655_ ( .A1(_00723_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_00853_ ) );
AOI211_X1 _16656_ ( .A(_00852_ ), .B(_00853_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_00790_ ), .ZN(_00854_ ) );
NAND3_X1 _16657_ ( .A1(_00792_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_00855_ ) );
NAND4_X1 _16658_ ( .A1(_00854_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00855_ ), .ZN(_00856_ ) );
NAND3_X1 _16659_ ( .A1(_00626_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_00857_ ) );
NAND3_X1 _16660_ ( .A1(fanout_net_11 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_00858_ ) );
AND2_X1 _16661_ ( .A1(_00857_ ), .A2(_00858_ ), .ZN(_00859_ ) );
NAND3_X1 _16662_ ( .A1(_00749_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_00860_ ) );
NAND3_X1 _16663_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_00861_ ) );
NAND4_X1 _16664_ ( .A1(_00859_ ), .A2(_00731_ ), .A3(_00860_ ), .A4(_00861_ ), .ZN(_00862_ ) );
NAND3_X1 _16665_ ( .A1(_00856_ ), .A2(_00624_ ), .A3(_00862_ ), .ZN(_00863_ ) );
NAND2_X1 _16666_ ( .A1(_00851_ ), .A2(_00863_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16667_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_00864_ ) );
AND3_X1 _16668_ ( .A1(_00625_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_00865_ ) );
AOI211_X1 _16669_ ( .A(_00864_ ), .B(_00865_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_06003_ ), .ZN(_00866_ ) );
NAND3_X1 _16670_ ( .A1(_00636_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_00867_ ) );
NAND4_X1 _16671_ ( .A1(_00866_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_00867_ ), .ZN(_00868_ ) );
NAND3_X1 _16672_ ( .A1(_00649_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_00869_ ) );
NAND3_X1 _16673_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_00870_ ) );
AND2_X1 _16674_ ( .A1(_00869_ ), .A2(_00870_ ), .ZN(_00871_ ) );
NAND3_X1 _16675_ ( .A1(_00632_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_00872_ ) );
NAND3_X1 _16676_ ( .A1(_00626_ ), .A2(_00632_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_00873_ ) );
NAND4_X1 _16677_ ( .A1(_00871_ ), .A2(_00653_ ), .A3(_00872_ ), .A4(_00873_ ), .ZN(_00874_ ) );
NAND3_X1 _16678_ ( .A1(_00868_ ), .A2(_00623_ ), .A3(_00874_ ), .ZN(_00875_ ) );
OAI21_X1 _16679_ ( .A(\myifu.state [2] ), .B1(_00609_ ), .B2(_03507_ ), .ZN(_00876_ ) );
NOR4_X1 _16680_ ( .A1(\myifu.data_in [11] ), .A2(_00669_ ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_00877_ ) );
OAI21_X1 _16681_ ( .A(_00875_ ), .B1(_00876_ ), .B2(_00877_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
OR4_X1 _16682_ ( .A1(_00669_ ), .A2(\myifu.data_in [10] ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_00878_ ) );
OAI211_X1 _16683_ ( .A(_00878_ ), .B(\myifu.state [2] ), .C1(_03498_ ), .C2(_00609_ ), .ZN(_00879_ ) );
AND3_X1 _16684_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_00880_ ) );
AND3_X1 _16685_ ( .A1(_00723_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_00881_ ) );
AOI211_X1 _16686_ ( .A(_00880_ ), .B(_00881_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_00790_ ), .ZN(_00882_ ) );
NAND3_X1 _16687_ ( .A1(_00792_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_00883_ ) );
NAND4_X1 _16688_ ( .A1(_00882_ ), .A2(_00616_ ), .A3(_00619_ ), .A4(_00883_ ), .ZN(_00884_ ) );
BUF_X4 _16689_ ( .A(_00625_ ), .Z(_00885_ ) );
NAND3_X1 _16690_ ( .A1(_00885_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_00886_ ) );
NAND3_X1 _16691_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_00887_ ) );
AND2_X1 _16692_ ( .A1(_00886_ ), .A2(_00887_ ), .ZN(_00888_ ) );
NAND3_X1 _16693_ ( .A1(_00749_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_00889_ ) );
NAND3_X1 _16694_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_00890_ ) );
NAND4_X1 _16695_ ( .A1(_00888_ ), .A2(_00731_ ), .A3(_00889_ ), .A4(_00890_ ), .ZN(_00891_ ) );
NAND3_X1 _16696_ ( .A1(_00884_ ), .A2(_00624_ ), .A3(_00891_ ), .ZN(_00892_ ) );
NAND2_X1 _16697_ ( .A1(_00879_ ), .A2(_00892_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
AOI21_X1 _16698_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_00893_ ) );
OAI211_X1 _16699_ ( .A(_00599_ ), .B(_00604_ ), .C1(_06050_ ), .C2(_00513_ ), .ZN(_00894_ ) );
NAND2_X1 _16700_ ( .A1(_00893_ ), .A2(_00894_ ), .ZN(_00895_ ) );
AND3_X1 _16701_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_00896_ ) );
AND3_X1 _16702_ ( .A1(_00723_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_00897_ ) );
AOI211_X1 _16703_ ( .A(_00896_ ), .B(_00897_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_00790_ ), .ZN(_00898_ ) );
BUF_X4 _16704_ ( .A(_00645_ ), .Z(_00899_ ) );
BUF_X4 _16705_ ( .A(_00617_ ), .Z(_00900_ ) );
NAND3_X1 _16706_ ( .A1(_00792_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_00901_ ) );
NAND4_X1 _16707_ ( .A1(_00898_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_00901_ ), .ZN(_00902_ ) );
NAND3_X1 _16708_ ( .A1(_00885_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_00903_ ) );
NAND3_X1 _16709_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_00904_ ) );
AND2_X1 _16710_ ( .A1(_00903_ ), .A2(_00904_ ), .ZN(_00905_ ) );
NAND3_X1 _16711_ ( .A1(_00749_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_00906_ ) );
NAND3_X1 _16712_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_00907_ ) );
NAND4_X1 _16713_ ( .A1(_00905_ ), .A2(_00731_ ), .A3(_00906_ ), .A4(_00907_ ), .ZN(_00908_ ) );
NAND3_X1 _16714_ ( .A1(_00902_ ), .A2(_00624_ ), .A3(_00908_ ), .ZN(_00909_ ) );
NAND2_X1 _16715_ ( .A1(_00895_ ), .A2(_00909_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
AOI21_X1 _16716_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00910_ ) );
NAND2_X1 _16717_ ( .A1(_00517_ ), .A2(_00519_ ), .ZN(_00911_ ) );
OAI211_X1 _16718_ ( .A(_00599_ ), .B(_00604_ ), .C1(_00911_ ), .C2(_00606_ ), .ZN(_00912_ ) );
NAND2_X1 _16719_ ( .A1(_00910_ ), .A2(_00912_ ), .ZN(_00913_ ) );
AND3_X1 _16720_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_00914_ ) );
AND3_X1 _16721_ ( .A1(_00723_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_00915_ ) );
AOI211_X1 _16722_ ( .A(_00914_ ), .B(_00915_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_00790_ ), .ZN(_00916_ ) );
NAND3_X1 _16723_ ( .A1(_00792_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_00917_ ) );
NAND4_X1 _16724_ ( .A1(_00916_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_00917_ ), .ZN(_00918_ ) );
BUF_X4 _16725_ ( .A(_00623_ ), .Z(_00919_ ) );
NAND3_X1 _16726_ ( .A1(_00885_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_00920_ ) );
NAND3_X1 _16727_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_00921_ ) );
AND2_X1 _16728_ ( .A1(_00920_ ), .A2(_00921_ ), .ZN(_00922_ ) );
NAND3_X1 _16729_ ( .A1(_00749_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_00923_ ) );
NAND3_X1 _16730_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_00924_ ) );
NAND4_X1 _16731_ ( .A1(_00922_ ), .A2(_00731_ ), .A3(_00923_ ), .A4(_00924_ ), .ZN(_00925_ ) );
NAND3_X1 _16732_ ( .A1(_00918_ ), .A2(_00919_ ), .A3(_00925_ ), .ZN(_00926_ ) );
NAND2_X1 _16733_ ( .A1(_00913_ ), .A2(_00926_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AOI21_X1 _16734_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00927_ ) );
OAI211_X1 _16735_ ( .A(_00599_ ), .B(_00604_ ), .C1(_06050_ ), .C2(_00522_ ), .ZN(_00928_ ) );
NAND2_X1 _16736_ ( .A1(_00927_ ), .A2(_00928_ ), .ZN(_00929_ ) );
AND3_X1 _16737_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_00930_ ) );
AND3_X1 _16738_ ( .A1(_00723_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_00931_ ) );
AOI211_X1 _16739_ ( .A(_00930_ ), .B(_00931_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00790_ ), .ZN(_00932_ ) );
NAND3_X1 _16740_ ( .A1(_00792_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_00933_ ) );
NAND4_X1 _16741_ ( .A1(_00932_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_00933_ ), .ZN(_00934_ ) );
NAND3_X1 _16742_ ( .A1(_00885_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_00935_ ) );
NAND3_X1 _16743_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_00936_ ) );
AND2_X1 _16744_ ( .A1(_00935_ ), .A2(_00936_ ), .ZN(_00937_ ) );
NAND3_X1 _16745_ ( .A1(_00749_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_00938_ ) );
NAND3_X1 _16746_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_00939_ ) );
NAND4_X1 _16747_ ( .A1(_00937_ ), .A2(_00731_ ), .A3(_00938_ ), .A4(_00939_ ), .ZN(_00940_ ) );
NAND3_X1 _16748_ ( .A1(_00934_ ), .A2(_00919_ ), .A3(_00940_ ), .ZN(_00941_ ) );
NAND2_X1 _16749_ ( .A1(_00929_ ), .A2(_00941_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
OAI211_X1 _16750_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00525_ ), .C2(_06049_ ), .ZN(_00942_ ) );
INV_X1 _16751_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00943_ ) );
OAI211_X1 _16752_ ( .A(_00942_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_00943_ ), .ZN(_00944_ ) );
AND3_X1 _16753_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_00945_ ) );
AND3_X1 _16754_ ( .A1(_00723_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_00946_ ) );
AOI211_X1 _16755_ ( .A(_00945_ ), .B(_00946_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00790_ ), .ZN(_00947_ ) );
NAND3_X1 _16756_ ( .A1(_00792_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_00948_ ) );
NAND4_X1 _16757_ ( .A1(_00947_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_00948_ ), .ZN(_00949_ ) );
NAND3_X1 _16758_ ( .A1(_00885_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_00950_ ) );
NAND3_X1 _16759_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_00951_ ) );
AND2_X1 _16760_ ( .A1(_00950_ ), .A2(_00951_ ), .ZN(_00952_ ) );
NAND3_X1 _16761_ ( .A1(_00749_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_00953_ ) );
NAND3_X1 _16762_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_00954_ ) );
NAND4_X1 _16763_ ( .A1(_00952_ ), .A2(_00731_ ), .A3(_00953_ ), .A4(_00954_ ), .ZN(_00955_ ) );
NAND3_X1 _16764_ ( .A1(_00949_ ), .A2(_00919_ ), .A3(_00955_ ), .ZN(_00956_ ) );
NAND2_X1 _16765_ ( .A1(_00944_ ), .A2(_00956_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
OAI211_X1 _16766_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00606_ ), .C2(_00528_ ), .ZN(_00957_ ) );
INV_X1 _16767_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00958_ ) );
OAI211_X1 _16768_ ( .A(_00957_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_00958_ ), .ZN(_00959_ ) );
AND3_X1 _16769_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_00960_ ) );
AND3_X1 _16770_ ( .A1(_00641_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_00961_ ) );
AOI211_X1 _16771_ ( .A(_00960_ ), .B(_00961_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00790_ ), .ZN(_00962_ ) );
NAND3_X1 _16772_ ( .A1(_00792_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_00963_ ) );
NAND4_X1 _16773_ ( .A1(_00962_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_00963_ ), .ZN(_00964_ ) );
NAND3_X1 _16774_ ( .A1(_00885_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_00965_ ) );
NAND3_X1 _16775_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_00966_ ) );
AND2_X1 _16776_ ( .A1(_00965_ ), .A2(_00966_ ), .ZN(_00967_ ) );
NAND3_X1 _16777_ ( .A1(_00749_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_00968_ ) );
NAND3_X1 _16778_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_00969_ ) );
NAND4_X1 _16779_ ( .A1(_00967_ ), .A2(_00654_ ), .A3(_00968_ ), .A4(_00969_ ), .ZN(_00970_ ) );
NAND3_X1 _16780_ ( .A1(_00964_ ), .A2(_00919_ ), .A3(_00970_ ), .ZN(_00971_ ) );
NAND2_X1 _16781_ ( .A1(_00959_ ), .A2(_00971_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _16782_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00972_ ) );
OAI211_X1 _16783_ ( .A(_00599_ ), .B(_00604_ ), .C1(_00531_ ), .C2(_00606_ ), .ZN(_00973_ ) );
NAND2_X1 _16784_ ( .A1(_00972_ ), .A2(_00973_ ), .ZN(_00974_ ) );
AND3_X1 _16785_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_00975_ ) );
AND3_X1 _16786_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_00976_ ) );
AOI211_X1 _16787_ ( .A(_00975_ ), .B(_00976_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00790_ ), .ZN(_00977_ ) );
NAND3_X1 _16788_ ( .A1(_00792_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_00978_ ) );
NAND4_X1 _16789_ ( .A1(_00977_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_00978_ ), .ZN(_00979_ ) );
NAND3_X1 _16790_ ( .A1(_00885_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_00980_ ) );
NAND3_X1 _16791_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_00981_ ) );
AND2_X1 _16792_ ( .A1(_00980_ ), .A2(_00981_ ), .ZN(_00982_ ) );
NAND3_X1 _16793_ ( .A1(_00646_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_00983_ ) );
NAND3_X1 _16794_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_00984_ ) );
NAND4_X1 _16795_ ( .A1(_00982_ ), .A2(_00654_ ), .A3(_00983_ ), .A4(_00984_ ), .ZN(_00985_ ) );
NAND3_X1 _16796_ ( .A1(_00979_ ), .A2(_00919_ ), .A3(_00985_ ), .ZN(_00986_ ) );
NAND2_X1 _16797_ ( .A1(_00974_ ), .A2(_00986_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
OAI211_X1 _16798_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00606_ ), .C2(_00534_ ), .ZN(_00987_ ) );
INV_X1 _16799_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00988_ ) );
OAI211_X1 _16800_ ( .A(_00987_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_00988_ ), .ZN(_00989_ ) );
AND3_X1 _16801_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_00990_ ) );
AND3_X1 _16802_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_00991_ ) );
AOI211_X1 _16803_ ( .A(_00990_ ), .B(_00991_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_00790_ ), .ZN(_00992_ ) );
NAND3_X1 _16804_ ( .A1(_00792_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_00993_ ) );
NAND4_X1 _16805_ ( .A1(_00992_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_00993_ ), .ZN(_00994_ ) );
NAND3_X1 _16806_ ( .A1(_00885_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_00995_ ) );
NAND3_X1 _16807_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_00996_ ) );
AND2_X1 _16808_ ( .A1(_00995_ ), .A2(_00996_ ), .ZN(_00997_ ) );
NAND3_X1 _16809_ ( .A1(_00646_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_00998_ ) );
NAND3_X1 _16810_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_00999_ ) );
NAND4_X1 _16811_ ( .A1(_00997_ ), .A2(_00654_ ), .A3(_00998_ ), .A4(_00999_ ), .ZN(_01000_ ) );
NAND3_X1 _16812_ ( .A1(_00994_ ), .A2(_00919_ ), .A3(_01000_ ), .ZN(_01001_ ) );
NAND2_X1 _16813_ ( .A1(_00989_ ), .A2(_01001_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
OAI211_X1 _16814_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00540_ ), .C2(_06049_ ), .ZN(_01002_ ) );
INV_X1 _16815_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01003_ ) );
OAI211_X1 _16816_ ( .A(_01002_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_01003_ ), .ZN(_01004_ ) );
AND3_X1 _16817_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01005_ ) );
AND3_X1 _16818_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01006_ ) );
AOI211_X1 _16819_ ( .A(_01005_ ), .B(_01006_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_00643_ ), .ZN(_01007_ ) );
NAND3_X1 _16820_ ( .A1(_00633_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01008_ ) );
NAND4_X1 _16821_ ( .A1(_01007_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_01008_ ), .ZN(_01009_ ) );
NAND3_X1 _16822_ ( .A1(_00885_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01010_ ) );
NAND3_X1 _16823_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01011_ ) );
AND2_X1 _16824_ ( .A1(_01010_ ), .A2(_01011_ ), .ZN(_01012_ ) );
NAND3_X1 _16825_ ( .A1(_00646_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01013_ ) );
NAND3_X1 _16826_ ( .A1(_00657_ ), .A2(_00655_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01014_ ) );
NAND4_X1 _16827_ ( .A1(_01012_ ), .A2(_00654_ ), .A3(_01013_ ), .A4(_01014_ ), .ZN(_01015_ ) );
NAND3_X1 _16828_ ( .A1(_01009_ ), .A2(_00919_ ), .A3(_01015_ ), .ZN(_01016_ ) );
NAND2_X1 _16829_ ( .A1(_01004_ ), .A2(_01016_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
OAI211_X1 _16830_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00606_ ), .C2(_00537_ ), .ZN(_01017_ ) );
OAI211_X1 _16831_ ( .A(_01017_ ), .B(\myifu.state [2] ), .C1(_00610_ ), .C2(_03523_ ), .ZN(_01018_ ) );
AND3_X1 _16832_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01019_ ) );
AND3_X1 _16833_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01020_ ) );
AOI211_X1 _16834_ ( .A(_01019_ ), .B(_01020_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00643_ ), .ZN(_01021_ ) );
NAND3_X1 _16835_ ( .A1(_00633_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01022_ ) );
NAND4_X1 _16836_ ( .A1(_01021_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_01022_ ), .ZN(_01023_ ) );
NAND3_X1 _16837_ ( .A1(_00885_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01024_ ) );
NAND3_X1 _16838_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01025_ ) );
AND2_X1 _16839_ ( .A1(_01024_ ), .A2(_01025_ ), .ZN(_01026_ ) );
NAND3_X1 _16840_ ( .A1(_00646_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01027_ ) );
NAND3_X1 _16841_ ( .A1(_00657_ ), .A2(_00655_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01028_ ) );
NAND4_X1 _16842_ ( .A1(_01026_ ), .A2(_00654_ ), .A3(_01027_ ), .A4(_01028_ ), .ZN(_01029_ ) );
NAND3_X1 _16843_ ( .A1(_01023_ ), .A2(_00919_ ), .A3(_01029_ ), .ZN(_01030_ ) );
NAND2_X1 _16844_ ( .A1(_01018_ ), .A2(_01030_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
AOI21_X1 _16845_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01031_ ) );
OAI211_X1 _16846_ ( .A(_00599_ ), .B(_00604_ ), .C1(_06050_ ), .C2(_00543_ ), .ZN(_01032_ ) );
NAND2_X1 _16847_ ( .A1(_01031_ ), .A2(_01032_ ), .ZN(_01033_ ) );
AND3_X1 _16848_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01034_ ) );
AND3_X1 _16849_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01035_ ) );
AOI211_X1 _16850_ ( .A(_01034_ ), .B(_01035_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_00643_ ), .ZN(_01036_ ) );
NAND3_X1 _16851_ ( .A1(_00633_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01037_ ) );
NAND4_X1 _16852_ ( .A1(_01036_ ), .A2(_00899_ ), .A3(_00900_ ), .A4(_01037_ ), .ZN(_01038_ ) );
NAND3_X1 _16853_ ( .A1(_00649_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01039_ ) );
NAND3_X1 _16854_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01040_ ) );
AND2_X1 _16855_ ( .A1(_01039_ ), .A2(_01040_ ), .ZN(_01041_ ) );
NAND3_X1 _16856_ ( .A1(_00646_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01042_ ) );
NAND3_X1 _16857_ ( .A1(_00657_ ), .A2(_00655_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01043_ ) );
NAND4_X1 _16858_ ( .A1(_01041_ ), .A2(_00654_ ), .A3(_01042_ ), .A4(_01043_ ), .ZN(_01044_ ) );
NAND3_X1 _16859_ ( .A1(_01038_ ), .A2(_00919_ ), .A3(_01044_ ), .ZN(_01045_ ) );
NAND2_X1 _16860_ ( .A1(_01033_ ), .A2(_01045_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
OAI211_X1 _16861_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00606_ ), .C2(_00546_ ), .ZN(_01046_ ) );
OAI211_X1 _16862_ ( .A(_01046_ ), .B(\myifu.state [2] ), .C1(_00609_ ), .C2(_03516_ ), .ZN(_01047_ ) );
AND3_X1 _16863_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01048_ ) );
AND3_X1 _16864_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01049_ ) );
AOI211_X1 _16865_ ( .A(_01048_ ), .B(_01049_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00643_ ), .ZN(_01050_ ) );
NAND3_X1 _16866_ ( .A1(_00633_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01051_ ) );
NAND4_X1 _16867_ ( .A1(_01050_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_01051_ ), .ZN(_01052_ ) );
NAND3_X1 _16868_ ( .A1(_00649_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01053_ ) );
NAND3_X1 _16869_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01054_ ) );
AND2_X1 _16870_ ( .A1(_01053_ ), .A2(_01054_ ), .ZN(_01055_ ) );
NAND3_X1 _16871_ ( .A1(_00646_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01056_ ) );
NAND3_X1 _16872_ ( .A1(_00657_ ), .A2(_00655_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01057_ ) );
NAND4_X1 _16873_ ( .A1(_01055_ ), .A2(_00654_ ), .A3(_01056_ ), .A4(_01057_ ), .ZN(_01058_ ) );
NAND3_X1 _16874_ ( .A1(_01052_ ), .A2(_00919_ ), .A3(_01058_ ), .ZN(_01059_ ) );
NAND2_X1 _16875_ ( .A1(_01047_ ), .A2(_01059_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
OAI211_X1 _16876_ ( .A(_00736_ ), .B(_00737_ ), .C1(_00606_ ), .C2(_00549_ ), .ZN(_01060_ ) );
OAI211_X1 _16877_ ( .A(_01060_ ), .B(\myifu.state [2] ), .C1(_00609_ ), .C2(_03476_ ), .ZN(_01061_ ) );
AND3_X1 _16878_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01062_ ) );
AND3_X1 _16879_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01063_ ) );
AOI211_X1 _16880_ ( .A(_01062_ ), .B(_01063_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_00643_ ), .ZN(_01064_ ) );
NAND3_X1 _16881_ ( .A1(_00633_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01065_ ) );
NAND4_X1 _16882_ ( .A1(_01064_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_01065_ ), .ZN(_01066_ ) );
NAND3_X1 _16883_ ( .A1(_00649_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01067_ ) );
NAND3_X1 _16884_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01068_ ) );
AND2_X1 _16885_ ( .A1(_01067_ ), .A2(_01068_ ), .ZN(_01069_ ) );
NAND3_X1 _16886_ ( .A1(_00646_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01070_ ) );
NAND3_X1 _16887_ ( .A1(_00657_ ), .A2(_00655_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01071_ ) );
NAND4_X1 _16888_ ( .A1(_01069_ ), .A2(_00654_ ), .A3(_01070_ ), .A4(_01071_ ), .ZN(_01072_ ) );
NAND3_X1 _16889_ ( .A1(_01066_ ), .A2(_00623_ ), .A3(_01072_ ), .ZN(_01073_ ) );
NAND2_X1 _16890_ ( .A1(_01061_ ), .A2(_01073_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
AOI21_X1 _16891_ ( .A(_00701_ ), .B1(_00703_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_01074_ ) );
OAI211_X1 _16892_ ( .A(_00599_ ), .B(_00604_ ), .C1(_00552_ ), .C2(_00606_ ), .ZN(_01075_ ) );
NAND2_X1 _16893_ ( .A1(_01074_ ), .A2(_01075_ ), .ZN(_01076_ ) );
AND3_X1 _16894_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01077_ ) );
AND3_X1 _16895_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01078_ ) );
AOI211_X1 _16896_ ( .A(_01077_ ), .B(_01078_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00643_ ), .ZN(_01079_ ) );
NAND3_X1 _16897_ ( .A1(_00633_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01080_ ) );
NAND4_X1 _16898_ ( .A1(_01079_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_01080_ ), .ZN(_01081_ ) );
NAND3_X1 _16899_ ( .A1(_00649_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01082_ ) );
NAND3_X1 _16900_ ( .A1(fanout_net_13 ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01083_ ) );
AND2_X1 _16901_ ( .A1(_01082_ ), .A2(_01083_ ), .ZN(_01084_ ) );
NAND3_X1 _16902_ ( .A1(_00646_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01085_ ) );
NAND3_X1 _16903_ ( .A1(_00657_ ), .A2(_00655_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01086_ ) );
NAND4_X1 _16904_ ( .A1(_01084_ ), .A2(_00654_ ), .A3(_01085_ ), .A4(_01086_ ), .ZN(_01087_ ) );
NAND3_X1 _16905_ ( .A1(_01081_ ), .A2(_00623_ ), .A3(_01087_ ), .ZN(_01088_ ) );
NAND2_X1 _16906_ ( .A1(_01076_ ), .A2(_01088_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
AND2_X1 _16907_ ( .A1(_00554_ ), .A2(_00555_ ), .ZN(_01089_ ) );
OAI211_X1 _16908_ ( .A(_00598_ ), .B(_00603_ ), .C1(_01089_ ), .C2(_01954_ ), .ZN(_01090_ ) );
NAND2_X1 _16909_ ( .A1(_01090_ ), .A2(\myifu.state [2] ), .ZN(_01091_ ) );
AOI21_X1 _16910_ ( .A(_01091_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00702_ ), .ZN(_01092_ ) );
AND3_X1 _16911_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01093_ ) );
AND3_X1 _16912_ ( .A1(_03746_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01094_ ) );
AOI211_X1 _16913_ ( .A(_01093_ ), .B(_01094_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_06003_ ), .ZN(_01095_ ) );
NAND3_X1 _16914_ ( .A1(_00635_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01096_ ) );
NAND4_X1 _16915_ ( .A1(_01095_ ), .A2(_00615_ ), .A3(_00617_ ), .A4(_01096_ ), .ZN(_01097_ ) );
NAND3_X1 _16916_ ( .A1(_03746_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01098_ ) );
NAND3_X1 _16917_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01099_ ) );
AND2_X1 _16918_ ( .A1(_01098_ ), .A2(_01099_ ), .ZN(_01100_ ) );
NAND3_X1 _16919_ ( .A1(_03755_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01101_ ) );
NAND3_X1 _16920_ ( .A1(_03747_ ), .A2(_03755_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01102_ ) );
NAND4_X1 _16921_ ( .A1(_01100_ ), .A2(_00653_ ), .A3(_01101_ ), .A4(_01102_ ), .ZN(_01103_ ) );
AND3_X1 _16922_ ( .A1(_01097_ ), .A2(_00622_ ), .A3(_01103_ ), .ZN(_01104_ ) );
OR2_X1 _16923_ ( .A1(_01092_ ), .A2(_01104_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
OAI211_X1 _16924_ ( .A(_00598_ ), .B(_00603_ ), .C1(_06049_ ), .C2(_00558_ ), .ZN(_01105_ ) );
NAND2_X1 _16925_ ( .A1(_01105_ ), .A2(\myifu.state [2] ), .ZN(_01106_ ) );
AOI21_X1 _16926_ ( .A(_01106_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00702_ ), .ZN(_01107_ ) );
AND3_X1 _16927_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01108_ ) );
AND3_X1 _16928_ ( .A1(_03746_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01109_ ) );
AOI211_X1 _16929_ ( .A(_01108_ ), .B(_01109_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_06003_ ), .ZN(_01110_ ) );
NAND3_X1 _16930_ ( .A1(_00635_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01111_ ) );
NAND4_X1 _16931_ ( .A1(_01110_ ), .A2(_00615_ ), .A3(_00617_ ), .A4(_01111_ ), .ZN(_01112_ ) );
NAND3_X1 _16932_ ( .A1(_03746_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01113_ ) );
NAND3_X1 _16933_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01114_ ) );
AND2_X1 _16934_ ( .A1(_01113_ ), .A2(_01114_ ), .ZN(_01115_ ) );
NAND3_X1 _16935_ ( .A1(_03755_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01116_ ) );
NAND3_X1 _16936_ ( .A1(_03747_ ), .A2(_03755_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01117_ ) );
NAND4_X1 _16937_ ( .A1(_01115_ ), .A2(_00630_ ), .A3(_01116_ ), .A4(_01117_ ), .ZN(_01118_ ) );
AND3_X1 _16938_ ( .A1(_01112_ ), .A2(_00622_ ), .A3(_01118_ ), .ZN(_01119_ ) );
OR2_X1 _16939_ ( .A1(_01107_ ), .A2(_01119_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
AND3_X1 _16940_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01120_ ) );
AND3_X1 _16941_ ( .A1(_00625_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01121_ ) );
AOI211_X1 _16942_ ( .A(_01120_ ), .B(_01121_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_06003_ ), .ZN(_01122_ ) );
NAND3_X1 _16943_ ( .A1(_00636_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01123_ ) );
NAND4_X1 _16944_ ( .A1(_01122_ ), .A2(_00645_ ), .A3(_00618_ ), .A4(_01123_ ), .ZN(_01124_ ) );
NAND3_X1 _16945_ ( .A1(_00649_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01125_ ) );
NAND3_X1 _16946_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01126_ ) );
AND2_X1 _16947_ ( .A1(_01125_ ), .A2(_01126_ ), .ZN(_01127_ ) );
NAND3_X1 _16948_ ( .A1(_00632_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01128_ ) );
NAND3_X1 _16949_ ( .A1(_00626_ ), .A2(_00632_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01129_ ) );
NAND4_X1 _16950_ ( .A1(_01127_ ), .A2(_00653_ ), .A3(_01128_ ), .A4(_01129_ ), .ZN(_01130_ ) );
NAND3_X1 _16951_ ( .A1(_01124_ ), .A2(_00623_ ), .A3(_01130_ ), .ZN(_01131_ ) );
INV_X1 _16952_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_01132_ ) );
OAI21_X1 _16953_ ( .A(\myifu.state [2] ), .B1(_00609_ ), .B2(_01132_ ), .ZN(_01133_ ) );
NOR4_X1 _16954_ ( .A1(\myifu.data_in [22] ), .A2(_00669_ ), .A3(_00602_ ), .A4(_00601_ ), .ZN(_01134_ ) );
OAI21_X1 _16955_ ( .A(_01131_ ), .B1(_01133_ ), .B2(_01134_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI21_X1 _16956_ ( .A(_03749_ ), .B1(_03630_ ), .B2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _16957_ ( .A1(_03819_ ), .A2(_03821_ ), .A3(_03830_ ), .A4(\myifu.state [2] ), .ZN(_01135_ ) );
INV_X1 _16958_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01136_ ) );
AND4_X1 _16959_ ( .A1(_01136_ ), .A2(_01869_ ), .A3(\myifu.state [0] ), .A4(_01933_ ), .ZN(_01137_ ) );
NOR2_X1 _16960_ ( .A1(_01137_ ), .A2(_00451_ ), .ZN(_01138_ ) );
AOI21_X1 _16961_ ( .A(reset ), .B1(_01135_ ), .B2(_01138_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _16962_ ( .A1(_05992_ ), .A2(_02027_ ), .ZN(_01139_ ) );
NAND3_X1 _16963_ ( .A1(_01139_ ), .A2(_01136_ ), .A3(_01967_ ), .ZN(_01140_ ) );
OAI211_X1 _16964_ ( .A(_01140_ ), .B(_03744_ ), .C1(_01136_ ), .C2(_01935_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _16965_ ( .A1(_03831_ ), .A2(_01570_ ), .A3(\myifu.state [2] ), .ZN(_01141_ ) );
NAND3_X1 _16966_ ( .A1(_05992_ ), .A2(\io_master_arburst [0] ), .A3(_02064_ ), .ZN(_01142_ ) );
NAND2_X1 _16967_ ( .A1(_01141_ ), .A2(_01142_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _16968_ ( .A1(_03819_ ), .A2(\myifu.state [2] ), .A3(_03830_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
NOR4_X1 _16969_ ( .A1(_00631_ ), .A2(_02063_ ), .A3(_06007_ ), .A4(_06008_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NOR4_X1 _16970_ ( .A1(_00631_ ), .A2(_02063_ ), .A3(_06007_ ), .A4(_00562_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _16971_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00631_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _16972_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(_03756_ ), .A4(_00631_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _16973_ ( .A1(_00631_ ), .A2(_02063_ ), .A3(_06006_ ), .A4(_06005_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _16974_ ( .A1(_03748_ ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00631_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
AND3_X1 _16975_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06004_ ), .A3(_00631_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _16976_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06004_ ), .A3(_00616_ ), .A4(_00619_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
NOR3_X1 _16977_ ( .A1(_02063_ ), .A2(_06005_ ), .A3(_06007_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
NOR3_X1 _16978_ ( .A1(_02063_ ), .A2(_06008_ ), .A3(_06007_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
NOR3_X1 _16979_ ( .A1(_02063_ ), .A2(_06007_ ), .A3(_00562_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
AND3_X1 _16980_ ( .A1(_02062_ ), .A2(_06004_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
AND2_X1 _16981_ ( .A1(_01934_ ), .A2(\myifu.state [0] ), .ZN(_01143_ ) );
INV_X1 _16982_ ( .A(_01143_ ), .ZN(_01144_ ) );
AOI21_X1 _16983_ ( .A(_00451_ ), .B1(\myidu.stall_quest_fencei ), .B2(\myifu.state [0] ), .ZN(_01145_ ) );
AND2_X1 _16984_ ( .A1(_00453_ ), .A2(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01146_ ) );
INV_X1 _16985_ ( .A(_01146_ ), .ZN(_01147_ ) );
NAND4_X1 _16986_ ( .A1(_01144_ ), .A2(_03215_ ), .A3(_01145_ ), .A4(_01147_ ), .ZN(_01148_ ) );
AOI221_X4 _16987_ ( .A(_01148_ ), .B1(_03831_ ), .B2(_01968_ ), .C1(_01139_ ), .C2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _16988_ ( .A1(_03618_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03215_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _16989_ ( .A(_00434_ ), .B(_00436_ ), .C1(_03075_ ), .C2(_03116_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
NAND4_X1 _16990_ ( .A1(_01147_ ), .A2(_01145_ ), .A3(_01535_ ), .A4(_03215_ ), .ZN(_01149_ ) );
INV_X1 _16991_ ( .A(_01934_ ), .ZN(_01150_ ) );
AOI21_X1 _16992_ ( .A(_01149_ ), .B1(_01150_ ), .B2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _16993_ ( .A(_06096_ ), .B(_03899_ ), .S(\mylsu.state [0] ), .Z(_01151_ ) );
NOR2_X1 _16994_ ( .A1(_06100_ ), .A2(_01151_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ) );
NOR3_X1 _16995_ ( .A1(_06100_ ), .A2(_03907_ ), .A3(_01151_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
AND3_X1 _16996_ ( .A1(_03897_ ), .A2(_02039_ ), .A3(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_01152_ ) );
NAND4_X1 _16997_ ( .A1(_05992_ ), .A2(\io_master_arid [1] ), .A3(_02048_ ), .A4(_01152_ ), .ZN(_01153_ ) );
AND2_X1 _16998_ ( .A1(_06099_ ), .A2(_03830_ ), .ZN(_01154_ ) );
OAI21_X1 _16999_ ( .A(_01153_ ), .B1(_01154_ ), .B2(_06029_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
BUF_X2 _17000_ ( .A(_02051_ ), .Z(_01155_ ) );
OAI211_X1 _17001_ ( .A(_01155_ ), .B(_06059_ ), .C1(io_master_wready ), .C2(io_master_awready ), .ZN(_01156_ ) );
NOR4_X1 _17002_ ( .A1(_02052_ ), .A2(_01156_ ), .A3(_02058_ ), .A4(_03906_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
INV_X1 _17003_ ( .A(io_master_wready ), .ZN(_01157_ ) );
NAND4_X1 _17004_ ( .A1(_03902_ ), .A2(\mylsu.state [2] ), .A3(_03904_ ), .A4(_01157_ ), .ZN(_01158_ ) );
AND3_X1 _17005_ ( .A1(_03894_ ), .A2(io_master_awready ), .A3(_03895_ ), .ZN(_01159_ ) );
AND3_X1 _17006_ ( .A1(_01159_ ), .A2(_01155_ ), .A3(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_01160_ ) );
INV_X1 _17007_ ( .A(_03846_ ), .ZN(_01161_ ) );
OAI211_X1 _17008_ ( .A(_01160_ ), .B(_01161_ ), .C1(_01157_ ), .C2(_05998_ ), .ZN(_01162_ ) );
OAI21_X1 _17009_ ( .A(_01158_ ), .B1(_02084_ ), .B2(_01162_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
AND2_X1 _17010_ ( .A1(_03896_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
AND2_X1 _17011_ ( .A1(_06010_ ), .A2(_02051_ ), .ZN(_01163_ ) );
AND2_X1 _17012_ ( .A1(_01163_ ), .A2(\mylsu.state [0] ), .ZN(_01164_ ) );
NAND4_X1 _17013_ ( .A1(_01164_ ), .A2(_02059_ ), .A3(io_master_wready ), .A4(io_master_awready ), .ZN(_01165_ ) );
NAND3_X1 _17014_ ( .A1(_03897_ ), .A2(\mylsu.state [2] ), .A3(io_master_wready ), .ZN(_01166_ ) );
NAND2_X1 _17015_ ( .A1(_01159_ ), .A2(\mylsu.state [4] ), .ZN(_01167_ ) );
NAND3_X1 _17016_ ( .A1(_06107_ ), .A2(\mylsu.state [1] ), .A3(_03897_ ), .ZN(_01168_ ) );
NAND4_X1 _17017_ ( .A1(_01165_ ), .A2(_01166_ ), .A3(_01167_ ), .A4(_01168_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
NOR3_X1 _17018_ ( .A1(_05993_ ), .A2(_02083_ ), .A3(_03846_ ), .ZN(_01169_ ) );
INV_X1 _17019_ ( .A(_02047_ ), .ZN(_01170_ ) );
NOR2_X1 _17020_ ( .A1(_02042_ ), .A2(_01170_ ), .ZN(_01171_ ) );
OAI21_X1 _17021_ ( .A(_01152_ ), .B1(_01169_ ), .B2(_01171_ ), .ZN(_01172_ ) );
OAI211_X1 _17022_ ( .A(_01164_ ), .B(_02052_ ), .C1(_02057_ ), .C2(_02055_ ), .ZN(_01173_ ) );
AOI22_X1 _17023_ ( .A1(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .A2(_03846_ ), .B1(\mylsu.state [1] ), .B2(_06106_ ), .ZN(_01174_ ) );
AND3_X1 _17024_ ( .A1(_03836_ ), .A2(_03896_ ), .A3(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_01175_ ) );
NAND3_X1 _17025_ ( .A1(_01175_ ), .A2(_02040_ ), .A3(_01161_ ), .ZN(_01176_ ) );
AND4_X1 _17026_ ( .A1(_03896_ ), .A2(_01173_ ), .A3(_01174_ ), .A4(_01176_ ), .ZN(_01177_ ) );
OR4_X1 _17027_ ( .A1(\EX_LS_typ [4] ), .A2(_06021_ ), .A3(_05996_ ), .A4(_06002_ ), .ZN(_01178_ ) );
NOR4_X1 _17028_ ( .A1(_03846_ ), .A2(_05996_ ), .A3(io_master_wready ), .A4(io_master_awready ), .ZN(_01179_ ) );
AND3_X1 _17029_ ( .A1(_01179_ ), .A2(_01155_ ), .A3(_06001_ ), .ZN(_01180_ ) );
NAND2_X1 _17030_ ( .A1(_02059_ ), .A2(_01180_ ), .ZN(_01181_ ) );
NAND4_X1 _17031_ ( .A1(_02058_ ), .A2(_06010_ ), .A3(\mylsu.state [0] ), .A4(_01155_ ), .ZN(_01182_ ) );
NAND4_X1 _17032_ ( .A1(_01177_ ), .A2(_01178_ ), .A3(_01181_ ), .A4(_01182_ ), .ZN(_01183_ ) );
AOI21_X1 _17033_ ( .A(_01183_ ), .B1(\mylsu.state [0] ), .B2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01184_ ) );
NAND3_X1 _17034_ ( .A1(_06099_ ), .A2(_03830_ ), .A3(_00283_ ), .ZN(_01185_ ) );
NAND3_X1 _17035_ ( .A1(_01172_ ), .A2(_01184_ ), .A3(_01185_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND4_X1 _17036_ ( .A1(_01155_ ), .A2(_03897_ ), .A3(_06009_ ), .A4(_05998_ ), .ZN(_01186_ ) );
NOR4_X1 _17037_ ( .A1(_01186_ ), .A2(_05996_ ), .A3(_01157_ ), .A4(_03846_ ), .ZN(_01187_ ) );
NAND2_X1 _17038_ ( .A1(_02059_ ), .A2(_01187_ ), .ZN(_01188_ ) );
NAND4_X1 _17039_ ( .A1(_03902_ ), .A2(\mylsu.state [4] ), .A3(_03904_ ), .A4(_05998_ ), .ZN(_01189_ ) );
NAND2_X1 _17040_ ( .A1(_01188_ ), .A2(_01189_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
MUX2_X1 _17041_ ( .A(\LS_WB_wdata_csreg [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_05879_ ), .Z(_01190_ ) );
INV_X1 _17042_ ( .A(_03847_ ), .ZN(_01191_ ) );
OR2_X1 _17043_ ( .A1(_03837_ ), .A2(_01191_ ), .ZN(_01192_ ) );
BUF_X4 _17044_ ( .A(_01192_ ), .Z(_01193_ ) );
BUF_X4 _17045_ ( .A(_01193_ ), .Z(_01194_ ) );
MUX2_X1 _17046_ ( .A(_01190_ ), .B(\EX_LS_pc [21] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
NAND2_X1 _17047_ ( .A1(\EX_LS_flag [2] ), .A2(\EX_LS_result_csreg_mem [20] ), .ZN(_01195_ ) );
OAI21_X1 _17048_ ( .A(_01195_ ), .B1(_03841_ ), .B2(_02079_ ), .ZN(_01196_ ) );
MUX2_X1 _17049_ ( .A(_01196_ ), .B(\EX_LS_pc [20] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
AOI21_X1 _17050_ ( .A(\EX_LS_pc [19] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01197_ ) );
MUX2_X1 _17051_ ( .A(\LS_WB_wdata_csreg [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_05736_ ), .Z(_01198_ ) );
NOR3_X1 _17052_ ( .A1(_03837_ ), .A2(_01191_ ), .A3(_01198_ ), .ZN(_01199_ ) );
NOR2_X1 _17053_ ( .A1(_01197_ ), .A2(_01199_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
AOI221_X4 _17054_ ( .A(_01193_ ), .B1(\LS_WB_wdata_csreg [18] ), .B2(_05387_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [18] ), .ZN(_01200_ ) );
AOI21_X1 _17055_ ( .A(\EX_LS_pc [18] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01201_ ) );
NOR2_X1 _17056_ ( .A1(_01200_ ), .A2(_01201_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
AOI21_X1 _17057_ ( .A(\EX_LS_pc [17] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01202_ ) );
MUX2_X1 _17058_ ( .A(\LS_WB_wdata_csreg [17] ), .B(\EX_LS_result_csreg_mem [17] ), .S(_05736_ ), .Z(_01203_ ) );
NOR3_X1 _17059_ ( .A1(_03837_ ), .A2(_01191_ ), .A3(_01203_ ), .ZN(_01204_ ) );
NOR2_X1 _17060_ ( .A1(_01202_ ), .A2(_01204_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _17061_ ( .A(\EX_LS_pc [16] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01205_ ) );
BUF_X4 _17062_ ( .A(_05232_ ), .Z(_01206_ ) );
OAI21_X1 _17063_ ( .A(_03848_ ), .B1(_01206_ ), .B2(_06138_ ), .ZN(_01207_ ) );
AOI221_X4 _17064_ ( .A(_01207_ ), .B1(\LS_WB_wdata_csreg [16] ), .B2(_01206_ ), .C1(_02084_ ), .C2(_01155_ ), .ZN(_01208_ ) );
NOR2_X1 _17065_ ( .A1(_01205_ ), .A2(_01208_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
AOI221_X4 _17066_ ( .A(_01193_ ), .B1(\LS_WB_wdata_csreg [15] ), .B2(_05387_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [15] ), .ZN(_01209_ ) );
AOI21_X1 _17067_ ( .A(\EX_LS_pc [15] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01210_ ) );
NOR2_X1 _17068_ ( .A1(_01209_ ), .A2(_01210_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _17069_ ( .A(\EX_LS_pc [14] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01211_ ) );
MUX2_X1 _17070_ ( .A(\LS_WB_wdata_csreg [14] ), .B(\EX_LS_result_csreg_mem [14] ), .S(_05736_ ), .Z(_01212_ ) );
NOR3_X1 _17071_ ( .A1(_03837_ ), .A2(_01191_ ), .A3(_01212_ ), .ZN(_01213_ ) );
NOR2_X1 _17072_ ( .A1(_01211_ ), .A2(_01213_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _17073_ ( .A(\LS_WB_wdata_csreg [13] ), .B(\EX_LS_result_csreg_mem [13] ), .S(_05879_ ), .Z(_01214_ ) );
MUX2_X1 _17074_ ( .A(_01214_ ), .B(\EX_LS_pc [13] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _17075_ ( .A(\LS_WB_wdata_csreg [12] ), .B(\EX_LS_result_csreg_mem [12] ), .S(_05879_ ), .Z(_01215_ ) );
MUX2_X1 _17076_ ( .A(_01215_ ), .B(\EX_LS_pc [12] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _17077_ ( .A(\EX_LS_pc [30] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01216_ ) );
MUX2_X1 _17078_ ( .A(\LS_WB_wdata_csreg [30] ), .B(\EX_LS_result_csreg_mem [30] ), .S(_03840_ ), .Z(_01217_ ) );
NOR3_X1 _17079_ ( .A1(_03837_ ), .A2(_01191_ ), .A3(_01217_ ), .ZN(_01218_ ) );
NOR2_X1 _17080_ ( .A1(_01216_ ), .A2(_01218_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _17081_ ( .A(\LS_WB_wdata_csreg [11] ), .B(\EX_LS_result_csreg_mem [11] ), .S(_05879_ ), .Z(_01219_ ) );
MUX2_X1 _17082_ ( .A(_01219_ ), .B(\EX_LS_pc [11] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _17083_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_05879_ ), .Z(_01220_ ) );
MUX2_X1 _17084_ ( .A(_01220_ ), .B(\EX_LS_pc [10] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _17085_ ( .A(\LS_WB_wdata_csreg [9] ), .B(\EX_LS_result_csreg_mem [9] ), .S(_05879_ ), .Z(_01221_ ) );
MUX2_X1 _17086_ ( .A(_01221_ ), .B(\EX_LS_pc [9] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _17087_ ( .A(\EX_LS_pc [8] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01222_ ) );
OAI21_X1 _17088_ ( .A(_03847_ ), .B1(_01206_ ), .B2(_06139_ ), .ZN(_01223_ ) );
AOI221_X4 _17089_ ( .A(_01223_ ), .B1(\LS_WB_wdata_csreg [8] ), .B2(_01206_ ), .C1(_02084_ ), .C2(_01155_ ), .ZN(_01224_ ) );
NOR2_X1 _17090_ ( .A1(_01222_ ), .A2(_01224_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _17091_ ( .A(\LS_WB_wdata_csreg [7] ), .B(\EX_LS_result_csreg_mem [7] ), .S(_05879_ ), .Z(_01225_ ) );
MUX2_X1 _17092_ ( .A(_01225_ ), .B(\EX_LS_pc [7] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _17093_ ( .A1(_03841_ ), .A2(_02081_ ), .B1(_03855_ ), .B2(_05719_ ), .ZN(_01226_ ) );
MUX2_X1 _17094_ ( .A(_01226_ ), .B(\EX_LS_pc [6] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
AOI21_X1 _17095_ ( .A(\EX_LS_pc [5] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01227_ ) );
OAI21_X1 _17096_ ( .A(_03847_ ), .B1(_01206_ ), .B2(_06111_ ), .ZN(_01228_ ) );
AOI221_X4 _17097_ ( .A(_01228_ ), .B1(\LS_WB_wdata_csreg [5] ), .B2(_01206_ ), .C1(_02084_ ), .C2(_01155_ ), .ZN(_01229_ ) );
NOR2_X1 _17098_ ( .A1(_01227_ ), .A2(_01229_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _17099_ ( .A(\LS_WB_wdata_csreg [4] ), .B(\EX_LS_result_csreg_mem [4] ), .S(_05879_ ), .Z(_01230_ ) );
MUX2_X1 _17100_ ( .A(_01230_ ), .B(\EX_LS_pc [4] ), .S(_01194_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
AOI21_X1 _17101_ ( .A(\EX_LS_pc [3] ), .B1(_03839_ ), .B2(_03849_ ), .ZN(_01231_ ) );
OAI21_X1 _17102_ ( .A(_03847_ ), .B1(_01206_ ), .B2(_06113_ ), .ZN(_01232_ ) );
AOI221_X4 _17103_ ( .A(_01232_ ), .B1(\LS_WB_wdata_csreg [3] ), .B2(_01206_ ), .C1(_02084_ ), .C2(_01155_ ), .ZN(_01233_ ) );
NOR2_X1 _17104_ ( .A1(_01231_ ), .A2(_01233_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
MUX2_X1 _17105_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\EX_LS_result_csreg_mem [2] ), .S(_05736_ ), .Z(_01234_ ) );
MUX2_X1 _17106_ ( .A(_01234_ ), .B(\EX_LS_pc [2] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _17107_ ( .A(\LS_WB_wdata_csreg [29] ), .B(\EX_LS_result_csreg_mem [29] ), .S(_05736_ ), .Z(_01235_ ) );
MUX2_X1 _17108_ ( .A(_01235_ ), .B(\EX_LS_pc [29] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _17109_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\EX_LS_result_csreg_mem [1] ), .S(_05736_ ), .Z(_01236_ ) );
MUX2_X1 _17110_ ( .A(_01236_ ), .B(\EX_LS_pc [1] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI221_X4 _17111_ ( .A(_01193_ ), .B1(_01941_ ), .B2(\LS_WB_wdata_csreg [0] ), .C1(\EX_LS_result_csreg_mem [0] ), .C2(_03841_ ), .ZN(_01237_ ) );
AOI21_X1 _17112_ ( .A(\EX_LS_pc [0] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01238_ ) );
NOR2_X1 _17113_ ( .A1(_01237_ ), .A2(_01238_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
AOI21_X1 _17114_ ( .A(\EX_LS_pc [28] ), .B1(_03838_ ), .B2(_03849_ ), .ZN(_01239_ ) );
OAI21_X1 _17115_ ( .A(_03847_ ), .B1(_05232_ ), .B2(_05618_ ), .ZN(_01240_ ) );
AOI221_X4 _17116_ ( .A(_01240_ ), .B1(\LS_WB_wdata_csreg [28] ), .B2(_01206_ ), .C1(_02084_ ), .C2(_01155_ ), .ZN(_01241_ ) );
NOR2_X1 _17117_ ( .A1(_01239_ ), .A2(_01241_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _17118_ ( .A(\LS_WB_wdata_csreg [27] ), .B(\EX_LS_result_csreg_mem [27] ), .S(_05736_ ), .Z(_01242_ ) );
MUX2_X1 _17119_ ( .A(_01242_ ), .B(\EX_LS_pc [27] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI21_X1 _17120_ ( .A(\EX_LS_pc [26] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01243_ ) );
MUX2_X1 _17121_ ( .A(\LS_WB_wdata_csreg [26] ), .B(\EX_LS_result_csreg_mem [26] ), .S(_03840_ ), .Z(_01244_ ) );
NOR3_X1 _17122_ ( .A1(_03837_ ), .A2(_01191_ ), .A3(_01244_ ), .ZN(_01245_ ) );
NOR2_X1 _17123_ ( .A1(_01243_ ), .A2(_01245_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI221_X4 _17124_ ( .A(_01193_ ), .B1(\LS_WB_wdata_csreg [25] ), .B2(_01941_ ), .C1(\EX_LS_result_csreg_mem [25] ), .C2(_03841_ ), .ZN(_01246_ ) );
AOI21_X1 _17125_ ( .A(\EX_LS_pc [25] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01247_ ) );
NOR2_X1 _17126_ ( .A1(_01246_ ), .A2(_01247_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI221_X4 _17127_ ( .A(_01192_ ), .B1(\LS_WB_wdata_csreg [24] ), .B2(_05387_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [24] ), .ZN(_01248_ ) );
AOI21_X1 _17128_ ( .A(\EX_LS_pc [24] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01249_ ) );
NOR2_X1 _17129_ ( .A1(_01248_ ), .A2(_01249_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _17130_ ( .A(\EX_LS_pc [23] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01250_ ) );
MUX2_X1 _17131_ ( .A(\LS_WB_wdata_csreg [23] ), .B(\EX_LS_result_csreg_mem [23] ), .S(_03840_ ), .Z(_01251_ ) );
NOR3_X1 _17132_ ( .A1(_03837_ ), .A2(_01191_ ), .A3(_01251_ ), .ZN(_01252_ ) );
NOR2_X1 _17133_ ( .A1(_01250_ ), .A2(_01252_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
AOI221_X4 _17134_ ( .A(_01192_ ), .B1(\LS_WB_wdata_csreg [22] ), .B2(_01206_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [22] ), .ZN(_01253_ ) );
AOI21_X1 _17135_ ( .A(\EX_LS_pc [22] ), .B1(_03838_ ), .B2(_03848_ ), .ZN(_01254_ ) );
NOR2_X1 _17136_ ( .A1(_01253_ ), .A2(_01254_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _17137_ ( .A(\LS_WB_wdata_csreg [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_05736_ ), .Z(_01255_ ) );
MUX2_X1 _17138_ ( .A(_01255_ ), .B(\EX_LS_pc [31] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17139_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01256_ ) );
INV_X1 _17140_ ( .A(_01256_ ), .ZN(_01257_ ) );
BUF_X2 _17141_ ( .A(_01257_ ), .Z(_01258_ ) );
OR3_X1 _17142_ ( .A1(_00491_ ), .A2(_06037_ ), .A3(_01258_ ), .ZN(_01259_ ) );
NAND3_X1 _17143_ ( .A1(_00457_ ), .A2(_01975_ ), .A3(_01258_ ), .ZN(_01260_ ) );
AND2_X2 _17144_ ( .A1(_01259_ ), .A2(_01260_ ), .ZN(_01261_ ) );
AND2_X1 _17145_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01262_ ) );
BUF_X2 _17146_ ( .A(_01262_ ), .Z(_01263_ ) );
INV_X1 _17147_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01264_ ) );
AND2_X1 _17148_ ( .A1(_01263_ ), .A2(_01264_ ), .ZN(_01265_ ) );
BUF_X2 _17149_ ( .A(_01265_ ), .Z(_01266_ ) );
AND2_X1 _17150_ ( .A1(_01261_ ), .A2(_01266_ ), .ZN(_01267_ ) );
AND2_X1 _17151_ ( .A1(_01264_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01268_ ) );
INV_X1 _17152_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_01269_ ) );
AND2_X1 _17153_ ( .A1(_01268_ ), .A2(_01269_ ), .ZN(_01270_ ) );
NAND2_X1 _17154_ ( .A1(_01269_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01271_ ) );
NOR2_X1 _17155_ ( .A1(_01271_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01272_ ) );
OR2_X1 _17156_ ( .A1(_01270_ ), .A2(_01272_ ), .ZN(_01273_ ) );
NOR2_X4 _17157_ ( .A1(_01267_ ), .A2(_01273_ ), .ZN(_01274_ ) );
AND2_X2 _17158_ ( .A1(_01262_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01275_ ) );
AOI211_X1 _17159_ ( .A(_06040_ ), .B(_01275_ ), .C1(_00464_ ), .C2(_00465_ ), .ZN(_01276_ ) );
OAI21_X1 _17160_ ( .A(_01274_ ), .B1(_01276_ ), .B2(_01266_ ), .ZN(_01277_ ) );
NOR2_X1 _17161_ ( .A1(_00491_ ), .A2(_06038_ ), .ZN(_01278_ ) );
NOR2_X1 _17162_ ( .A1(_06045_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01279_ ) );
NOR2_X1 _17163_ ( .A1(_00558_ ), .A2(_06038_ ), .ZN(_01280_ ) );
NOR2_X1 _17164_ ( .A1(_06042_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01281_ ) );
AOI22_X1 _17165_ ( .A1(_01278_ ), .A2(_01279_ ), .B1(_01280_ ), .B2(_01281_ ), .ZN(_01282_ ) );
NOR3_X1 _17166_ ( .A1(_00911_ ), .A2(_06038_ ), .A3(_01258_ ), .ZN(_01283_ ) );
INV_X1 _17167_ ( .A(_01283_ ), .ZN(_01284_ ) );
NAND4_X1 _17168_ ( .A1(_00457_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_01975_ ), .ZN(_01285_ ) );
AND3_X2 _17169_ ( .A1(_01282_ ), .A2(_01284_ ), .A3(_01285_ ), .ZN(_01286_ ) );
INV_X1 _17170_ ( .A(_01270_ ), .ZN(_01287_ ) );
NOR2_X1 _17171_ ( .A1(_01286_ ), .A2(_01287_ ), .ZN(_01288_ ) );
NOR2_X1 _17172_ ( .A1(_01288_ ), .A2(_06096_ ), .ZN(_01289_ ) );
AOI22_X1 _17173_ ( .A1(_01277_ ), .A2(_01289_ ), .B1(_06096_ ), .B2(_04474_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
INV_X1 _17174_ ( .A(_01275_ ), .ZN(_01290_ ) );
AND2_X2 _17175_ ( .A1(_01274_ ), .A2(_01290_ ), .ZN(_01291_ ) );
NOR2_X2 _17176_ ( .A1(_00471_ ), .A2(_06036_ ), .ZN(_01292_ ) );
OAI21_X1 _17177_ ( .A(_01291_ ), .B1(_01263_ ), .B2(_01292_ ), .ZN(_01293_ ) );
INV_X1 _17178_ ( .A(_01288_ ), .ZN(_01294_ ) );
BUF_X4 _17179_ ( .A(_01294_ ), .Z(_01295_ ) );
NAND2_X1 _17180_ ( .A1(_01293_ ), .A2(_01295_ ), .ZN(_01296_ ) );
MUX2_X1 _17181_ ( .A(\EX_LS_result_reg [20] ), .B(_01296_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
INV_X1 _17182_ ( .A(_01274_ ), .ZN(_01297_ ) );
NOR2_X2 _17183_ ( .A1(_00475_ ), .A2(_06037_ ), .ZN(_01298_ ) );
AOI21_X1 _17184_ ( .A(_01266_ ), .B1(_01298_ ), .B2(_01290_ ), .ZN(_01299_ ) );
OAI21_X1 _17185_ ( .A(_01294_ ), .B1(_01297_ ), .B2(_01299_ ), .ZN(_01300_ ) );
MUX2_X1 _17186_ ( .A(\EX_LS_result_reg [19] ), .B(_01300_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NOR2_X1 _17187_ ( .A1(_00478_ ), .A2(_06036_ ), .ZN(_01301_ ) );
OAI21_X1 _17188_ ( .A(_01291_ ), .B1(_01263_ ), .B2(_01301_ ), .ZN(_01302_ ) );
NAND2_X1 _17189_ ( .A1(_01302_ ), .A2(_01295_ ), .ZN(_01303_ ) );
MUX2_X1 _17190_ ( .A(\EX_LS_result_reg [18] ), .B(_01303_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NOR2_X2 _17191_ ( .A1(_00481_ ), .A2(_06037_ ), .ZN(_01304_ ) );
AOI21_X1 _17192_ ( .A(_01266_ ), .B1(_01304_ ), .B2(_01290_ ), .ZN(_01305_ ) );
OAI21_X1 _17193_ ( .A(_01294_ ), .B1(_01297_ ), .B2(_01305_ ), .ZN(_01306_ ) );
MUX2_X1 _17194_ ( .A(\EX_LS_result_reg [17] ), .B(_01306_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
AND4_X1 _17195_ ( .A1(\io_master_arid [1] ), .A2(_00484_ ), .A3(_00488_ ), .A4(_01290_ ), .ZN(_01307_ ) );
OAI21_X1 _17196_ ( .A(_01274_ ), .B1(_01266_ ), .B2(_01307_ ), .ZN(_01308_ ) );
NAND2_X1 _17197_ ( .A1(_01308_ ), .A2(_01295_ ), .ZN(_01309_ ) );
MUX2_X1 _17198_ ( .A(\EX_LS_result_reg [16] ), .B(_01309_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
INV_X1 _17199_ ( .A(_01262_ ), .ZN(_01310_ ) );
AOI21_X1 _17200_ ( .A(_01310_ ), .B1(_01259_ ), .B2(_01260_ ), .ZN(_01311_ ) );
NOR3_X1 _17201_ ( .A1(_01270_ ), .A2(_01263_ ), .A3(_01272_ ), .ZN(_01312_ ) );
AOI21_X1 _17202_ ( .A(_01311_ ), .B1(_01278_ ), .B2(_01312_ ), .ZN(_01313_ ) );
AOI22_X1 _17203_ ( .A1(_01289_ ), .A2(_01313_ ), .B1(_06096_ ), .B2(_04597_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
BUF_X4 _17204_ ( .A(_01256_ ), .Z(_01314_ ) );
NOR2_X1 _17205_ ( .A1(_01310_ ), .A2(_01314_ ), .ZN(_01315_ ) );
NOR2_X1 _17206_ ( .A1(_06039_ ), .A2(_01315_ ), .ZN(_01316_ ) );
INV_X1 _17207_ ( .A(_01273_ ), .ZN(_01317_ ) );
AND2_X1 _17208_ ( .A1(_01316_ ), .A2(_01317_ ), .ZN(_01318_ ) );
AND3_X1 _17209_ ( .A1(_00493_ ), .A2(_00495_ ), .A3(_01318_ ), .ZN(_01319_ ) );
NOR2_X1 _17210_ ( .A1(_00671_ ), .A2(_06038_ ), .ZN(_01320_ ) );
AOI21_X1 _17211_ ( .A(_01319_ ), .B1(_01320_ ), .B2(_01315_ ), .ZN(_01321_ ) );
BUF_X4 _17212_ ( .A(_01287_ ), .Z(_01322_ ) );
OAI21_X1 _17213_ ( .A(_01321_ ), .B1(_01286_ ), .B2(_01322_ ), .ZN(_01323_ ) );
MUX2_X1 _17214_ ( .A(\EX_LS_result_reg [14] ), .B(_01323_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
AND4_X1 _17215_ ( .A1(\io_master_arid [1] ), .A2(_00502_ ), .A3(_00504_ ), .A4(_01315_ ), .ZN(_01324_ ) );
AND3_X1 _17216_ ( .A1(_00496_ ), .A2(_00498_ ), .A3(_01316_ ), .ZN(_01325_ ) );
OAI21_X1 _17217_ ( .A(_01317_ ), .B1(_01324_ ), .B2(_01325_ ), .ZN(_01326_ ) );
OAI21_X1 _17218_ ( .A(_01326_ ), .B1(_01286_ ), .B2(_01322_ ), .ZN(_01327_ ) );
MUX2_X1 _17219_ ( .A(\EX_LS_result_reg [13] ), .B(_01327_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
NOR3_X1 _17220_ ( .A1(_00501_ ), .A2(_06040_ ), .A3(_01315_ ), .ZN(_01328_ ) );
NOR4_X1 _17221_ ( .A1(_00537_ ), .A2(_06039_ ), .A3(_01310_ ), .A4(_01314_ ), .ZN(_01329_ ) );
OAI21_X1 _17222_ ( .A(_01317_ ), .B1(_01328_ ), .B2(_01329_ ), .ZN(_01330_ ) );
OAI21_X1 _17223_ ( .A(_01330_ ), .B1(_01286_ ), .B2(_01322_ ), .ZN(_01331_ ) );
MUX2_X1 _17224_ ( .A(\EX_LS_result_reg [12] ), .B(_01331_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
OAI21_X1 _17225_ ( .A(_01291_ ), .B1(_01263_ ), .B2(_01320_ ), .ZN(_01332_ ) );
NAND2_X1 _17226_ ( .A1(_01332_ ), .A2(_01295_ ), .ZN(_01333_ ) );
MUX2_X1 _17227_ ( .A(\EX_LS_result_reg [30] ), .B(_01333_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _17228_ ( .A1(_00505_ ), .A2(_00507_ ), .A3(_01318_ ), .ZN(_01334_ ) );
NOR2_X2 _17229_ ( .A1(_00546_ ), .A2(_06037_ ), .ZN(_01335_ ) );
NAND2_X1 _17230_ ( .A1(_01335_ ), .A2(_01315_ ), .ZN(_01336_ ) );
OAI211_X1 _17231_ ( .A(_01334_ ), .B(_01336_ ), .C1(_01286_ ), .C2(_01322_ ), .ZN(_01337_ ) );
MUX2_X1 _17232_ ( .A(\EX_LS_result_reg [11] ), .B(_01337_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
NAND3_X1 _17233_ ( .A1(_00508_ ), .A2(_00510_ ), .A3(_01318_ ), .ZN(_01338_ ) );
NOR2_X2 _17234_ ( .A1(_00549_ ), .A2(_06038_ ), .ZN(_01339_ ) );
NAND2_X1 _17235_ ( .A1(_01339_ ), .A2(_01315_ ), .ZN(_01340_ ) );
OAI211_X1 _17236_ ( .A(_01338_ ), .B(_01340_ ), .C1(_01286_ ), .C2(_01322_ ), .ZN(_01341_ ) );
MUX2_X1 _17237_ ( .A(\EX_LS_result_reg [10] ), .B(_01341_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
NOR4_X1 _17238_ ( .A1(_00552_ ), .A2(_06039_ ), .A3(_01310_ ), .A4(_01314_ ), .ZN(_01342_ ) );
NOR3_X1 _17239_ ( .A1(_00513_ ), .A2(_06040_ ), .A3(_01315_ ), .ZN(_01343_ ) );
OAI21_X1 _17240_ ( .A(_01317_ ), .B1(_01342_ ), .B2(_01343_ ), .ZN(_01344_ ) );
OAI21_X1 _17241_ ( .A(_01344_ ), .B1(_01286_ ), .B2(_01322_ ), .ZN(_01345_ ) );
MUX2_X1 _17242_ ( .A(\EX_LS_result_reg [9] ), .B(_01345_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NOR2_X1 _17243_ ( .A1(_01089_ ), .A2(_06040_ ), .ZN(_01346_ ) );
NAND2_X1 _17244_ ( .A1(_01346_ ), .A2(_01315_ ), .ZN(_01347_ ) );
NAND3_X1 _17245_ ( .A1(_00514_ ), .A2(_00516_ ), .A3(_01318_ ), .ZN(_01348_ ) );
OAI211_X1 _17246_ ( .A(_01347_ ), .B(_01348_ ), .C1(_01286_ ), .C2(_01322_ ), .ZN(_01349_ ) );
MUX2_X1 _17247_ ( .A(\EX_LS_result_reg [8] ), .B(_01349_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
INV_X1 _17248_ ( .A(_01265_ ), .ZN(_01350_ ) );
NOR3_X1 _17249_ ( .A1(_00558_ ), .A2(_06039_ ), .A3(_01314_ ), .ZN(_01351_ ) );
INV_X1 _17250_ ( .A(_01351_ ), .ZN(_01352_ ) );
AOI21_X1 _17251_ ( .A(_01290_ ), .B1(_01352_ ), .B2(_01284_ ), .ZN(_01353_ ) );
AND4_X1 _17252_ ( .A1(\io_master_arid [1] ), .A2(_00517_ ), .A3(_00519_ ), .A4(_01290_ ), .ZN(_01354_ ) );
OAI21_X1 _17253_ ( .A(_01350_ ), .B1(_01353_ ), .B2(_01354_ ), .ZN(_01355_ ) );
OAI21_X1 _17254_ ( .A(_01266_ ), .B1(_01351_ ), .B2(_01283_ ), .ZN(_01356_ ) );
AOI21_X1 _17255_ ( .A(_01272_ ), .B1(_01355_ ), .B2(_01356_ ), .ZN(_01357_ ) );
NOR3_X1 _17256_ ( .A1(_01286_ ), .A2(\mylsu.typ_tmp [2] ), .A3(_01271_ ), .ZN(_01358_ ) );
OAI21_X1 _17257_ ( .A(_01322_ ), .B1(_01357_ ), .B2(_01358_ ), .ZN(_01359_ ) );
NAND2_X1 _17258_ ( .A1(_01359_ ), .A2(_01295_ ), .ZN(_01360_ ) );
MUX2_X1 _17259_ ( .A(\EX_LS_result_reg [7] ), .B(_01360_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
OR3_X1 _17260_ ( .A1(_00522_ ), .A2(_06039_ ), .A3(_01258_ ), .ZN(_01361_ ) );
AND4_X1 _17261_ ( .A1(_01975_ ), .A2(_00493_ ), .A3(_00495_ ), .A4(_01279_ ), .ZN(_01362_ ) );
AND3_X2 _17262_ ( .A1(_00559_ ), .A2(_00561_ ), .A3(_01975_ ), .ZN(_01363_ ) );
INV_X1 _17263_ ( .A(_01281_ ), .ZN(_01364_ ) );
MUX2_X1 _17264_ ( .A(_01363_ ), .B(_01320_ ), .S(_01364_ ), .Z(_01365_ ) );
INV_X1 _17265_ ( .A(_01279_ ), .ZN(_01366_ ) );
AOI21_X1 _17266_ ( .A(_01362_ ), .B1(_01365_ ), .B2(_01366_ ), .ZN(_01367_ ) );
OAI21_X1 _17267_ ( .A(_01361_ ), .B1(_01367_ ), .B2(_01314_ ), .ZN(_01368_ ) );
NOR2_X2 _17268_ ( .A1(_00522_ ), .A2(_06037_ ), .ZN(_01369_ ) );
MUX2_X2 _17269_ ( .A(_01363_ ), .B(_01369_ ), .S(_01256_ ), .Z(_01370_ ) );
MUX2_X2 _17270_ ( .A(_01369_ ), .B(_01370_ ), .S(_01275_ ), .Z(_01371_ ) );
MUX2_X1 _17271_ ( .A(_01370_ ), .B(_01371_ ), .S(_01350_ ), .Z(_01372_ ) );
MUX2_X1 _17272_ ( .A(_01372_ ), .B(_01368_ ), .S(_01272_ ), .Z(_01373_ ) );
MUX2_X1 _17273_ ( .A(_01368_ ), .B(_01373_ ), .S(_01322_ ), .Z(_01374_ ) );
MUX2_X1 _17274_ ( .A(\EX_LS_result_reg [6] ), .B(_01374_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _17275_ ( .A1(_06096_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01375_ ) );
NOR2_X1 _17276_ ( .A1(_01312_ ), .A2(_01314_ ), .ZN(_01376_ ) );
INV_X1 _17277_ ( .A(_01376_ ), .ZN(_01377_ ) );
NAND2_X1 _17278_ ( .A1(_00525_ ), .A2(_01377_ ), .ZN(_01378_ ) );
AND2_X1 _17279_ ( .A1(_01273_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01379_ ) );
NOR2_X1 _17280_ ( .A1(_01377_ ), .A2(_01379_ ), .ZN(_01380_ ) );
NAND3_X1 _17281_ ( .A1(_00464_ ), .A2(_00465_ ), .A3(_01380_ ), .ZN(_01381_ ) );
NAND4_X1 _17282_ ( .A1(_01378_ ), .A2(\mylsu.state [3] ), .A3(\io_master_arid [1] ), .A4(_01381_ ), .ZN(_01382_ ) );
NAND3_X1 _17283_ ( .A1(_00502_ ), .A2(\mylsu.araddr_tmp [1] ), .A3(_00504_ ), .ZN(_01383_ ) );
NAND3_X1 _17284_ ( .A1(_00496_ ), .A2(_06042_ ), .A3(_00498_ ), .ZN(_01384_ ) );
AND3_X1 _17285_ ( .A1(_01383_ ), .A2(_01384_ ), .A3(_01379_ ), .ZN(_01385_ ) );
OAI21_X1 _17286_ ( .A(_01375_ ), .B1(_01382_ ), .B2(_01385_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
OR3_X1 _17287_ ( .A1(_00528_ ), .A2(_06039_ ), .A3(_01258_ ), .ZN(_01386_ ) );
NOR3_X1 _17288_ ( .A1(_00501_ ), .A2(_06038_ ), .A3(_01366_ ), .ZN(_01387_ ) );
NOR2_X1 _17289_ ( .A1(_00537_ ), .A2(_06038_ ), .ZN(_01388_ ) );
MUX2_X1 _17290_ ( .A(_01388_ ), .B(_01292_ ), .S(_01281_ ), .Z(_01389_ ) );
AOI21_X1 _17291_ ( .A(_01387_ ), .B1(_01389_ ), .B2(_01366_ ), .ZN(_01390_ ) );
OAI21_X1 _17292_ ( .A(_01386_ ), .B1(_01390_ ), .B2(_01314_ ), .ZN(_01391_ ) );
NOR2_X2 _17293_ ( .A1(_00528_ ), .A2(_06037_ ), .ZN(_01392_ ) );
MUX2_X2 _17294_ ( .A(_01392_ ), .B(_01292_ ), .S(_01258_ ), .Z(_01393_ ) );
MUX2_X2 _17295_ ( .A(_01392_ ), .B(_01393_ ), .S(_01275_ ), .Z(_01394_ ) );
MUX2_X1 _17296_ ( .A(_01393_ ), .B(_01394_ ), .S(_01350_ ), .Z(_01395_ ) );
MUX2_X1 _17297_ ( .A(_01395_ ), .B(_01391_ ), .S(_01272_ ), .Z(_01396_ ) );
MUX2_X1 _17298_ ( .A(_01391_ ), .B(_01396_ ), .S(_01322_ ), .Z(_01397_ ) );
MUX2_X1 _17299_ ( .A(\EX_LS_result_reg [4] ), .B(_01397_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
OR3_X1 _17300_ ( .A1(_00531_ ), .A2(_06039_ ), .A3(_01258_ ), .ZN(_01398_ ) );
AND4_X1 _17301_ ( .A1(_01975_ ), .A2(_00505_ ), .A3(_00507_ ), .A4(_01279_ ), .ZN(_01399_ ) );
MUX2_X1 _17302_ ( .A(_01335_ ), .B(_01298_ ), .S(_01281_ ), .Z(_01400_ ) );
AOI21_X1 _17303_ ( .A(_01399_ ), .B1(_01400_ ), .B2(_01366_ ), .ZN(_01401_ ) );
OAI21_X1 _17304_ ( .A(_01398_ ), .B1(_01401_ ), .B2(_01314_ ), .ZN(_01402_ ) );
NOR2_X2 _17305_ ( .A1(_00531_ ), .A2(_06037_ ), .ZN(_01403_ ) );
MUX2_X2 _17306_ ( .A(_01403_ ), .B(_01298_ ), .S(_01258_ ), .Z(_01404_ ) );
MUX2_X2 _17307_ ( .A(_01403_ ), .B(_01404_ ), .S(_01275_ ), .Z(_01405_ ) );
MUX2_X1 _17308_ ( .A(_01404_ ), .B(_01405_ ), .S(_01350_ ), .Z(_01406_ ) );
MUX2_X1 _17309_ ( .A(_01406_ ), .B(_01402_ ), .S(_01272_ ), .Z(_01407_ ) );
MUX2_X1 _17310_ ( .A(_01402_ ), .B(_01407_ ), .S(_01287_ ), .Z(_01408_ ) );
MUX2_X1 _17311_ ( .A(\EX_LS_result_reg [3] ), .B(_01408_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
OR3_X1 _17312_ ( .A1(_00534_ ), .A2(_06039_ ), .A3(_01258_ ), .ZN(_01409_ ) );
AND4_X1 _17313_ ( .A1(_01975_ ), .A2(_00508_ ), .A3(_00510_ ), .A4(_01279_ ), .ZN(_01410_ ) );
MUX2_X1 _17314_ ( .A(_01339_ ), .B(_01301_ ), .S(_01281_ ), .Z(_01411_ ) );
AOI21_X1 _17315_ ( .A(_01410_ ), .B1(_01411_ ), .B2(_01366_ ), .ZN(_01412_ ) );
OAI21_X1 _17316_ ( .A(_01409_ ), .B1(_01412_ ), .B2(_01314_ ), .ZN(_01413_ ) );
NOR2_X1 _17317_ ( .A1(_00534_ ), .A2(_06037_ ), .ZN(_01414_ ) );
MUX2_X2 _17318_ ( .A(_01414_ ), .B(_01301_ ), .S(_01257_ ), .Z(_01415_ ) );
MUX2_X2 _17319_ ( .A(_01414_ ), .B(_01415_ ), .S(_01275_ ), .Z(_01416_ ) );
MUX2_X1 _17320_ ( .A(_01415_ ), .B(_01416_ ), .S(_01350_ ), .Z(_01417_ ) );
MUX2_X1 _17321_ ( .A(_01417_ ), .B(_01413_ ), .S(_01272_ ), .Z(_01418_ ) );
MUX2_X1 _17322_ ( .A(_01413_ ), .B(_01418_ ), .S(_01287_ ), .Z(_01419_ ) );
MUX2_X1 _17323_ ( .A(\EX_LS_result_reg [2] ), .B(_01419_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
AND4_X1 _17324_ ( .A1(\io_master_arid [1] ), .A2(_00502_ ), .A3(_00504_ ), .A4(_01310_ ), .ZN(_01420_ ) );
OAI21_X1 _17325_ ( .A(_01274_ ), .B1(_01266_ ), .B2(_01420_ ), .ZN(_01421_ ) );
NAND2_X1 _17326_ ( .A1(_01421_ ), .A2(_01295_ ), .ZN(_01422_ ) );
MUX2_X1 _17327_ ( .A(\EX_LS_result_reg [29] ), .B(_01422_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
OR3_X1 _17328_ ( .A1(_00540_ ), .A2(_06039_ ), .A3(_01258_ ), .ZN(_01423_ ) );
NOR3_X1 _17329_ ( .A1(_00513_ ), .A2(_06038_ ), .A3(_01366_ ), .ZN(_01424_ ) );
NOR2_X2 _17330_ ( .A1(_00552_ ), .A2(_06038_ ), .ZN(_01425_ ) );
MUX2_X2 _17331_ ( .A(_01304_ ), .B(_01425_ ), .S(_01364_ ), .Z(_01426_ ) );
AOI21_X1 _17332_ ( .A(_01424_ ), .B1(_01426_ ), .B2(_01366_ ), .ZN(_01427_ ) );
OAI21_X2 _17333_ ( .A(_01423_ ), .B1(_01427_ ), .B2(_01314_ ), .ZN(_01428_ ) );
NOR2_X2 _17334_ ( .A1(_00540_ ), .A2(_06037_ ), .ZN(_01429_ ) );
MUX2_X2 _17335_ ( .A(_01429_ ), .B(_01304_ ), .S(_01257_ ), .Z(_01430_ ) );
MUX2_X2 _17336_ ( .A(_01429_ ), .B(_01430_ ), .S(_01275_ ), .Z(_01431_ ) );
MUX2_X1 _17337_ ( .A(_01430_ ), .B(_01431_ ), .S(_01350_ ), .Z(_01432_ ) );
MUX2_X1 _17338_ ( .A(_01432_ ), .B(_01428_ ), .S(_01272_ ), .Z(_01433_ ) );
MUX2_X1 _17339_ ( .A(_01428_ ), .B(_01433_ ), .S(_01287_ ), .Z(_01434_ ) );
MUX2_X1 _17340_ ( .A(\EX_LS_result_reg [1] ), .B(_01434_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
AOI211_X1 _17341_ ( .A(_06095_ ), .B(_06040_ ), .C1(_00769_ ), .C2(_01380_ ), .ZN(_01435_ ) );
NAND2_X1 _17342_ ( .A1(_00543_ ), .A2(_01377_ ), .ZN(_01436_ ) );
NAND2_X1 _17343_ ( .A1(_01435_ ), .A2(_01436_ ), .ZN(_01437_ ) );
MUX2_X1 _17344_ ( .A(_01089_ ), .B(_00605_ ), .S(_06042_ ), .Z(_01438_ ) );
AOI21_X1 _17345_ ( .A(_01437_ ), .B1(_01379_ ), .B2(_01438_ ), .ZN(_01439_ ) );
AND2_X1 _17346_ ( .A1(_06096_ ), .A2(\EX_LS_result_reg [0] ), .ZN(_01440_ ) );
OR2_X1 _17347_ ( .A1(_01439_ ), .A2(_01440_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
NOR3_X1 _17348_ ( .A1(_00537_ ), .A2(_06040_ ), .A3(_01275_ ), .ZN(_01441_ ) );
OAI21_X1 _17349_ ( .A(_01274_ ), .B1(_01266_ ), .B2(_01441_ ), .ZN(_01442_ ) );
NAND2_X1 _17350_ ( .A1(_01442_ ), .A2(_01295_ ), .ZN(_01443_ ) );
MUX2_X1 _17351_ ( .A(\EX_LS_result_reg [28] ), .B(_01443_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
OAI21_X1 _17352_ ( .A(_01291_ ), .B1(_01263_ ), .B2(_01335_ ), .ZN(_01444_ ) );
AOI22_X1 _17353_ ( .A1(_01444_ ), .A2(_01289_ ), .B1(_06096_ ), .B2(_04197_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
NOR3_X1 _17354_ ( .A1(_00549_ ), .A2(_06040_ ), .A3(_01263_ ), .ZN(_01445_ ) );
OAI21_X1 _17355_ ( .A(_01274_ ), .B1(_01266_ ), .B2(_01445_ ), .ZN(_01446_ ) );
AOI22_X1 _17356_ ( .A1(_01446_ ), .A2(_01289_ ), .B1(_06096_ ), .B2(_04222_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
OAI21_X1 _17357_ ( .A(_01291_ ), .B1(_01263_ ), .B2(_01425_ ), .ZN(_01447_ ) );
AOI22_X1 _17358_ ( .A1(_01447_ ), .A2(_01289_ ), .B1(_06096_ ), .B2(_04246_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
OAI21_X1 _17359_ ( .A(_01291_ ), .B1(_01263_ ), .B2(_01346_ ), .ZN(_01448_ ) );
NAND2_X1 _17360_ ( .A1(_01448_ ), .A2(_01295_ ), .ZN(_01449_ ) );
MUX2_X1 _17361_ ( .A(\EX_LS_result_reg [24] ), .B(_01449_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
OAI21_X1 _17362_ ( .A(_01291_ ), .B1(_01263_ ), .B2(_01280_ ), .ZN(_01450_ ) );
NAND2_X1 _17363_ ( .A1(_01450_ ), .A2(_01295_ ), .ZN(_01451_ ) );
MUX2_X1 _17364_ ( .A(\EX_LS_result_reg [23] ), .B(_01451_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _17365_ ( .A1(_01274_ ), .A2(_01290_ ), .A3(_01363_ ), .ZN(_01452_ ) );
OR3_X1 _17366_ ( .A1(_01261_ ), .A2(_01350_ ), .A3(_01273_ ), .ZN(_01453_ ) );
NAND3_X1 _17367_ ( .A1(_01452_ ), .A2(_01294_ ), .A3(_01453_ ), .ZN(_01454_ ) );
MUX2_X1 _17368_ ( .A(\EX_LS_result_reg [22] ), .B(_01454_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17369_ ( .A1(_00457_ ), .A2(\io_master_arid [1] ), .A3(_01310_ ), .ZN(_01455_ ) );
OAI21_X1 _17370_ ( .A(_01274_ ), .B1(_01266_ ), .B2(_01455_ ), .ZN(_01456_ ) );
NAND2_X1 _17371_ ( .A1(_01456_ ), .A2(_01295_ ), .ZN(_01457_ ) );
MUX2_X1 _17372_ ( .A(\EX_LS_result_reg [31] ), .B(_01457_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
INV_X1 _17373_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01458_ ) );
NOR2_X1 _17374_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(\LS_WB_waddr_reg [2] ), .ZN(_01459_ ) );
INV_X1 _17375_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01460_ ) );
INV_X1 _17376_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01461_ ) );
NAND3_X1 _17377_ ( .A1(_01459_ ), .A2(_01460_ ), .A3(_01461_ ), .ZN(_01462_ ) );
AND2_X1 _17378_ ( .A1(_01535_ ), .A2(LS_WB_wen_reg ), .ZN(_01463_ ) );
NAND2_X1 _17379_ ( .A1(_01462_ ), .A2(_01463_ ), .ZN(_01464_ ) );
BUF_X4 _17380_ ( .A(_01464_ ), .Z(_01465_ ) );
NOR2_X1 _17381_ ( .A1(_01465_ ), .A2(_01461_ ), .ZN(_01466_ ) );
INV_X1 _17382_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01467_ ) );
NOR2_X1 _17383_ ( .A1(_01465_ ), .A2(_01467_ ), .ZN(_01468_ ) );
AND4_X1 _17384_ ( .A1(_01458_ ), .A2(_01466_ ), .A3(_01468_ ), .A4(_01460_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _17385_ ( .A1(_01464_ ), .A2(_01460_ ), .ZN(_01469_ ) );
AND4_X1 _17386_ ( .A1(_01458_ ), .A2(_01469_ ), .A3(_01468_ ), .A4(_01461_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
AOI21_X1 _17387_ ( .A(_01465_ ), .B1(_01460_ ), .B2(_01461_ ), .ZN(_01470_ ) );
NOR4_X1 _17388_ ( .A1(_01470_ ), .A2(_01458_ ), .A3(_01467_ ), .A4(_01465_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
CLKBUF_X1 _17389_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
AOI21_X1 _17390_ ( .A(_01465_ ), .B1(_01458_ ), .B2(_01467_ ), .ZN(_01471_ ) );
NOR4_X1 _17391_ ( .A1(_01471_ ), .A2(_01469_ ), .A3(_01461_ ), .A4(_01465_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
NOR4_X1 _17392_ ( .A1(_01471_ ), .A2(_01466_ ), .A3(_01460_ ), .A4(_01465_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17393_ ( .A1(_01471_ ), .A2(_01460_ ), .A3(_01461_ ), .A4(_01465_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17394_ ( .A1(_01458_ ), .A2(_01469_ ), .A3(_01468_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
NOR4_X1 _17395_ ( .A1(_01470_ ), .A2(_01468_ ), .A3(_01458_ ), .A4(_01465_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR2_X1 _17396_ ( .A1(_01464_ ), .A2(_01458_ ), .ZN(_01472_ ) );
AND4_X1 _17397_ ( .A1(_01467_ ), .A2(_01466_ ), .A3(_01472_ ), .A4(_01460_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17398_ ( .A1(_01467_ ), .A2(_01469_ ), .A3(_01472_ ), .A4(_01461_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17399_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01466_ ), .A3(_01472_ ), .A4(_01460_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17400_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01469_ ), .A3(_01472_ ), .A4(_01461_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17401_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(_01469_ ), .A3(_01468_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17402_ ( .A1(_01467_ ), .A2(_01469_ ), .A3(_01472_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17403_ ( .A1(_01470_ ), .A2(_01472_ ), .A3(_01467_ ), .A4(_01465_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17404_ ( .A1(_01938_ ), .A2(_01570_ ), .A3(_01945_ ), .ZN(_01473_ ) );
NAND2_X1 _17405_ ( .A1(_01473_ ), .A2(_01570_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17406_ ( .A(reset ), .B(_01938_ ), .C1(_01939_ ), .C2(_01959_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17407_ ( .A(_01462_ ), .Z(_01474_ ) );
CLKBUF_X2 _17408_ ( .A(_01463_ ), .Z(_01475_ ) );
AND3_X1 _17409_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17410_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17411_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17412_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17413_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17414_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17415_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17416_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17417_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17418_ ( .A1(_01474_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01475_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17419_ ( .A(_01462_ ), .Z(_01476_ ) );
CLKBUF_X2 _17420_ ( .A(_01463_ ), .Z(_01477_ ) );
AND3_X1 _17421_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17422_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17423_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17424_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17425_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17426_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17427_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17428_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17429_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17430_ ( .A1(_01476_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01477_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17431_ ( .A(_01462_ ), .Z(_01478_ ) );
CLKBUF_X2 _17432_ ( .A(_01463_ ), .Z(_01479_ ) );
AND3_X1 _17433_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17434_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17435_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17436_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17437_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17438_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17439_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17440_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17441_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17442_ ( .A1(_01478_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01479_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17443_ ( .A1(_01462_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01463_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17444_ ( .A1(_01462_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01463_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_D ) );
AND3_X1 _17445_ ( .A1(_01624_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17446_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01480_ ) );
AND2_X1 _17447_ ( .A1(_01480_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01481_ ) );
INV_X1 _17448_ ( .A(_01481_ ), .ZN(_01482_ ) );
NOR2_X1 _17449_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01483_ ) );
OAI211_X1 _17450_ ( .A(_01535_ ), .B(\mysc.state [0] ), .C1(_01482_ ), .C2(_01483_ ), .ZN(_01484_ ) );
INV_X1 _17451_ ( .A(_01484_ ), .ZN(_01485_ ) );
OR3_X1 _17452_ ( .A1(_01485_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17453_ ( .A1(_01482_ ), .A2(reset ), .A3(_01483_ ), .ZN(_01486_ ) );
NAND2_X1 _17454_ ( .A1(_01486_ ), .A2(\mysc.state [0] ), .ZN(_01487_ ) );
OR3_X1 _17455_ ( .A1(_03882_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01488_ ) );
NAND2_X1 _17456_ ( .A1(_01487_ ), .A2(_01488_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17457_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07961_ ) );
CLKGATE_X1 _17458_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07962_ ) );
CLKGATE_X1 _17459_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07963_ ) );
CLKGATE_X1 _17460_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07964_ ) );
CLKGATE_X1 _17461_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07965_ ) );
CLKGATE_X1 _17462_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_07966_ ) );
CLKGATE_X1 _17463_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_07967_ ) );
CLKGATE_X1 _17464_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_07968_ ) );
CLKGATE_X1 _17465_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_07969_ ) );
CLKGATE_X1 _17466_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_07970_ ) );
CLKGATE_X1 _17467_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_07971_ ) );
CLKGATE_X1 _17468_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07972_ ) );
CLKGATE_X1 _17469_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07973_ ) );
CLKGATE_X1 _17470_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_07974_ ) );
CLKGATE_X1 _17471_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_07975_ ) );
CLKGATE_X1 _17472_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07976_ ) );
CLKGATE_X1 _17473_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07977_ ) );
CLKGATE_X1 _17474_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_07978_ ) );
CLKGATE_X1 _17475_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_07979_ ) );
CLKGATE_X1 _17476_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ), .GCK(_07980_ ) );
CLKGATE_X1 _17477_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .GCK(_07981_ ) );
CLKGATE_X1 _17478_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_07982_ ) );
CLKGATE_X1 _17479_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_07983_ ) );
CLKGATE_X1 _17480_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_07984_ ) );
CLKGATE_X1 _17481_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_07985_ ) );
CLKGATE_X1 _17482_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_07986_ ) );
CLKGATE_X1 _17483_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_07987_ ) );
CLKGATE_X1 _17484_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_07988_ ) );
CLKGATE_X1 _17485_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_07989_ ) );
CLKGATE_X1 _17486_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_07990_ ) );
CLKGATE_X1 _17487_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_07991_ ) );
CLKGATE_X1 _17488_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_07992_ ) );
CLKGATE_X1 _17489_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_07993_ ) );
CLKGATE_X1 _17490_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_07994_ ) );
CLKGATE_X1 _17491_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_07995_ ) );
CLKGATE_X1 _17492_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07996_ ) );
CLKGATE_X1 _17493_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07997_ ) );
CLKGATE_X1 _17494_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07998_ ) );
CLKGATE_X1 _17495_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07999_ ) );
CLKGATE_X1 _17496_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08000_ ) );
CLKGATE_X1 _17497_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08001_ ) );
CLKGATE_X1 _17498_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08002_ ) );
CLKGATE_X1 _17499_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08003_ ) );
CLKGATE_X1 _17500_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08004_ ) );
CLKGATE_X1 _17501_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08005_ ) );
CLKGATE_X1 _17502_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08006_ ) );
CLKGATE_X1 _17503_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08007_ ) );
CLKGATE_X1 _17504_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08008_ ) );
CLKGATE_X1 _17505_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08009_ ) );
CLKGATE_X1 _17506_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08010_ ) );
CLKGATE_X1 _17507_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08011_ ) );
CLKGATE_X1 _17508_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_08012_ ) );
CLKGATE_X1 _17509_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08013_ ) );
CLKGATE_X1 _17510_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08014_ ) );
CLKGATE_X1 _17511_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08015_ ) );
CLKGATE_X1 _17512_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08016_ ) );
CLKGATE_X1 _17513_ ( .CK(clock ), .E(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08017_ ) );
CLKGATE_X1 _17514_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_08018_ ) );
CLKGATE_X1 _17515_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ), .GCK(_08019_ ) );
CLKGATE_X1 _17516_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08020_ ) );
CLKGATE_X1 _17517_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08021_ ) );
CLKGATE_X1 _17518_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08022_ ) );
CLKGATE_X1 _17519_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08023_ ) );
CLKGATE_X1 _17520_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08024_ ) );
CLKGATE_X1 _17521_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08025_ ) );
LOGIC1_X1 _17522_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17523_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08255_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08256_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08257_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08258_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08259_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08260_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08261_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08262_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08263_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08264_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08265_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08266_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08267_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08268_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08269_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08270_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08271_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08272_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08273_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08274_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08275_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08276_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08277_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08278_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08279_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08280_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08281_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08282_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08283_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08284_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08285_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08025_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08286_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08024_ ), .Q(\mtvec [31] ), .QN(_08287_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08024_ ), .Q(\mtvec [30] ), .QN(_08288_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08024_ ), .Q(\mtvec [21] ), .QN(_08289_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08024_ ), .Q(\mtvec [20] ), .QN(_08290_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08024_ ), .Q(\mtvec [19] ), .QN(_08291_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08024_ ), .Q(\mtvec [18] ), .QN(_08292_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08024_ ), .Q(\mtvec [17] ), .QN(_08293_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08024_ ), .Q(\mtvec [16] ), .QN(_08294_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08024_ ), .Q(\mtvec [15] ), .QN(_08295_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08024_ ), .Q(\mtvec [14] ), .QN(_08296_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08024_ ), .Q(\mtvec [13] ), .QN(_08297_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08024_ ), .Q(\mtvec [12] ), .QN(_08298_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08024_ ), .Q(\mtvec [29] ), .QN(_08299_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08024_ ), .Q(\mtvec [11] ), .QN(_08300_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08024_ ), .Q(\mtvec [10] ), .QN(_08301_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08024_ ), .Q(\mtvec [9] ), .QN(_08302_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08024_ ), .Q(\mtvec [8] ), .QN(_08303_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08024_ ), .Q(\mtvec [7] ), .QN(_08304_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08024_ ), .Q(\mtvec [6] ), .QN(_08305_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08024_ ), .Q(\mtvec [5] ), .QN(_08306_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08024_ ), .Q(\mtvec [4] ), .QN(_08307_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08024_ ), .Q(\mtvec [3] ), .QN(_08308_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08024_ ), .Q(\mtvec [2] ), .QN(_08309_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08024_ ), .Q(\mtvec [28] ), .QN(_08310_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08024_ ), .Q(\mtvec [1] ), .QN(_08311_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08024_ ), .Q(\mtvec [0] ), .QN(_08312_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08024_ ), .Q(\mtvec [27] ), .QN(_08313_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08024_ ), .Q(\mtvec [26] ), .QN(_08314_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08024_ ), .Q(\mtvec [25] ), .QN(_08315_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08024_ ), .Q(\mtvec [24] ), .QN(_08316_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08024_ ), .Q(\mtvec [23] ), .QN(_08317_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08024_ ), .Q(\mtvec [22] ), .QN(_08318_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08023_ ), .Q(\mepc [31] ), .QN(_08319_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08023_ ), .Q(\mepc [30] ), .QN(_08320_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08023_ ), .Q(\mepc [21] ), .QN(_08321_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08023_ ), .Q(\mepc [20] ), .QN(_08322_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08023_ ), .Q(\mepc [19] ), .QN(_08323_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08023_ ), .Q(\mepc [18] ), .QN(_08324_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08023_ ), .Q(\mepc [17] ), .QN(_08325_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08023_ ), .Q(\mepc [16] ), .QN(_08326_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08023_ ), .Q(\mepc [15] ), .QN(_08327_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08023_ ), .Q(\mepc [14] ), .QN(_08328_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08023_ ), .Q(\mepc [13] ), .QN(_08329_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08023_ ), .Q(\mepc [12] ), .QN(_08330_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08023_ ), .Q(\mepc [29] ), .QN(_08331_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08023_ ), .Q(\mepc [11] ), .QN(_08332_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08023_ ), .Q(\mepc [10] ), .QN(_08333_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08023_ ), .Q(\mepc [9] ), .QN(_08334_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08023_ ), .Q(\mepc [8] ), .QN(_08335_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08023_ ), .Q(\mepc [7] ), .QN(_08336_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08023_ ), .Q(\mepc [6] ), .QN(_08337_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08023_ ), .Q(\mepc [5] ), .QN(_08338_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08023_ ), .Q(\mepc [4] ), .QN(_08339_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08023_ ), .Q(\mepc [3] ), .QN(_08340_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08023_ ), .Q(\mepc [2] ), .QN(_08341_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08023_ ), .Q(\mepc [28] ), .QN(_08342_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08023_ ), .Q(\mepc [1] ), .QN(_08343_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08023_ ), .Q(\mepc [0] ), .QN(_08344_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08023_ ), .Q(\mepc [27] ), .QN(_08345_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08023_ ), .Q(\mepc [26] ), .QN(_08346_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08023_ ), .Q(\mepc [25] ), .QN(_08347_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08023_ ), .Q(\mepc [24] ), .QN(_08348_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08023_ ), .Q(\mepc [23] ), .QN(_08349_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08023_ ), .Q(\mepc [22] ), .QN(_08350_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08351_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08352_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08353_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08254_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08253_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08252_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08251_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08250_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08249_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08248_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08247_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08246_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08245_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08244_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08243_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08242_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08241_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08240_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08239_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08238_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08237_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08236_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08235_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08234_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08233_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00086_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08232_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00087_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08231_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00088_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08230_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00089_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08229_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00090_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08228_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00091_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08227_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00092_ ), .CK(_08022_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08354_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PP0__Q ( .D(_00093_ ), .CK(clock ), .Q(excp_written ), .QN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08226_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08355_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08356_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08357_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08358_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08359_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08360_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08361_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08362_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08363_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08364_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08365_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08366_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08367_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08368_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08369_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08370_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08371_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08372_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08373_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08374_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08375_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08376_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08377_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08378_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08379_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08380_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08381_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08382_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08383_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08384_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08021_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08225_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00094_ ), .CK(_08020_ ), .Q(\myec.state [1] ), .QN(_08224_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00095_ ), .CK(_08020_ ), .Q(\myec.state [0] ), .QN(_08385_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PN0__Q ( .D(_00096_ ), .CK(clock ), .Q(check_quest ), .QN(_08386_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08223_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08387_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08388_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08389_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08390_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08391_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08392_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08393_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08394_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08395_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08396_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08222_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00097_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08221_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00098_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08220_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00099_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08219_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00100_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08218_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00101_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08217_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00102_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08216_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00103_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08215_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00104_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08214_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00105_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08213_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00106_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08212_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00107_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08211_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00108_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08210_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00109_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08209_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00110_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08208_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00111_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08207_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00112_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08206_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00113_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08205_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00114_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08204_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00115_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08203_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00116_ ), .CK(_08019_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08202_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q ( .D(_00117_ ), .CK(_08018_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08201_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_1 ( .D(_00118_ ), .CK(_08018_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08200_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_2 ( .D(_00119_ ), .CK(_08018_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08199_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_3 ( .D(_00120_ ), .CK(_08018_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08198_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_4 ( .D(_00121_ ), .CK(_08018_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08197_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q ( .D(_00122_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [30] ), .QN(_08196_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_1 ( .D(_00123_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [29] ), .QN(_08195_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_10 ( .D(_00124_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [20] ), .QN(_08194_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_11 ( .D(_00125_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [19] ), .QN(_08193_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_12 ( .D(_00126_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [18] ), .QN(_08192_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_13 ( .D(_00127_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [17] ), .QN(_08191_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_14 ( .D(_00128_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [16] ), .QN(_08190_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_15 ( .D(_00129_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [15] ), .QN(_08189_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_16 ( .D(_00130_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [14] ), .QN(_08188_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_17 ( .D(_00131_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [13] ), .QN(_08187_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_18 ( .D(_00132_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [12] ), .QN(_08186_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_19 ( .D(_00133_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [11] ), .QN(_08185_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_2 ( .D(_00134_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [28] ), .QN(_08184_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_20 ( .D(_00135_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [10] ), .QN(_08183_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_21 ( .D(_00136_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [9] ), .QN(_08182_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_22 ( .D(_00137_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [8] ), .QN(_08181_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_23 ( .D(_00138_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [7] ), .QN(_08180_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_24 ( .D(_00139_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [6] ), .QN(_08179_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_25 ( .D(_00140_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [5] ), .QN(_08178_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_26 ( .D(_00141_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [4] ), .QN(_08177_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_27 ( .D(_00142_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [3] ), .QN(_08176_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_28 ( .D(_00143_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [2] ), .QN(_08175_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_29 ( .D(_00144_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [1] ), .QN(_08174_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_3 ( .D(_00145_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [27] ), .QN(_08173_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_30 ( .D(_00146_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [0] ), .QN(_08172_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_4 ( .D(_00147_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [26] ), .QN(_08171_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_5 ( .D(_00148_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [25] ), .QN(_08170_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_6 ( .D(_00149_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [24] ), .QN(_08169_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_7 ( .D(_00150_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [23] ), .QN(_08168_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_8 ( .D(_00151_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [22] ), .QN(_08167_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_9 ( .D(_00152_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [21] ), .QN(_08166_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN1P__Q ( .D(_00153_ ), .CK(_08017_ ), .Q(\myexu.pc_jump [31] ), .QN(_08165_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q ( .D(_00154_ ), .CK(_08018_ ), .Q(\EX_LS_pc [31] ), .QN(_08164_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_1 ( .D(_00155_ ), .CK(_08018_ ), .Q(\EX_LS_pc [30] ), .QN(_08163_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_10 ( .D(_00156_ ), .CK(_08018_ ), .Q(\EX_LS_pc [21] ), .QN(_08162_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_11 ( .D(_00157_ ), .CK(_08018_ ), .Q(\EX_LS_pc [20] ), .QN(_08161_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_12 ( .D(_00158_ ), .CK(_08018_ ), .Q(\EX_LS_pc [19] ), .QN(_08160_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_13 ( .D(_00159_ ), .CK(_08018_ ), .Q(\EX_LS_pc [18] ), .QN(_08159_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_14 ( .D(_00160_ ), .CK(_08018_ ), .Q(\EX_LS_pc [17] ), .QN(_08158_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_15 ( .D(_00161_ ), .CK(_08018_ ), .Q(\EX_LS_pc [16] ), .QN(_08157_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_16 ( .D(_00162_ ), .CK(_08018_ ), .Q(\EX_LS_pc [15] ), .QN(_08156_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_17 ( .D(_00163_ ), .CK(_08018_ ), .Q(\EX_LS_pc [14] ), .QN(_08155_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_18 ( .D(_00164_ ), .CK(_08018_ ), .Q(\EX_LS_pc [13] ), .QN(_08154_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_19 ( .D(_00165_ ), .CK(_08018_ ), .Q(\EX_LS_pc [12] ), .QN(_08153_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_2 ( .D(_00166_ ), .CK(_08018_ ), .Q(\EX_LS_pc [29] ), .QN(_08152_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_20 ( .D(_00167_ ), .CK(_08018_ ), .Q(\EX_LS_pc [11] ), .QN(_08151_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_21 ( .D(_00168_ ), .CK(_08018_ ), .Q(\EX_LS_pc [10] ), .QN(_08150_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_22 ( .D(_00169_ ), .CK(_08018_ ), .Q(\EX_LS_pc [9] ), .QN(_08149_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_23 ( .D(_00170_ ), .CK(_08018_ ), .Q(\EX_LS_pc [8] ), .QN(_08148_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_24 ( .D(_00171_ ), .CK(_08018_ ), .Q(\EX_LS_pc [7] ), .QN(_08147_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_25 ( .D(_00172_ ), .CK(_08018_ ), .Q(\EX_LS_pc [6] ), .QN(_08146_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_26 ( .D(_00173_ ), .CK(_08018_ ), .Q(\EX_LS_pc [5] ), .QN(_08145_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_27 ( .D(_00174_ ), .CK(_08018_ ), .Q(\EX_LS_pc [4] ), .QN(_08144_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_28 ( .D(_00175_ ), .CK(_08018_ ), .Q(\EX_LS_pc [3] ), .QN(_08143_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_29 ( .D(_00176_ ), .CK(_08018_ ), .Q(\EX_LS_pc [2] ), .QN(_08142_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_3 ( .D(_00177_ ), .CK(_08018_ ), .Q(\EX_LS_pc [28] ), .QN(_08141_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_30 ( .D(_00178_ ), .CK(_08018_ ), .Q(\EX_LS_pc [1] ), .QN(_08140_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_31 ( .D(_00179_ ), .CK(_08018_ ), .Q(\EX_LS_pc [0] ), .QN(_08139_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_4 ( .D(_00180_ ), .CK(_08018_ ), .Q(\EX_LS_pc [27] ), .QN(_08138_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_5 ( .D(_00181_ ), .CK(_08018_ ), .Q(\EX_LS_pc [26] ), .QN(_08137_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_6 ( .D(_00182_ ), .CK(_08018_ ), .Q(\EX_LS_pc [25] ), .QN(_08136_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_7 ( .D(_00183_ ), .CK(_08018_ ), .Q(\EX_LS_pc [24] ), .QN(_08135_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_8 ( .D(_00184_ ), .CK(_08018_ ), .Q(\EX_LS_pc [23] ), .QN(_08134_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_9 ( .D(_00185_ ), .CK(_08018_ ), .Q(\EX_LS_pc [22] ), .QN(_08397_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08398_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08399_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08400_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08401_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08402_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08403_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08404_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08405_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08406_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08407_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08408_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08409_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08410_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08411_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08412_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08413_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08414_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08415_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08416_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08417_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08418_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08419_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08420_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08421_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08422_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08423_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08424_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08425_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08426_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08427_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08428_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08019_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08429_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08019_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PN0__Q ( .D(_00187_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q ( .D(_00186_ ), .CK(_08018_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_1 ( .D(_00188_ ), .CK(_08018_ ), .Q(\EX_LS_flag [1] ), .QN(_08133_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_2 ( .D(_00189_ ), .CK(_08018_ ), .Q(\EX_LS_flag [0] ), .QN(_08132_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_3 ( .D(_00190_ ), .CK(_08018_ ), .Q(\EX_LS_typ [4] ), .QN(_08131_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_4 ( .D(_00191_ ), .CK(_08018_ ), .Q(\EX_LS_typ [3] ), .QN(_08130_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_5 ( .D(_00192_ ), .CK(_08018_ ), .Q(\EX_LS_typ [2] ), .QN(_08129_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_6 ( .D(_00193_ ), .CK(_08018_ ), .Q(\EX_LS_typ [1] ), .QN(_08128_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_7 ( .D(_00194_ ), .CK(_08018_ ), .Q(\EX_LS_typ [0] ), .QN(_08127_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00195_ ), .CK(_08016_ ), .Q(\ID_EX_csr [11] ), .QN(_08126_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00196_ ), .CK(_08016_ ), .Q(\ID_EX_csr [10] ), .QN(_08125_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00197_ ), .CK(_08016_ ), .Q(\ID_EX_csr [1] ), .QN(_08124_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00198_ ), .CK(_08016_ ), .Q(\ID_EX_csr [0] ), .QN(_08123_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00199_ ), .CK(_08016_ ), .Q(\ID_EX_csr [9] ), .QN(_08122_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00200_ ), .CK(_08016_ ), .Q(\ID_EX_csr [8] ), .QN(_08121_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00201_ ), .CK(_08016_ ), .Q(\ID_EX_csr [7] ), .QN(_08120_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00202_ ), .CK(_08016_ ), .Q(\ID_EX_csr [6] ), .QN(_08119_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00203_ ), .CK(_08016_ ), .Q(\ID_EX_csr [5] ), .QN(_08118_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00204_ ), .CK(_08016_ ), .Q(\ID_EX_csr [4] ), .QN(_08117_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00205_ ), .CK(_08016_ ), .Q(\ID_EX_csr [3] ), .QN(_08116_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00206_ ), .CK(_08016_ ), .Q(\ID_EX_csr [2] ), .QN(_08115_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00207_ ), .CK(_08015_ ), .Q(exception_quest_IDU ), .QN(_08114_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00208_ ), .CK(_08014_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08013_ ), .Q(\ID_EX_imm [31] ), .QN(_08430_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08013_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08013_ ), .Q(\ID_EX_imm [21] ), .QN(_08431_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08013_ ), .Q(\ID_EX_imm [20] ), .QN(_08432_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08013_ ), .Q(\ID_EX_imm [19] ), .QN(_08433_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08013_ ), .Q(\ID_EX_imm [18] ), .QN(_08434_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08013_ ), .Q(\ID_EX_imm [17] ), .QN(_08435_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08013_ ), .Q(\ID_EX_imm [16] ), .QN(_08436_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08013_ ), .Q(\ID_EX_imm [15] ), .QN(_08437_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08013_ ), .Q(\ID_EX_imm [14] ), .QN(_08438_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08013_ ), .Q(\ID_EX_imm [13] ), .QN(_08439_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08013_ ), .Q(\ID_EX_imm [12] ), .QN(_08440_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08013_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08013_ ), .Q(\ID_EX_imm [11] ), .QN(_08441_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08013_ ), .Q(\ID_EX_imm [10] ), .QN(_08442_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08013_ ), .Q(\ID_EX_imm [9] ), .QN(_08443_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08013_ ), .Q(\ID_EX_imm [8] ), .QN(_08444_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08013_ ), .Q(\ID_EX_imm [7] ), .QN(_08445_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08013_ ), .Q(\ID_EX_imm [6] ), .QN(_08446_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08013_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08013_ ), .Q(\ID_EX_imm [4] ), .QN(_08447_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08013_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08013_ ), .Q(\ID_EX_imm [2] ), .QN(_08448_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08013_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08013_ ), .Q(\ID_EX_imm [1] ), .QN(_08449_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08013_ ), .Q(\ID_EX_imm [0] ), .QN(_08450_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08013_ ), .Q(\ID_EX_imm [27] ), .QN(_08451_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08013_ ), .Q(\ID_EX_imm [26] ), .QN(_08452_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08013_ ), .Q(\ID_EX_imm [25] ), .QN(_08453_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08013_ ), .Q(\ID_EX_imm [24] ), .QN(_08454_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08013_ ), .Q(\ID_EX_imm [23] ), .QN(_08455_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08013_ ), .Q(\ID_EX_imm [22] ), .QN(_08456_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08012_ ), .Q(\ID_EX_pc [31] ), .QN(_08457_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08012_ ), .Q(\ID_EX_pc [30] ), .QN(_08458_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08012_ ), .Q(\ID_EX_pc [21] ), .QN(_08459_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08012_ ), .Q(\ID_EX_pc [20] ), .QN(_08460_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08012_ ), .Q(\ID_EX_pc [19] ), .QN(_08461_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08012_ ), .Q(\ID_EX_pc [18] ), .QN(_08462_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08012_ ), .Q(\ID_EX_pc [17] ), .QN(_08463_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08012_ ), .Q(\ID_EX_pc [16] ), .QN(_08464_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08012_ ), .Q(\ID_EX_pc [15] ), .QN(_08465_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08012_ ), .Q(\ID_EX_pc [14] ), .QN(_08466_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08012_ ), .Q(\ID_EX_pc [13] ), .QN(_08467_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08012_ ), .Q(\ID_EX_pc [12] ), .QN(_08468_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08012_ ), .Q(\ID_EX_pc [29] ), .QN(_08469_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08012_ ), .Q(\ID_EX_pc [11] ), .QN(_08470_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08012_ ), .Q(\ID_EX_pc [10] ), .QN(_08471_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08012_ ), .Q(\ID_EX_pc [9] ), .QN(_08472_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08012_ ), .Q(\ID_EX_pc [8] ), .QN(_08473_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08012_ ), .Q(\ID_EX_pc [7] ), .QN(_08474_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08012_ ), .Q(\ID_EX_pc [6] ), .QN(_08475_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08012_ ), .Q(\ID_EX_pc [5] ), .QN(_08476_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08012_ ), .Q(\ID_EX_pc [4] ), .QN(_08477_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08012_ ), .Q(\ID_EX_pc [3] ), .QN(_08478_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08012_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08012_ ), .Q(\ID_EX_pc [28] ), .QN(_08479_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08012_ ), .Q(\ID_EX_pc [1] ), .QN(_08480_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08012_ ), .Q(\ID_EX_pc [0] ), .QN(_08481_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08012_ ), .Q(\ID_EX_pc [27] ), .QN(_08482_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08012_ ), .Q(\ID_EX_pc [26] ), .QN(_08483_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08012_ ), .Q(\ID_EX_pc [25] ), .QN(_08484_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08012_ ), .Q(\ID_EX_pc [24] ), .QN(_08485_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08012_ ), .Q(\ID_EX_pc [23] ), .QN(_08486_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08012_ ), .Q(\ID_EX_pc [22] ), .QN(_08113_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00209_ ), .CK(_08011_ ), .Q(\ID_EX_rd [4] ), .QN(_08112_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00210_ ), .CK(_08011_ ), .Q(\ID_EX_rd [3] ), .QN(_08111_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00211_ ), .CK(_08011_ ), .Q(\ID_EX_rd [2] ), .QN(_08110_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00212_ ), .CK(_08011_ ), .Q(\ID_EX_rd [1] ), .QN(_08109_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00213_ ), .CK(_08011_ ), .Q(\ID_EX_rd [0] ), .QN(_08108_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00214_ ), .CK(_08010_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08107_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00215_ ), .CK(_08010_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08106_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00217_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08104_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00216_ ), .CK(_08010_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08105_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00219_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08102_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00218_ ), .CK(_08010_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08103_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00221_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08100_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00220_ ), .CK(_08010_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08101_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00223_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08098_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00222_ ), .CK(_08009_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08099_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00224_ ), .CK(_08009_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08097_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00226_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08095_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00225_ ), .CK(_08009_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08096_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00228_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08093_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00227_ ), .CK(_08009_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08094_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00230_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08091_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00229_ ), .CK(_08009_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08092_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00232_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08089_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_08008_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08090_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00233_ ), .CK(_08007_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08088_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08488_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00234_ ), .CK(_08006_ ), .Q(\ID_EX_typ [7] ), .QN(_08487_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00235_ ), .CK(_08006_ ), .Q(\ID_EX_typ [6] ), .QN(_08087_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00236_ ), .CK(_08006_ ), .Q(\ID_EX_typ [5] ), .QN(_08086_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00237_ ), .CK(_08006_ ), .Q(\ID_EX_typ [4] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00238_ ), .CK(_08006_ ), .Q(\ID_EX_typ [3] ), .QN(_08085_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00239_ ), .CK(_08006_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00240_ ), .CK(_08006_ ), .Q(\ID_EX_typ [1] ), .QN(_08084_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00241_ ), .CK(_08006_ ), .Q(\ID_EX_typ [0] ), .QN(_08489_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08005_ ), .Q(check_assert ), .QN(_08490_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08004_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08004_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08004_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08004_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08004_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08004_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08004_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08004_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08004_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08004_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08004_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08004_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08004_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08004_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08004_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08004_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08004_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08004_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08004_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08004_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08004_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08004_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08004_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08004_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08004_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08004_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08004_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08004_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08004_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08004_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08004_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08004_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08491_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08492_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08493_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08494_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08495_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08496_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08497_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08498_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08499_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08500_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08501_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08502_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08503_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08504_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08505_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08506_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08507_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08508_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08509_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08510_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08511_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08512_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08513_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08514_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08515_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08516_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08517_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08518_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08519_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08520_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08521_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08003_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08522_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08523_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08524_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08525_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08526_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08527_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08528_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08529_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08530_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08531_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08532_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08533_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08534_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08535_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08536_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08537_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08538_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08539_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08540_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08541_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08542_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08543_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08544_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08545_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08546_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08547_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08548_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08549_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08550_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08551_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08552_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08553_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08002_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08554_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08555_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08556_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08557_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08558_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08559_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08560_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08561_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08562_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08563_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08564_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08565_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08566_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08567_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08001_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08000_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07999_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07998_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07997_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07996_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07995_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07994_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07993_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07992_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08083_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00242_ ), .CK(_07991_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08082_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00243_ ), .CK(_07990_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08081_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00244_ ), .CK(_07989_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_07988_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08080_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_07987_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_07986_ ), .Q(\IF_ID_pc [30] ), .QN(_08079_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00247_ ), .CK(_07986_ ), .Q(\IF_ID_pc [21] ), .QN(_08078_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00248_ ), .CK(_07986_ ), .Q(\IF_ID_pc [20] ), .QN(_08077_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00249_ ), .CK(_07986_ ), .Q(\IF_ID_pc [19] ), .QN(_08076_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00250_ ), .CK(_07986_ ), .Q(\IF_ID_pc [18] ), .QN(_08075_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00251_ ), .CK(_07986_ ), .Q(\IF_ID_pc [17] ), .QN(_08074_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00252_ ), .CK(_07986_ ), .Q(\IF_ID_pc [16] ), .QN(_08073_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00253_ ), .CK(_07986_ ), .Q(\IF_ID_pc [15] ), .QN(_08072_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00254_ ), .CK(_07986_ ), .Q(\IF_ID_pc [14] ), .QN(_08071_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00255_ ), .CK(_07986_ ), .Q(\IF_ID_pc [13] ), .QN(_08070_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00256_ ), .CK(_07986_ ), .Q(\IF_ID_pc [12] ), .QN(_08069_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00257_ ), .CK(_07986_ ), .Q(\IF_ID_pc [29] ), .QN(_08068_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00258_ ), .CK(_07986_ ), .Q(\IF_ID_pc [11] ), .QN(_08067_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00259_ ), .CK(_07986_ ), .Q(\IF_ID_pc [10] ), .QN(_08066_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00260_ ), .CK(_07986_ ), .Q(\IF_ID_pc [9] ), .QN(_08065_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00261_ ), .CK(_07986_ ), .Q(\IF_ID_pc [8] ), .QN(_08064_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00262_ ), .CK(_07986_ ), .Q(\IF_ID_pc [7] ), .QN(_08063_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00263_ ), .CK(_07986_ ), .Q(\IF_ID_pc [6] ), .QN(_08062_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00264_ ), .CK(_07986_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00265_ ), .CK(_07986_ ), .Q(\IF_ID_pc [4] ), .QN(_08061_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00267_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08060_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00266_ ), .CK(_07986_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00269_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08058_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00268_ ), .CK(_07986_ ), .Q(\IF_ID_pc [2] ), .QN(_08059_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00270_ ), .CK(_07986_ ), .Q(\IF_ID_pc [28] ), .QN(_08057_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00271_ ), .CK(_07986_ ), .Q(\IF_ID_pc [1] ), .QN(_08056_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00272_ ), .CK(_07986_ ), .Q(\IF_ID_pc [27] ), .QN(_08055_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00273_ ), .CK(_07986_ ), .Q(\IF_ID_pc [26] ), .QN(_08054_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00274_ ), .CK(_07986_ ), .Q(\IF_ID_pc [25] ), .QN(_08053_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00275_ ), .CK(_07986_ ), .Q(\IF_ID_pc [24] ), .QN(_08052_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00276_ ), .CK(_07986_ ), .Q(\IF_ID_pc [23] ), .QN(_08051_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00277_ ), .CK(_07986_ ), .Q(\IF_ID_pc [22] ), .QN(_08050_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00278_ ), .CK(_07986_ ), .Q(\IF_ID_pc [31] ), .QN(_08049_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08856_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08048_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00279_ ), .CK(_07985_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08855_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00281_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00280_ ), .CK(_07984_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08047_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08857_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08858_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08859_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08860_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08861_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08862_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08863_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08864_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08865_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08866_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08867_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08868_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08869_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08870_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08871_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08872_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08873_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08874_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08875_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08876_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08877_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08878_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08879_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08880_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08881_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08882_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08883_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08884_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08885_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08886_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08887_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07983_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08888_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08889_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08890_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08891_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08892_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08893_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08894_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08895_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08896_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08897_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08898_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08899_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08900_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08901_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08902_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08903_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08904_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08905_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08906_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08907_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08908_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08909_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08910_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08911_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08912_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08913_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08914_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08915_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08916_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08917_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08918_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08919_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07982_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08046_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PN0P__Q ( .D(_00282_ ), .CK(_07981_ ), .Q(LS_WB_pc ), .QN(_08045_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PN0P__Q ( .D(_00283_ ), .CK(_07980_ ), .Q(\mylsu.previous_load_done ), .QN(_08920_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08921_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08922_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08923_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_07983_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_07983_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08924_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_07983_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08044_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00284_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08043_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00285_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08042_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00286_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08041_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00287_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08040_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00288_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08039_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00289_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08038_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00290_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08037_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00291_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08036_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00292_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08035_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00293_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08034_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00294_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08033_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00295_ ), .CK(_07983_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08925_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_07983_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08926_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_07983_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08927_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_07983_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08928_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_07983_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08929_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08930_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08931_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08932_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08933_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08934_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08935_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08936_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08937_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08938_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08939_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08940_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08941_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08942_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08943_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08944_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08945_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08946_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08947_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08948_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08949_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08950_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08951_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08952_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08953_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08954_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08955_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08956_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08957_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08958_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08959_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08960_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_07983_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08961_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08962_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_08963_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_08964_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_08965_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_08966_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_08967_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_08968_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_08969_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_08970_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_08971_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_08972_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_08973_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_08974_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_08975_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_08976_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_08977_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_08978_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_08979_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_08980_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_08981_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_08982_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_08983_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_08984_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_08985_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_08986_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_08987_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_08988_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_08989_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_08990_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_08991_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_08992_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_07979_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08032_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q ( .D(_00296_ ), .CK(_07978_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_B ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_1 ( .D(_00297_ ), .CK(_07978_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08031_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_2 ( .D(_00298_ ), .CK(_07978_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08030_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_3 ( .D(_00299_ ), .CK(_07978_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08029_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_4 ( .D(_00300_ ), .CK(_07978_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08028_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_5 ( .D(_00301_ ), .CK(_07978_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08027_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PN0P__Q ( .D(_00302_ ), .CK(_07978_ ), .Q(LS_WB_wen_reg ), .QN(_08993_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_08994_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_08995_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07977_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07976_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07975_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07974_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07973_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07972_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07971_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07970_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07969_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07968_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07967_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07966_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07965_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07964_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07963_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07962_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00303_ ), .CK(_07961_ ), .Q(loaduse_clear ), .QN(_08996_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_08997_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_08998_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08026_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(fanout_net_22 ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(fanout_net_22 ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(fanout_net_22 ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(fanout_net_22 ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(fanout_net_22 ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(fanout_net_35 ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(fanout_net_35 ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(fanout_net_35 ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(fanout_net_35 ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(fanout_net_35 ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_40 ) );

endmodule
