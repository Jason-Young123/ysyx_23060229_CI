//Generate the verilog at 2025-09-29T16:31:17 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire _09036_ ;
wire _09037_ ;
wire _09038_ ;
wire _09039_ ;
wire _09040_ ;
wire _09041_ ;
wire _09042_ ;
wire _09043_ ;
wire _09044_ ;
wire _09045_ ;
wire _09046_ ;
wire _09047_ ;
wire _09048_ ;
wire _09049_ ;
wire _09050_ ;
wire _09051_ ;
wire _09052_ ;
wire _09053_ ;
wire _09054_ ;
wire _09055_ ;
wire _09056_ ;
wire _09057_ ;
wire _09058_ ;
wire _09059_ ;
wire _09060_ ;
wire _09061_ ;
wire _09062_ ;
wire _09063_ ;
wire _09064_ ;
wire _09065_ ;
wire _09066_ ;
wire _09067_ ;
wire _09068_ ;
wire _09069_ ;
wire _09070_ ;
wire _09071_ ;
wire _09072_ ;
wire _09073_ ;
wire _09074_ ;
wire _09075_ ;
wire _09076_ ;
wire _09077_ ;
wire _09078_ ;
wire _09079_ ;
wire _09080_ ;
wire _09081_ ;
wire _09082_ ;
wire _09083_ ;
wire _09084_ ;
wire _09085_ ;
wire _09086_ ;
wire _09087_ ;
wire _09088_ ;
wire _09089_ ;
wire _09090_ ;
wire _09091_ ;
wire _09092_ ;
wire _09093_ ;
wire _09094_ ;
wire _09095_ ;
wire _09096_ ;
wire _09097_ ;
wire _09098_ ;
wire _09099_ ;
wire _09100_ ;
wire _09101_ ;
wire _09102_ ;
wire _09103_ ;
wire _09104_ ;
wire _09105_ ;
wire _09106_ ;
wire _09107_ ;
wire _09108_ ;
wire _09109_ ;
wire _09110_ ;
wire _09111_ ;
wire _09112_ ;
wire _09113_ ;
wire _09114_ ;
wire _09115_ ;
wire _09116_ ;
wire _09117_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[4]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[5]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[6]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data[7]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.tag[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_D ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

INV_X1 _09118_ ( .A(\LS_WB_wdata_csreg [31] ), .ZN(_01663_ ) );
NOR2_X1 _09119_ ( .A1(_01663_ ), .A2(fanout_net_1 ), .ZN(_00000_ ) );
INV_X2 _09120_ ( .A(fanout_net_1 ), .ZN(_01664_ ) );
BUF_X4 _09121_ ( .A(_01664_ ), .Z(_01665_ ) );
AND3_X4 _09122_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01666_ ) );
AND3_X4 _09123_ ( .A1(_01666_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01667_ ) );
AND3_X4 _09124_ ( .A1(_01667_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01668_ ) );
AND3_X4 _09125_ ( .A1(_01668_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01669_ ) );
AND3_X4 _09126_ ( .A1(_01669_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01670_ ) );
AND3_X4 _09127_ ( .A1(_01670_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01671_ ) );
AND3_X4 _09128_ ( .A1(_01671_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01672_ ) );
AND3_X4 _09129_ ( .A1(_01672_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01673_ ) );
AND3_X4 _09130_ ( .A1(_01673_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01674_ ) );
AND3_X4 _09131_ ( .A1(_01674_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01675_ ) );
AND3_X4 _09132_ ( .A1(_01675_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01676_ ) );
AND3_X4 _09133_ ( .A1(_01676_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01677_ ) );
AND3_X4 _09134_ ( .A1(_01677_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01678_ ) );
AND2_X4 _09135_ ( .A1(_01678_ ), .A2(\myclint.mtime [27] ), .ZN(_01679_ ) );
AND2_X1 _09136_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01680_ ) );
AND2_X1 _09137_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01681_ ) );
AND4_X4 _09138_ ( .A1(\myclint.mtime [33] ), .A2(_01679_ ), .A3(_01680_ ), .A4(_01681_ ), .ZN(_01682_ ) );
AND3_X4 _09139_ ( .A1(_01682_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01683_ ) );
AND3_X4 _09140_ ( .A1(_01683_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [35] ), .ZN(_01684_ ) );
AND3_X4 _09141_ ( .A1(_01684_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [37] ), .ZN(_01685_ ) );
AND2_X4 _09142_ ( .A1(_01685_ ), .A2(\myclint.mtime [39] ), .ZN(_01686_ ) );
AND2_X1 _09143_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01687_ ) );
AND2_X4 _09144_ ( .A1(_01686_ ), .A2(_01687_ ), .ZN(_01688_ ) );
AND2_X2 _09145_ ( .A1(\myclint.mtime [42] ), .A2(\myclint.mtime [43] ), .ZN(_01689_ ) );
AND2_X4 _09146_ ( .A1(_01688_ ), .A2(_01689_ ), .ZN(_01690_ ) );
AND2_X1 _09147_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01691_ ) );
AND3_X1 _09148_ ( .A1(_01691_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01692_ ) );
NAND2_X4 _09149_ ( .A1(_01690_ ), .A2(_01692_ ), .ZN(_01693_ ) );
AND2_X1 _09150_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01694_ ) );
INV_X1 _09151_ ( .A(_01694_ ), .ZN(_01695_ ) );
NOR2_X4 _09152_ ( .A1(_01693_ ), .A2(_01695_ ), .ZN(_01696_ ) );
AND2_X1 _09153_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01697_ ) );
AND2_X4 _09154_ ( .A1(_01696_ ), .A2(_01697_ ), .ZN(_01698_ ) );
AND2_X1 _09155_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01699_ ) );
AND2_X4 _09156_ ( .A1(_01698_ ), .A2(_01699_ ), .ZN(_01700_ ) );
AND2_X1 _09157_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01701_ ) );
AND2_X4 _09158_ ( .A1(_01700_ ), .A2(_01701_ ), .ZN(_01702_ ) );
AND2_X1 _09159_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01703_ ) );
AND2_X4 _09160_ ( .A1(_01702_ ), .A2(_01703_ ), .ZN(_01704_ ) );
AND2_X1 _09161_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01705_ ) );
AND2_X4 _09162_ ( .A1(_01704_ ), .A2(_01705_ ), .ZN(_01706_ ) );
NAND3_X4 _09163_ ( .A1(_01706_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01707_ ) );
NOR2_X2 _09164_ ( .A1(_01707_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01708_ ) );
OAI21_X1 _09165_ ( .A(_01665_ ), .B1(_01708_ ), .B2(\myclint.mtime [63] ), .ZN(_01709_ ) );
AND2_X2 _09166_ ( .A1(_01679_ ), .A2(_01681_ ), .ZN(_01710_ ) );
AND2_X1 _09167_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01711_ ) );
AND3_X2 _09168_ ( .A1(_01710_ ), .A2(_01711_ ), .A3(_01680_ ), .ZN(_01712_ ) );
AND3_X4 _09169_ ( .A1(_01712_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01713_ ) );
NAND2_X4 _09170_ ( .A1(_01713_ ), .A2(\myclint.mtime [36] ), .ZN(_01714_ ) );
INV_X1 _09171_ ( .A(\myclint.mtime [38] ), .ZN(_01715_ ) );
INV_X1 _09172_ ( .A(\myclint.mtime [37] ), .ZN(_01716_ ) );
NOR3_X2 _09173_ ( .A1(_01714_ ), .A2(_01715_ ), .A3(_01716_ ), .ZN(_01717_ ) );
AND2_X2 _09174_ ( .A1(_01717_ ), .A2(\myclint.mtime [39] ), .ZN(_01718_ ) );
AND2_X2 _09175_ ( .A1(_01718_ ), .A2(_01687_ ), .ZN(_01719_ ) );
AND2_X2 _09176_ ( .A1(_01719_ ), .A2(_01689_ ), .ZN(_01720_ ) );
AND2_X2 _09177_ ( .A1(_01720_ ), .A2(_01692_ ), .ZN(_01721_ ) );
AND2_X2 _09178_ ( .A1(_01721_ ), .A2(_01694_ ), .ZN(_01722_ ) );
AND2_X2 _09179_ ( .A1(_01722_ ), .A2(_01697_ ), .ZN(_01723_ ) );
AND2_X2 _09180_ ( .A1(_01723_ ), .A2(_01699_ ), .ZN(_01724_ ) );
AND2_X2 _09181_ ( .A1(_01724_ ), .A2(_01701_ ), .ZN(_01725_ ) );
AND2_X2 _09182_ ( .A1(_01725_ ), .A2(_01703_ ), .ZN(_01726_ ) );
AND2_X2 _09183_ ( .A1(_01726_ ), .A2(_01705_ ), .ZN(_01727_ ) );
NAND3_X1 _09184_ ( .A1(_01727_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01728_ ) );
NOR2_X1 _09185_ ( .A1(_01728_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01729_ ) );
AOI21_X1 _09186_ ( .A(_01709_ ), .B1(\myclint.mtime [63] ), .B2(_01729_ ), .ZN(_00001_ ) );
AND2_X1 _09187_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_01730_ ) );
AND3_X1 _09188_ ( .A1(_01730_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01731_ ) );
AND4_X1 _09189_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01732_ ) );
AND2_X1 _09190_ ( .A1(_01731_ ), .A2(_01732_ ), .ZN(_01733_ ) );
AND2_X1 _09191_ ( .A1(\myclint.mtime [24] ), .A2(\myclint.mtime [25] ), .ZN(_01734_ ) );
AND3_X1 _09192_ ( .A1(_01734_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [27] ), .ZN(_01735_ ) );
NAND4_X1 _09193_ ( .A1(_01733_ ), .A2(_01680_ ), .A3(_01681_ ), .A4(_01735_ ), .ZN(_01736_ ) );
AND2_X1 _09194_ ( .A1(_01666_ ), .A2(\myclint.mtime [3] ), .ZN(_01737_ ) );
AND4_X1 _09195_ ( .A1(\myclint.mtime [6] ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [5] ), .A4(\myclint.mtime [7] ), .ZN(_01738_ ) );
AND2_X1 _09196_ ( .A1(_01737_ ), .A2(_01738_ ), .ZN(_01739_ ) );
AND4_X1 _09197_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01740_ ) );
AND2_X1 _09198_ ( .A1(\myclint.mtime [10] ), .A2(\myclint.mtime [11] ), .ZN(_01741_ ) );
AND4_X1 _09199_ ( .A1(\myclint.mtime [8] ), .A2(_01740_ ), .A3(\myclint.mtime [9] ), .A4(_01741_ ), .ZN(_01742_ ) );
NAND2_X1 _09200_ ( .A1(_01739_ ), .A2(_01742_ ), .ZN(_01743_ ) );
NOR2_X1 _09201_ ( .A1(_01736_ ), .A2(_01743_ ), .ZN(_01744_ ) );
AND3_X1 _09202_ ( .A1(_01711_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01745_ ) );
AND2_X1 _09203_ ( .A1(_01689_ ), .A2(_01687_ ), .ZN(_01746_ ) );
AND4_X1 _09204_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01747_ ) );
AND4_X1 _09205_ ( .A1(_01692_ ), .A2(_01745_ ), .A3(_01746_ ), .A4(_01747_ ), .ZN(_01748_ ) );
AND2_X1 _09206_ ( .A1(_01744_ ), .A2(_01748_ ), .ZN(_01749_ ) );
AND4_X1 _09207_ ( .A1(_01701_ ), .A2(_01699_ ), .A3(_01697_ ), .A4(_01694_ ), .ZN(_01750_ ) );
AND2_X1 _09208_ ( .A1(_01749_ ), .A2(_01750_ ), .ZN(_01751_ ) );
AND4_X1 _09209_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01752_ ) );
AND2_X1 _09210_ ( .A1(_01751_ ), .A2(_01752_ ), .ZN(_01753_ ) );
AND3_X1 _09211_ ( .A1(_01753_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01754_ ) );
XNOR2_X1 _09212_ ( .A(_01754_ ), .B(\myclint.mtime [62] ), .ZN(_01755_ ) );
NOR2_X1 _09213_ ( .A1(_01755_ ), .A2(fanout_net_1 ), .ZN(_00002_ ) );
INV_X1 _09214_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01756_ ) );
AND4_X1 _09215_ ( .A1(_01756_ ), .A2(_01722_ ), .A3(\myclint.mtime [53] ), .A4(_01697_ ), .ZN(_01757_ ) );
BUF_X4 _09216_ ( .A(_01664_ ), .Z(_01758_ ) );
AND3_X1 _09217_ ( .A1(_01696_ ), .A2(_01756_ ), .A3(_01697_ ), .ZN(_01759_ ) );
OAI21_X1 _09218_ ( .A(_01758_ ), .B1(_01759_ ), .B2(\myclint.mtime [53] ), .ZN(_01760_ ) );
NOR2_X1 _09219_ ( .A1(_01757_ ), .A2(_01760_ ), .ZN(_00003_ ) );
AND2_X1 _09220_ ( .A1(_01697_ ), .A2(_01694_ ), .ZN(_01761_ ) );
AND2_X1 _09221_ ( .A1(_01749_ ), .A2(_01761_ ), .ZN(_01762_ ) );
XNOR2_X1 _09222_ ( .A(_01762_ ), .B(\myclint.mtime [52] ), .ZN(_01763_ ) );
NOR2_X1 _09223_ ( .A1(_01763_ ), .A2(fanout_net_1 ), .ZN(_00004_ ) );
NOR3_X1 _09224_ ( .A1(_01693_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01695_ ), .ZN(_01764_ ) );
OAI21_X1 _09225_ ( .A(_01665_ ), .B1(_01764_ ), .B2(\myclint.mtime [51] ), .ZN(_01765_ ) );
INV_X1 _09226_ ( .A(_01721_ ), .ZN(_01766_ ) );
NOR3_X1 _09227_ ( .A1(_01766_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01695_ ), .ZN(_01767_ ) );
AOI21_X1 _09228_ ( .A(_01765_ ), .B1(_01767_ ), .B2(\myclint.mtime [51] ), .ZN(_00005_ ) );
INV_X1 _09229_ ( .A(_01744_ ), .ZN(_01768_ ) );
INV_X1 _09230_ ( .A(_01748_ ), .ZN(_01769_ ) );
OR4_X1 _09231_ ( .A1(\myclint.mtime [50] ), .A2(_01768_ ), .A3(_01695_ ), .A4(_01769_ ), .ZN(_01770_ ) );
AND3_X1 _09232_ ( .A1(_01744_ ), .A2(_01694_ ), .A3(_01748_ ), .ZN(_01771_ ) );
INV_X1 _09233_ ( .A(_01771_ ), .ZN(_01772_ ) );
NAND2_X1 _09234_ ( .A1(_01772_ ), .A2(\myclint.mtime [50] ), .ZN(_01773_ ) );
AOI21_X1 _09235_ ( .A(fanout_net_1 ), .B1(_01770_ ), .B2(_01773_ ), .ZN(_00006_ ) );
INV_X1 _09236_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01774_ ) );
AND4_X1 _09237_ ( .A1(\myclint.mtime [49] ), .A2(_01720_ ), .A3(_01774_ ), .A4(_01692_ ), .ZN(_01775_ ) );
AND3_X1 _09238_ ( .A1(_01690_ ), .A2(_01774_ ), .A3(_01692_ ), .ZN(_01776_ ) );
OAI21_X1 _09239_ ( .A(_01758_ ), .B1(_01776_ ), .B2(\myclint.mtime [49] ), .ZN(_01777_ ) );
NOR2_X1 _09240_ ( .A1(_01775_ ), .A2(_01777_ ), .ZN(_00007_ ) );
OAI21_X1 _09241_ ( .A(\myclint.mtime [48] ), .B1(_01768_ ), .B2(_01769_ ), .ZN(_01778_ ) );
OR4_X1 _09242_ ( .A1(\myclint.mtime [48] ), .A2(_01736_ ), .A3(_01769_ ), .A4(_01743_ ), .ZN(_01779_ ) );
AOI21_X1 _09243_ ( .A(fanout_net_1 ), .B1(_01778_ ), .B2(_01779_ ), .ZN(_00008_ ) );
NAND3_X1 _09244_ ( .A1(_01688_ ), .A2(_01691_ ), .A3(_01689_ ), .ZN(_01780_ ) );
NOR2_X1 _09245_ ( .A1(_01780_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01781_ ) );
OAI21_X1 _09246_ ( .A(_01665_ ), .B1(_01781_ ), .B2(\myclint.mtime [47] ), .ZN(_01782_ ) );
NAND3_X1 _09247_ ( .A1(_01719_ ), .A2(\myclint.mtime [44] ), .A3(_01689_ ), .ZN(_01783_ ) );
INV_X1 _09248_ ( .A(\myclint.mtime [45] ), .ZN(_01784_ ) );
NOR3_X1 _09249_ ( .A1(_01783_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01784_ ), .ZN(_01785_ ) );
AOI21_X1 _09250_ ( .A(_01782_ ), .B1(_01785_ ), .B2(\myclint.mtime [47] ), .ZN(_00009_ ) );
AND2_X1 _09251_ ( .A1(_01745_ ), .A2(_01747_ ), .ZN(_01786_ ) );
AND2_X1 _09252_ ( .A1(_01744_ ), .A2(_01786_ ), .ZN(_01787_ ) );
AND3_X1 _09253_ ( .A1(_01787_ ), .A2(_01691_ ), .A3(_01746_ ), .ZN(_01788_ ) );
XNOR2_X1 _09254_ ( .A(_01788_ ), .B(\myclint.mtime [46] ), .ZN(_01789_ ) );
NOR2_X1 _09255_ ( .A1(_01789_ ), .A2(fanout_net_1 ), .ZN(_00010_ ) );
INV_X1 _09256_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01790_ ) );
NAND3_X1 _09257_ ( .A1(_01688_ ), .A2(_01790_ ), .A3(_01689_ ), .ZN(_01791_ ) );
AOI21_X1 _09258_ ( .A(fanout_net_1 ), .B1(_01791_ ), .B2(_01784_ ), .ZN(_01792_ ) );
NAND4_X1 _09259_ ( .A1(_01719_ ), .A2(\myclint.mtime [45] ), .A3(_01790_ ), .A4(_01689_ ), .ZN(_01793_ ) );
AND2_X1 _09260_ ( .A1(_01792_ ), .A2(_01793_ ), .ZN(_00011_ ) );
AND2_X1 _09261_ ( .A1(_01787_ ), .A2(_01746_ ), .ZN(_01794_ ) );
XNOR2_X1 _09262_ ( .A(_01794_ ), .B(\myclint.mtime [44] ), .ZN(_01795_ ) );
NOR2_X1 _09263_ ( .A1(_01795_ ), .A2(fanout_net_1 ), .ZN(_00012_ ) );
INV_X1 _09264_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01796_ ) );
AND4_X1 _09265_ ( .A1(\myclint.mtime [61] ), .A2(_01726_ ), .A3(_01796_ ), .A4(_01705_ ), .ZN(_01797_ ) );
AND3_X1 _09266_ ( .A1(_01704_ ), .A2(_01796_ ), .A3(_01705_ ), .ZN(_01798_ ) );
OAI21_X1 _09267_ ( .A(_01758_ ), .B1(_01798_ ), .B2(\myclint.mtime [61] ), .ZN(_01799_ ) );
NOR2_X1 _09268_ ( .A1(_01797_ ), .A2(_01799_ ), .ZN(_00013_ ) );
NAND3_X1 _09269_ ( .A1(_01744_ ), .A2(_01687_ ), .A3(_01786_ ), .ZN(_01800_ ) );
OR3_X1 _09270_ ( .A1(_01800_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [43] ), .ZN(_01801_ ) );
OAI21_X1 _09271_ ( .A(\myclint.mtime [43] ), .B1(_01800_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01802_ ) );
AOI21_X1 _09272_ ( .A(fanout_net_1 ), .B1(_01801_ ), .B2(_01802_ ), .ZN(_00014_ ) );
OR2_X1 _09273_ ( .A1(_01800_ ), .A2(\myclint.mtime [42] ), .ZN(_01803_ ) );
NAND2_X1 _09274_ ( .A1(_01800_ ), .A2(\myclint.mtime [42] ), .ZN(_01804_ ) );
AOI21_X1 _09275_ ( .A(fanout_net_1 ), .B1(_01803_ ), .B2(_01804_ ), .ZN(_00015_ ) );
INV_X1 _09276_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01805_ ) );
AND4_X1 _09277_ ( .A1(\myclint.mtime [41] ), .A2(_01717_ ), .A3(_01805_ ), .A4(\myclint.mtime [39] ), .ZN(_01806_ ) );
AND3_X1 _09278_ ( .A1(_01685_ ), .A2(_01805_ ), .A3(\myclint.mtime [39] ), .ZN(_01807_ ) );
OAI21_X1 _09279_ ( .A(_01758_ ), .B1(_01807_ ), .B2(\myclint.mtime [41] ), .ZN(_01808_ ) );
NOR2_X1 _09280_ ( .A1(_01806_ ), .A2(_01808_ ), .ZN(_00016_ ) );
XNOR2_X1 _09281_ ( .A(_01787_ ), .B(\myclint.mtime [40] ), .ZN(_01809_ ) );
NOR2_X1 _09282_ ( .A1(_01809_ ), .A2(fanout_net_1 ), .ZN(_00017_ ) );
NOR3_X1 _09283_ ( .A1(_01714_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01716_ ), .ZN(_01810_ ) );
AND2_X1 _09284_ ( .A1(_01810_ ), .A2(\myclint.mtime [39] ), .ZN(_01811_ ) );
OAI21_X1 _09285_ ( .A(_01758_ ), .B1(_01810_ ), .B2(\myclint.mtime [39] ), .ZN(_01812_ ) );
NOR2_X1 _09286_ ( .A1(_01811_ ), .A2(_01812_ ), .ZN(_00018_ ) );
BUF_X2 _09287_ ( .A(_01664_ ), .Z(_01813_ ) );
NAND4_X1 _09288_ ( .A1(_01679_ ), .A2(\myclint.mtime [33] ), .A3(_01680_ ), .A4(_01681_ ), .ZN(_01814_ ) );
INV_X1 _09289_ ( .A(\myclint.mtime [32] ), .ZN(_01815_ ) );
NOR2_X1 _09290_ ( .A1(_01814_ ), .A2(_01815_ ), .ZN(_01816_ ) );
AND3_X1 _09291_ ( .A1(_01816_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01817_ ) );
AND3_X1 _09292_ ( .A1(_01817_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .ZN(_01818_ ) );
OAI21_X1 _09293_ ( .A(_01813_ ), .B1(_01818_ ), .B2(\myclint.mtime [38] ), .ZN(_01819_ ) );
NOR2_X1 _09294_ ( .A1(_01819_ ), .A2(_01685_ ), .ZN(_00019_ ) );
INV_X1 _09295_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01820_ ) );
NAND3_X1 _09296_ ( .A1(_01683_ ), .A2(_01820_ ), .A3(\myclint.mtime [35] ), .ZN(_01821_ ) );
AOI21_X1 _09297_ ( .A(fanout_net_1 ), .B1(_01821_ ), .B2(_01716_ ), .ZN(_01822_ ) );
AND2_X1 _09298_ ( .A1(_01712_ ), .A2(\myclint.mtime [34] ), .ZN(_01823_ ) );
NAND4_X1 _09299_ ( .A1(_01823_ ), .A2(\myclint.mtime [37] ), .A3(_01820_ ), .A4(\myclint.mtime [35] ), .ZN(_01824_ ) );
AND2_X1 _09300_ ( .A1(_01822_ ), .A2(_01824_ ), .ZN(_00020_ ) );
OAI21_X1 _09301_ ( .A(_01813_ ), .B1(_01817_ ), .B2(\myclint.mtime [36] ), .ZN(_01825_ ) );
NOR2_X1 _09302_ ( .A1(_01825_ ), .A2(_01684_ ), .ZN(_00021_ ) );
INV_X1 _09303_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01826_ ) );
AND3_X1 _09304_ ( .A1(_01712_ ), .A2(_01826_ ), .A3(\myclint.mtime [35] ), .ZN(_01827_ ) );
NOR3_X1 _09305_ ( .A1(_01814_ ), .A2(_01815_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01828_ ) );
OAI21_X1 _09306_ ( .A(_01758_ ), .B1(_01828_ ), .B2(\myclint.mtime [35] ), .ZN(_01829_ ) );
NOR2_X1 _09307_ ( .A1(_01827_ ), .A2(_01829_ ), .ZN(_00022_ ) );
OAI21_X1 _09308_ ( .A(_01813_ ), .B1(_01816_ ), .B2(\myclint.mtime [34] ), .ZN(_01830_ ) );
NOR2_X1 _09309_ ( .A1(_01830_ ), .A2(_01683_ ), .ZN(_00023_ ) );
XNOR2_X1 _09310_ ( .A(_01753_ ), .B(\myclint.mtime [60] ), .ZN(_01831_ ) );
NOR2_X1 _09311_ ( .A1(_01831_ ), .A2(fanout_net_1 ), .ZN(_00024_ ) );
INV_X1 _09312_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01832_ ) );
AND3_X1 _09313_ ( .A1(_01710_ ), .A2(_01832_ ), .A3(_01680_ ), .ZN(_01833_ ) );
AND2_X1 _09314_ ( .A1(_01833_ ), .A2(\myclint.mtime [33] ), .ZN(_01834_ ) );
OAI21_X1 _09315_ ( .A(_01758_ ), .B1(_01833_ ), .B2(\myclint.mtime [33] ), .ZN(_01835_ ) );
NOR2_X1 _09316_ ( .A1(_01834_ ), .A2(_01835_ ), .ZN(_00025_ ) );
AND4_X1 _09317_ ( .A1(_01680_ ), .A2(_01733_ ), .A3(_01681_ ), .A4(_01735_ ), .ZN(_01836_ ) );
AND2_X1 _09318_ ( .A1(_01739_ ), .A2(_01742_ ), .ZN(_01837_ ) );
NAND3_X1 _09319_ ( .A1(_01836_ ), .A2(_01815_ ), .A3(_01837_ ), .ZN(_01838_ ) );
OAI21_X1 _09320_ ( .A(\myclint.mtime [32] ), .B1(_01736_ ), .B2(_01743_ ), .ZN(_01839_ ) );
AOI21_X1 _09321_ ( .A(fanout_net_1 ), .B1(_01838_ ), .B2(_01839_ ), .ZN(_00026_ ) );
AND2_X1 _09322_ ( .A1(_01837_ ), .A2(_01733_ ), .ZN(_01840_ ) );
NAND3_X1 _09323_ ( .A1(_01840_ ), .A2(_01681_ ), .A3(_01735_ ), .ZN(_01841_ ) );
OR3_X1 _09324_ ( .A1(_01841_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [31] ), .ZN(_01842_ ) );
OAI21_X1 _09325_ ( .A(\myclint.mtime [31] ), .B1(_01841_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01843_ ) );
AOI21_X1 _09326_ ( .A(fanout_net_1 ), .B1(_01842_ ), .B2(_01843_ ), .ZN(_00027_ ) );
OR2_X1 _09327_ ( .A1(_01841_ ), .A2(\myclint.mtime [30] ), .ZN(_01844_ ) );
NAND2_X1 _09328_ ( .A1(_01841_ ), .A2(\myclint.mtime [30] ), .ZN(_01845_ ) );
AOI21_X1 _09329_ ( .A(fanout_net_1 ), .B1(_01844_ ), .B2(_01845_ ), .ZN(_00028_ ) );
INV_X1 _09330_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01846_ ) );
AND3_X1 _09331_ ( .A1(_01678_ ), .A2(_01846_ ), .A3(\myclint.mtime [27] ), .ZN(_01847_ ) );
AND2_X1 _09332_ ( .A1(_01847_ ), .A2(\myclint.mtime [29] ), .ZN(_01848_ ) );
OAI21_X1 _09333_ ( .A(_01665_ ), .B1(_01847_ ), .B2(\myclint.mtime [29] ), .ZN(_01849_ ) );
NOR2_X1 _09334_ ( .A1(_01848_ ), .A2(_01849_ ), .ZN(_00029_ ) );
NAND2_X1 _09335_ ( .A1(_01840_ ), .A2(_01735_ ), .ZN(_01850_ ) );
OR2_X1 _09336_ ( .A1(_01850_ ), .A2(\myclint.mtime [28] ), .ZN(_01851_ ) );
NAND2_X1 _09337_ ( .A1(_01850_ ), .A2(\myclint.mtime [28] ), .ZN(_01852_ ) );
AOI21_X1 _09338_ ( .A(fanout_net_1 ), .B1(_01851_ ), .B2(_01852_ ), .ZN(_00030_ ) );
INV_X1 _09339_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01853_ ) );
AND3_X1 _09340_ ( .A1(_01677_ ), .A2(_01853_ ), .A3(\myclint.mtime [25] ), .ZN(_01854_ ) );
AND2_X1 _09341_ ( .A1(_01854_ ), .A2(\myclint.mtime [27] ), .ZN(_01855_ ) );
OAI21_X1 _09342_ ( .A(_01665_ ), .B1(_01854_ ), .B2(\myclint.mtime [27] ), .ZN(_01856_ ) );
NOR2_X1 _09343_ ( .A1(_01855_ ), .A2(_01856_ ), .ZN(_00031_ ) );
BUF_X4 _09344_ ( .A(_01664_ ), .Z(_01857_ ) );
AND2_X1 _09345_ ( .A1(_01677_ ), .A2(\myclint.mtime [25] ), .ZN(_01858_ ) );
OAI21_X1 _09346_ ( .A(_01857_ ), .B1(_01858_ ), .B2(\myclint.mtime [26] ), .ZN(_01859_ ) );
NOR2_X1 _09347_ ( .A1(_01859_ ), .A2(_01678_ ), .ZN(_00032_ ) );
INV_X1 _09348_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01860_ ) );
AND3_X1 _09349_ ( .A1(_01676_ ), .A2(_01860_ ), .A3(\myclint.mtime [23] ), .ZN(_01861_ ) );
AND2_X1 _09350_ ( .A1(_01861_ ), .A2(\myclint.mtime [25] ), .ZN(_01862_ ) );
OAI21_X1 _09351_ ( .A(_01665_ ), .B1(_01861_ ), .B2(\myclint.mtime [25] ), .ZN(_01863_ ) );
NOR2_X1 _09352_ ( .A1(_01862_ ), .A2(_01863_ ), .ZN(_00033_ ) );
AND2_X1 _09353_ ( .A1(_01676_ ), .A2(\myclint.mtime [23] ), .ZN(_01864_ ) );
OAI21_X1 _09354_ ( .A(_01857_ ), .B1(_01864_ ), .B2(\myclint.mtime [24] ), .ZN(_01865_ ) );
NOR2_X1 _09355_ ( .A1(_01865_ ), .A2(_01677_ ), .ZN(_00034_ ) );
INV_X1 _09356_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01866_ ) );
AND4_X1 _09357_ ( .A1(_01866_ ), .A2(_01725_ ), .A3(\myclint.mtime [59] ), .A4(_01703_ ), .ZN(_01867_ ) );
AND3_X1 _09358_ ( .A1(_01702_ ), .A2(_01866_ ), .A3(_01703_ ), .ZN(_01868_ ) );
OAI21_X1 _09359_ ( .A(_01665_ ), .B1(_01868_ ), .B2(\myclint.mtime [59] ), .ZN(_01869_ ) );
NOR2_X1 _09360_ ( .A1(_01867_ ), .A2(_01869_ ), .ZN(_00035_ ) );
AND2_X1 _09361_ ( .A1(_01837_ ), .A2(_01731_ ), .ZN(_01870_ ) );
NAND3_X1 _09362_ ( .A1(_01870_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01871_ ) );
OR3_X1 _09363_ ( .A1(_01871_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01872_ ) );
OAI21_X1 _09364_ ( .A(\myclint.mtime [23] ), .B1(_01871_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01873_ ) );
AOI21_X1 _09365_ ( .A(fanout_net_1 ), .B1(_01872_ ), .B2(_01873_ ), .ZN(_00036_ ) );
AND2_X1 _09366_ ( .A1(_01675_ ), .A2(\myclint.mtime [21] ), .ZN(_01874_ ) );
OAI21_X1 _09367_ ( .A(_01857_ ), .B1(_01874_ ), .B2(\myclint.mtime [22] ), .ZN(_01875_ ) );
NOR2_X1 _09368_ ( .A1(_01875_ ), .A2(_01676_ ), .ZN(_00037_ ) );
INV_X1 _09369_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01876_ ) );
AND3_X1 _09370_ ( .A1(_01674_ ), .A2(_01876_ ), .A3(\myclint.mtime [19] ), .ZN(_01877_ ) );
AND2_X1 _09371_ ( .A1(_01877_ ), .A2(\myclint.mtime [21] ), .ZN(_01878_ ) );
OAI21_X1 _09372_ ( .A(_01665_ ), .B1(_01877_ ), .B2(\myclint.mtime [21] ), .ZN(_01879_ ) );
NOR2_X1 _09373_ ( .A1(_01878_ ), .A2(_01879_ ), .ZN(_00038_ ) );
AND2_X1 _09374_ ( .A1(_01674_ ), .A2(\myclint.mtime [19] ), .ZN(_01880_ ) );
OAI21_X1 _09375_ ( .A(_01857_ ), .B1(_01880_ ), .B2(\myclint.mtime [20] ), .ZN(_01881_ ) );
NOR2_X1 _09376_ ( .A1(_01881_ ), .A2(_01675_ ), .ZN(_00039_ ) );
NAND3_X1 _09377_ ( .A1(_01837_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01882_ ) );
OR3_X1 _09378_ ( .A1(_01882_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01883_ ) );
OAI21_X1 _09379_ ( .A(\myclint.mtime [19] ), .B1(_01882_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01884_ ) );
AOI21_X1 _09380_ ( .A(fanout_net_1 ), .B1(_01883_ ), .B2(_01884_ ), .ZN(_00040_ ) );
AND2_X1 _09381_ ( .A1(_01673_ ), .A2(\myclint.mtime [17] ), .ZN(_01885_ ) );
OAI21_X1 _09382_ ( .A(_01857_ ), .B1(_01885_ ), .B2(\myclint.mtime [18] ), .ZN(_01886_ ) );
NOR2_X1 _09383_ ( .A1(_01886_ ), .A2(_01674_ ), .ZN(_00041_ ) );
INV_X1 _09384_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01887_ ) );
AND3_X1 _09385_ ( .A1(_01672_ ), .A2(_01887_ ), .A3(\myclint.mtime [15] ), .ZN(_01888_ ) );
AND2_X1 _09386_ ( .A1(_01888_ ), .A2(\myclint.mtime [17] ), .ZN(_01889_ ) );
OAI21_X1 _09387_ ( .A(_01665_ ), .B1(_01888_ ), .B2(\myclint.mtime [17] ), .ZN(_01890_ ) );
NOR2_X1 _09388_ ( .A1(_01889_ ), .A2(_01890_ ), .ZN(_00042_ ) );
AND2_X1 _09389_ ( .A1(_01672_ ), .A2(\myclint.mtime [15] ), .ZN(_01891_ ) );
OAI21_X1 _09390_ ( .A(_01857_ ), .B1(_01891_ ), .B2(\myclint.mtime [16] ), .ZN(_01892_ ) );
NOR2_X1 _09391_ ( .A1(_01892_ ), .A2(_01673_ ), .ZN(_00043_ ) );
AND3_X1 _09392_ ( .A1(_01741_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01893_ ) );
AND2_X1 _09393_ ( .A1(_01739_ ), .A2(_01893_ ), .ZN(_01894_ ) );
NAND3_X1 _09394_ ( .A1(_01894_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01895_ ) );
OR3_X1 _09395_ ( .A1(_01895_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01896_ ) );
OAI21_X1 _09396_ ( .A(\myclint.mtime [15] ), .B1(_01895_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01897_ ) );
AOI21_X1 _09397_ ( .A(fanout_net_1 ), .B1(_01896_ ), .B2(_01897_ ), .ZN(_00044_ ) );
AND2_X1 _09398_ ( .A1(_01671_ ), .A2(\myclint.mtime [13] ), .ZN(_01898_ ) );
OAI21_X1 _09399_ ( .A(_01857_ ), .B1(_01898_ ), .B2(\myclint.mtime [14] ), .ZN(_01899_ ) );
NOR2_X1 _09400_ ( .A1(_01899_ ), .A2(_01672_ ), .ZN(_00045_ ) );
NAND3_X1 _09401_ ( .A1(_01749_ ), .A2(_01703_ ), .A3(_01750_ ), .ZN(_01900_ ) );
OR2_X1 _09402_ ( .A1(_01900_ ), .A2(\myclint.mtime [58] ), .ZN(_01901_ ) );
NAND2_X1 _09403_ ( .A1(_01900_ ), .A2(\myclint.mtime [58] ), .ZN(_01902_ ) );
AOI21_X1 _09404_ ( .A(fanout_net_1 ), .B1(_01901_ ), .B2(_01902_ ), .ZN(_00046_ ) );
INV_X1 _09405_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01903_ ) );
NAND3_X1 _09406_ ( .A1(_01739_ ), .A2(_01903_ ), .A3(_01893_ ), .ZN(_01904_ ) );
OR2_X1 _09407_ ( .A1(_01904_ ), .A2(\myclint.mtime [13] ), .ZN(_01905_ ) );
NAND2_X1 _09408_ ( .A1(_01904_ ), .A2(\myclint.mtime [13] ), .ZN(_01906_ ) );
AOI21_X1 _09409_ ( .A(fanout_net_1 ), .B1(_01905_ ), .B2(_01906_ ), .ZN(_00047_ ) );
AND2_X1 _09410_ ( .A1(_01670_ ), .A2(\myclint.mtime [11] ), .ZN(_01907_ ) );
OAI21_X1 _09411_ ( .A(_01857_ ), .B1(_01907_ ), .B2(\myclint.mtime [12] ), .ZN(_01908_ ) );
NOR2_X1 _09412_ ( .A1(_01908_ ), .A2(_01671_ ), .ZN(_00048_ ) );
NAND3_X1 _09413_ ( .A1(_01739_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01909_ ) );
OR3_X1 _09414_ ( .A1(_01909_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_01910_ ) );
OAI21_X1 _09415_ ( .A(\myclint.mtime [11] ), .B1(_01909_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01911_ ) );
AOI21_X1 _09416_ ( .A(fanout_net_1 ), .B1(_01910_ ), .B2(_01911_ ), .ZN(_00049_ ) );
AND2_X1 _09417_ ( .A1(_01669_ ), .A2(\myclint.mtime [9] ), .ZN(_01912_ ) );
OAI21_X1 _09418_ ( .A(_01857_ ), .B1(_01912_ ), .B2(\myclint.mtime [10] ), .ZN(_01913_ ) );
NOR2_X1 _09419_ ( .A1(_01913_ ), .A2(_01670_ ), .ZN(_00050_ ) );
AND2_X1 _09420_ ( .A1(_01668_ ), .A2(\myclint.mtime [7] ), .ZN(_01914_ ) );
INV_X1 _09421_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01915_ ) );
AND3_X1 _09422_ ( .A1(_01914_ ), .A2(\myclint.mtime [9] ), .A3(_01915_ ), .ZN(_01916_ ) );
AOI21_X1 _09423_ ( .A(\myclint.mtime [9] ), .B1(_01914_ ), .B2(_01915_ ), .ZN(_01917_ ) );
NOR3_X1 _09424_ ( .A1(_01916_ ), .A2(_01917_ ), .A3(fanout_net_1 ), .ZN(_00051_ ) );
OAI21_X1 _09425_ ( .A(_01857_ ), .B1(_01914_ ), .B2(\myclint.mtime [8] ), .ZN(_01918_ ) );
NOR2_X1 _09426_ ( .A1(_01918_ ), .A2(_01669_ ), .ZN(_00052_ ) );
AND2_X1 _09427_ ( .A1(_01667_ ), .A2(\myclint.mtime [5] ), .ZN(_01919_ ) );
INV_X1 _09428_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01920_ ) );
AND3_X1 _09429_ ( .A1(_01919_ ), .A2(_01920_ ), .A3(\myclint.mtime [7] ), .ZN(_01921_ ) );
AOI21_X1 _09430_ ( .A(\myclint.mtime [7] ), .B1(_01919_ ), .B2(_01920_ ), .ZN(_01922_ ) );
NOR3_X1 _09431_ ( .A1(_01921_ ), .A2(_01922_ ), .A3(fanout_net_1 ), .ZN(_00053_ ) );
OAI21_X1 _09432_ ( .A(_01758_ ), .B1(_01919_ ), .B2(\myclint.mtime [6] ), .ZN(_01923_ ) );
NOR2_X1 _09433_ ( .A1(_01923_ ), .A2(_01668_ ), .ZN(_00054_ ) );
INV_X1 _09434_ ( .A(_01737_ ), .ZN(_01924_ ) );
OR3_X1 _09435_ ( .A1(_01924_ ), .A2(\myclint.mtime [5] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01925_ ) );
OAI21_X1 _09436_ ( .A(\myclint.mtime [5] ), .B1(_01924_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01926_ ) );
AOI21_X1 _09437_ ( .A(fanout_net_1 ), .B1(_01925_ ), .B2(_01926_ ), .ZN(_00055_ ) );
OAI21_X1 _09438_ ( .A(_01758_ ), .B1(_01737_ ), .B2(\myclint.mtime [4] ), .ZN(_01927_ ) );
NOR2_X1 _09439_ ( .A1(_01927_ ), .A2(_01667_ ), .ZN(_00056_ ) );
INV_X1 _09440_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01928_ ) );
AND4_X1 _09441_ ( .A1(\myclint.mtime [57] ), .A2(_01724_ ), .A3(_01928_ ), .A4(_01701_ ), .ZN(_01929_ ) );
AND3_X1 _09442_ ( .A1(_01700_ ), .A2(_01928_ ), .A3(_01701_ ), .ZN(_01930_ ) );
OAI21_X1 _09443_ ( .A(_01665_ ), .B1(_01930_ ), .B2(\myclint.mtime [57] ), .ZN(_01931_ ) );
NOR2_X1 _09444_ ( .A1(_01929_ ), .A2(_01931_ ), .ZN(_00057_ ) );
AND2_X1 _09445_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01932_ ) );
INV_X1 _09446_ ( .A(_01932_ ), .ZN(_01933_ ) );
OR3_X1 _09447_ ( .A1(_01933_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01934_ ) );
OAI21_X1 _09448_ ( .A(\myclint.mtime [3] ), .B1(_01933_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01935_ ) );
AOI21_X1 _09449_ ( .A(fanout_net_1 ), .B1(_01934_ ), .B2(_01935_ ), .ZN(_00058_ ) );
AOI21_X1 _09450_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01936_ ) );
NOR3_X1 _09451_ ( .A1(_01666_ ), .A2(_01936_ ), .A3(fanout_net_1 ), .ZN(_00059_ ) );
NOR2_X1 _09452_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01937_ ) );
NOR3_X1 _09453_ ( .A1(_01932_ ), .A2(_01937_ ), .A3(fanout_net_1 ), .ZN(_00060_ ) );
INV_X1 _09454_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_01938_ ) );
NOR2_X1 _09455_ ( .A1(_01938_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
XNOR2_X1 _09456_ ( .A(_01751_ ), .B(\myclint.mtime [56] ), .ZN(_01939_ ) );
NOR2_X1 _09457_ ( .A1(_01939_ ), .A2(fanout_net_2 ), .ZN(_00062_ ) );
NAND2_X1 _09458_ ( .A1(_01698_ ), .A2(_01699_ ), .ZN(_01940_ ) );
NOR2_X1 _09459_ ( .A1(_01940_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01941_ ) );
OAI21_X1 _09460_ ( .A(_01664_ ), .B1(_01941_ ), .B2(\myclint.mtime [55] ), .ZN(_01942_ ) );
INV_X1 _09461_ ( .A(_01724_ ), .ZN(_01943_ ) );
NOR2_X1 _09462_ ( .A1(_01943_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01944_ ) );
AOI21_X1 _09463_ ( .A(_01942_ ), .B1(_01944_ ), .B2(\myclint.mtime [55] ), .ZN(_00063_ ) );
NAND3_X1 _09464_ ( .A1(_01749_ ), .A2(_01699_ ), .A3(_01761_ ), .ZN(_01945_ ) );
OR2_X1 _09465_ ( .A1(_01945_ ), .A2(\myclint.mtime [54] ), .ZN(_01946_ ) );
NAND2_X1 _09466_ ( .A1(_01945_ ), .A2(\myclint.mtime [54] ), .ZN(_01947_ ) );
AOI21_X1 _09467_ ( .A(fanout_net_2 ), .B1(_01946_ ), .B2(_01947_ ), .ZN(_00064_ ) );
MUX2_X1 _09468_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(fanout_net_42 ), .Z(_01948_ ) );
MUX2_X1 _09469_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(fanout_net_42 ), .Z(_01949_ ) );
MUX2_X2 _09470_ ( .A(_01948_ ), .B(_01949_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01950_ ) );
INV_X1 _09471_ ( .A(\IF_ID_pc [21] ), .ZN(_01951_ ) );
MUX2_X1 _09472_ ( .A(\myifu.myicache.tag[0][4] ), .B(\myifu.myicache.tag[1][4] ), .S(fanout_net_42 ), .Z(_01952_ ) );
INV_X32 _09473_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01953_ ) );
BUF_X32 _09474_ ( .A(_01953_ ), .Z(_01954_ ) );
BUF_X16 _09475_ ( .A(_01954_ ), .Z(_01955_ ) );
NAND2_X1 _09476_ ( .A1(_01952_ ), .A2(_01955_ ), .ZN(_01956_ ) );
MUX2_X1 _09477_ ( .A(\myifu.myicache.tag[2][4] ), .B(\myifu.myicache.tag[3][4] ), .S(fanout_net_42 ), .Z(_01957_ ) );
NAND2_X1 _09478_ ( .A1(_01957_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01958_ ) );
NAND2_X1 _09479_ ( .A1(_01956_ ), .A2(_01958_ ), .ZN(_01959_ ) );
INV_X1 _09480_ ( .A(\IF_ID_pc [9] ), .ZN(_01960_ ) );
AOI22_X1 _09481_ ( .A1(_01950_ ), .A2(_01951_ ), .B1(_01959_ ), .B2(_01960_ ), .ZN(_01961_ ) );
INV_X32 _09482_ ( .A(fanout_net_42 ), .ZN(_01962_ ) );
OR2_X1 _09483_ ( .A1(_01962_ ), .A2(\myifu.myicache.tag[1][2] ), .ZN(_01963_ ) );
OAI211_X1 _09484_ ( .A(_01963_ ), .B(_01954_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][2] ), .ZN(_01964_ ) );
OR2_X1 _09485_ ( .A1(_01962_ ), .A2(\myifu.myicache.tag[3][2] ), .ZN(_01965_ ) );
OAI211_X1 _09486_ ( .A(_01965_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[2][2] ), .ZN(_01966_ ) );
NAND2_X1 _09487_ ( .A1(_01964_ ), .A2(_01966_ ), .ZN(_01967_ ) );
INV_X1 _09488_ ( .A(_01967_ ), .ZN(_01968_ ) );
OAI221_X1 _09489_ ( .A(_01961_ ), .B1(_01960_ ), .B2(_01959_ ), .C1(\IF_ID_pc [7] ), .C2(_01968_ ), .ZN(_01969_ ) );
MUX2_X1 _09490_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(fanout_net_42 ), .Z(_01970_ ) );
OR2_X1 _09491_ ( .A1(_01970_ ), .A2(_01955_ ), .ZN(_01971_ ) );
MUX2_X1 _09492_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(fanout_net_42 ), .Z(_01972_ ) );
OAI21_X1 _09493_ ( .A(_01971_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01972_ ), .ZN(_01973_ ) );
NAND2_X1 _09494_ ( .A1(_01973_ ), .A2(\IF_ID_pc [20] ), .ZN(_01974_ ) );
INV_X1 _09495_ ( .A(\IF_ID_pc [12] ), .ZN(_01975_ ) );
MUX2_X1 _09496_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(fanout_net_42 ), .Z(_01976_ ) );
MUX2_X1 _09497_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(fanout_net_42 ), .Z(_01977_ ) );
MUX2_X1 _09498_ ( .A(_01976_ ), .B(_01977_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01978_ ) );
OAI21_X1 _09499_ ( .A(_01974_ ), .B1(_01975_ ), .B2(_01978_ ), .ZN(_01979_ ) );
MUX2_X1 _09500_ ( .A(\myifu.myicache.tag[0][3] ), .B(\myifu.myicache.tag[1][3] ), .S(fanout_net_42 ), .Z(_01980_ ) );
MUX2_X1 _09501_ ( .A(\myifu.myicache.tag[2][3] ), .B(\myifu.myicache.tag[3][3] ), .S(fanout_net_42 ), .Z(_01981_ ) );
MUX2_X2 _09502_ ( .A(_01980_ ), .B(_01981_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01982_ ) );
INV_X1 _09503_ ( .A(\IF_ID_pc [8] ), .ZN(_01983_ ) );
NOR2_X1 _09504_ ( .A1(_01982_ ), .A2(_01983_ ), .ZN(_01984_ ) );
AND2_X1 _09505_ ( .A1(_01978_ ), .A2(_01975_ ), .ZN(_01985_ ) );
NOR4_X1 _09506_ ( .A1(_01969_ ), .A2(_01979_ ), .A3(_01984_ ), .A4(_01985_ ), .ZN(_01986_ ) );
OR2_X4 _09507_ ( .A1(_01962_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01987_ ) );
OAI211_X1 _09508_ ( .A(_01987_ ), .B(_01953_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01988_ ) );
OR2_X4 _09509_ ( .A1(fanout_net_42 ), .A2(\myifu.myicache.tag[2][12] ), .ZN(_01989_ ) );
OAI211_X1 _09510_ ( .A(_01989_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01962_ ), .C2(\myifu.myicache.tag[3][12] ), .ZN(_01990_ ) );
NAND2_X1 _09511_ ( .A1(_01988_ ), .A2(_01990_ ), .ZN(_01991_ ) );
INV_X1 _09512_ ( .A(_01991_ ), .ZN(_01992_ ) );
INV_X1 _09513_ ( .A(\IF_ID_pc [15] ), .ZN(_01993_ ) );
OR2_X1 _09514_ ( .A1(fanout_net_42 ), .A2(\myifu.myicache.tag[0][10] ), .ZN(_01994_ ) );
OAI211_X1 _09515_ ( .A(_01994_ ), .B(_01954_ ), .C1(_01962_ ), .C2(\myifu.myicache.tag[1][10] ), .ZN(_01995_ ) );
OR2_X1 _09516_ ( .A1(fanout_net_42 ), .A2(\myifu.myicache.tag[2][10] ), .ZN(_01996_ ) );
OAI211_X1 _09517_ ( .A(_01996_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01962_ ), .C2(\myifu.myicache.tag[3][10] ), .ZN(_01997_ ) );
NAND2_X1 _09518_ ( .A1(_01995_ ), .A2(_01997_ ), .ZN(_01998_ ) );
OAI22_X1 _09519_ ( .A1(_01992_ ), .A2(\IF_ID_pc [17] ), .B1(_01993_ ), .B2(_01998_ ), .ZN(_01999_ ) );
AOI221_X1 _09520_ ( .A(_01999_ ), .B1(_01993_ ), .B2(_01998_ ), .C1(\IF_ID_pc [7] ), .C2(_01968_ ), .ZN(_02000_ ) );
MUX2_X1 _09521_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(fanout_net_42 ), .Z(_02001_ ) );
MUX2_X1 _09522_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_42 ), .Z(_02002_ ) );
MUX2_X2 _09523_ ( .A(_02001_ ), .B(_02002_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02003_ ) );
INV_X1 _09524_ ( .A(\IF_ID_pc [25] ), .ZN(_02004_ ) );
OR2_X1 _09525_ ( .A1(_02003_ ), .A2(_02004_ ), .ZN(_02005_ ) );
MUX2_X1 _09526_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_42 ), .Z(_02006_ ) );
OR2_X1 _09527_ ( .A1(_02006_ ), .A2(_01955_ ), .ZN(_02007_ ) );
MUX2_X1 _09528_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_42 ), .Z(_02008_ ) );
OAI21_X1 _09529_ ( .A(_02007_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_02008_ ), .ZN(_02009_ ) );
NAND2_X1 _09530_ ( .A1(_02009_ ), .A2(\IF_ID_pc [16] ), .ZN(_02010_ ) );
MUX2_X1 _09531_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(fanout_net_42 ), .Z(_02011_ ) );
OR2_X2 _09532_ ( .A1(_02011_ ), .A2(_01954_ ), .ZN(_02012_ ) );
MUX2_X1 _09533_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(fanout_net_42 ), .Z(_02013_ ) );
OAI21_X1 _09534_ ( .A(_02012_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_02013_ ), .ZN(_02014_ ) );
AOI22_X1 _09535_ ( .A1(_02014_ ), .A2(\IF_ID_pc [27] ), .B1(_01992_ ), .B2(\IF_ID_pc [17] ), .ZN(_02015_ ) );
AND4_X1 _09536_ ( .A1(_02000_ ), .A2(_02005_ ), .A3(_02010_ ), .A4(_02015_ ), .ZN(_02016_ ) );
MUX2_X1 _09537_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(fanout_net_42 ), .Z(_02017_ ) );
OR2_X2 _09538_ ( .A1(_02017_ ), .A2(_01954_ ), .ZN(_02018_ ) );
MUX2_X1 _09539_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(fanout_net_42 ), .Z(_02019_ ) );
OAI21_X1 _09540_ ( .A(_02018_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_02019_ ), .ZN(_02020_ ) );
INV_X1 _09541_ ( .A(_02020_ ), .ZN(_02021_ ) );
INV_X1 _09542_ ( .A(\IF_ID_pc [10] ), .ZN(_02022_ ) );
AOI22_X1 _09543_ ( .A1(_02021_ ), .A2(_02022_ ), .B1(_01983_ ), .B2(_01982_ ), .ZN(_02023_ ) );
INV_X1 _09544_ ( .A(\IF_ID_pc [14] ), .ZN(_02024_ ) );
MUX2_X1 _09545_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(fanout_net_42 ), .Z(_02025_ ) );
MUX2_X1 _09546_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(fanout_net_42 ), .Z(_02026_ ) );
MUX2_X2 _09547_ ( .A(_02025_ ), .B(_02026_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02027_ ) );
OAI221_X1 _09548_ ( .A(_02023_ ), .B1(_02024_ ), .B2(_02027_ ), .C1(\IF_ID_pc [16] ), .C2(_02009_ ), .ZN(_02028_ ) );
MUX2_X1 _09549_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(fanout_net_42 ), .Z(_02029_ ) );
MUX2_X1 _09550_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(fanout_net_42 ), .Z(_02030_ ) );
MUX2_X1 _09551_ ( .A(_02029_ ), .B(_02030_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02031_ ) );
INV_X1 _09552_ ( .A(\IF_ID_pc [23] ), .ZN(_02032_ ) );
OR2_X2 _09553_ ( .A1(_02031_ ), .A2(_02032_ ), .ZN(_02033_ ) );
OAI221_X1 _09554_ ( .A(_02033_ ), .B1(_01951_ ), .B2(_01950_ ), .C1(_02021_ ), .C2(_02022_ ), .ZN(_02034_ ) );
NOR2_X1 _09555_ ( .A1(_02028_ ), .A2(_02034_ ), .ZN(_02035_ ) );
MUX2_X1 _09556_ ( .A(\myifu.myicache.tag[2][8] ), .B(\myifu.myicache.tag[3][8] ), .S(fanout_net_42 ), .Z(_02036_ ) );
AND2_X1 _09557_ ( .A1(_02036_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_02037_ ) );
MUX2_X1 _09558_ ( .A(\myifu.myicache.tag[0][8] ), .B(\myifu.myicache.tag[1][8] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02038_ ) );
AOI21_X1 _09559_ ( .A(_02037_ ), .B1(_01955_ ), .B2(_02038_ ), .ZN(_02039_ ) );
AOI22_X1 _09560_ ( .A1(_02039_ ), .A2(\IF_ID_pc [13] ), .B1(_02004_ ), .B2(_02003_ ), .ZN(_02040_ ) );
NAND2_X1 _09561_ ( .A1(_02031_ ), .A2(_02032_ ), .ZN(_02041_ ) );
INV_X1 _09562_ ( .A(\IF_ID_pc [31] ), .ZN(_02042_ ) );
MUX2_X1 _09563_ ( .A(\myifu.myicache.tag[0][26] ), .B(\myifu.myicache.tag[1][26] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02043_ ) );
MUX2_X1 _09564_ ( .A(\myifu.myicache.tag[2][26] ), .B(\myifu.myicache.tag[3][26] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02044_ ) );
MUX2_X1 _09565_ ( .A(_02043_ ), .B(_02044_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02045_ ) );
OAI211_X1 _09566_ ( .A(_02040_ ), .B(_02041_ ), .C1(_02042_ ), .C2(_02045_ ), .ZN(_02046_ ) );
AND2_X1 _09567_ ( .A1(_02045_ ), .A2(_02042_ ), .ZN(_02047_ ) );
NOR2_X1 _09568_ ( .A1(_02039_ ), .A2(\IF_ID_pc [13] ), .ZN(_02048_ ) );
NAND2_X1 _09569_ ( .A1(_02027_ ), .A2(_02024_ ), .ZN(_02049_ ) );
OAI21_X1 _09570_ ( .A(_02049_ ), .B1(_01973_ ), .B2(\IF_ID_pc [20] ), .ZN(_02050_ ) );
NOR4_X2 _09571_ ( .A1(_02046_ ), .A2(_02047_ ), .A3(_02048_ ), .A4(_02050_ ), .ZN(_02051_ ) );
AND4_X2 _09572_ ( .A1(_01986_ ), .A2(_02016_ ), .A3(_02035_ ), .A4(_02051_ ), .ZN(_02052_ ) );
BUF_X16 _09573_ ( .A(_01962_ ), .Z(_02053_ ) );
OR2_X4 _09574_ ( .A1(_02053_ ), .A2(\myifu.myicache.tag[3][23] ), .ZN(_02054_ ) );
OAI211_X1 _09575_ ( .A(_02054_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][23] ), .ZN(_02055_ ) );
INV_X1 _09576_ ( .A(\IF_ID_pc [28] ), .ZN(_02056_ ) );
OR2_X1 _09577_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][23] ), .ZN(_02057_ ) );
OAI211_X1 _09578_ ( .A(_02057_ ), .B(_01955_ ), .C1(_02053_ ), .C2(\myifu.myicache.tag[1][23] ), .ZN(_02058_ ) );
AND3_X1 _09579_ ( .A1(_02055_ ), .A2(_02056_ ), .A3(_02058_ ), .ZN(_02059_ ) );
AOI21_X1 _09580_ ( .A(_02056_ ), .B1(_02055_ ), .B2(_02058_ ), .ZN(_02060_ ) );
BUF_X32 _09581_ ( .A(_01962_ ), .Z(_02061_ ) );
OR2_X4 _09582_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[3][14] ), .ZN(_02062_ ) );
OAI211_X1 _09583_ ( .A(_02062_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][14] ), .ZN(_02063_ ) );
INV_X1 _09584_ ( .A(\IF_ID_pc [19] ), .ZN(_02064_ ) );
OR2_X1 _09585_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][14] ), .ZN(_02065_ ) );
OAI211_X1 _09586_ ( .A(_02065_ ), .B(_01955_ ), .C1(_02053_ ), .C2(\myifu.myicache.tag[1][14] ), .ZN(_02066_ ) );
AND3_X1 _09587_ ( .A1(_02063_ ), .A2(_02064_ ), .A3(_02066_ ), .ZN(_02067_ ) );
AOI21_X1 _09588_ ( .A(_02064_ ), .B1(_02063_ ), .B2(_02066_ ), .ZN(_02068_ ) );
OAI22_X1 _09589_ ( .A1(_02059_ ), .A2(_02060_ ), .B1(_02067_ ), .B2(_02068_ ), .ZN(_02069_ ) );
OR2_X4 _09590_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[1][0] ), .ZN(_02070_ ) );
OAI211_X2 _09591_ ( .A(_02070_ ), .B(_01954_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][0] ), .ZN(_02071_ ) );
OR2_X4 _09592_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[3][0] ), .ZN(_02072_ ) );
OAI211_X2 _09593_ ( .A(_02072_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][0] ), .ZN(_02073_ ) );
AND2_X4 _09594_ ( .A1(_02071_ ), .A2(_02073_ ), .ZN(_02074_ ) );
XOR2_X2 _09595_ ( .A(_02074_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .Z(_02075_ ) );
OR2_X4 _09596_ ( .A1(_02053_ ), .A2(\myifu.myicache.tag[1][17] ), .ZN(_02076_ ) );
OAI211_X1 _09597_ ( .A(_02076_ ), .B(_01955_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][17] ), .ZN(_02077_ ) );
OR2_X1 _09598_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][17] ), .ZN(_02078_ ) );
OAI211_X1 _09599_ ( .A(_02078_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02053_ ), .C2(\myifu.myicache.tag[3][17] ), .ZN(_02079_ ) );
AND3_X1 _09600_ ( .A1(_02077_ ), .A2(_02079_ ), .A3(\IF_ID_pc [22] ), .ZN(_02080_ ) );
AOI21_X1 _09601_ ( .A(\IF_ID_pc [22] ), .B1(_02077_ ), .B2(_02079_ ), .ZN(_02081_ ) );
OR4_X2 _09602_ ( .A1(_02069_ ), .A2(_02075_ ), .A3(_02080_ ), .A4(_02081_ ), .ZN(_02082_ ) );
OR2_X4 _09603_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[1][24] ), .ZN(_02083_ ) );
OAI211_X2 _09604_ ( .A(_02083_ ), .B(_01954_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][24] ), .ZN(_02084_ ) );
OR2_X4 _09605_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[3][24] ), .ZN(_02085_ ) );
OAI211_X2 _09606_ ( .A(_02085_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][24] ), .ZN(_02086_ ) );
INV_X1 _09607_ ( .A(\IF_ID_pc [29] ), .ZN(_02087_ ) );
AND3_X1 _09608_ ( .A1(_02084_ ), .A2(_02086_ ), .A3(_02087_ ), .ZN(_02088_ ) );
AOI21_X1 _09609_ ( .A(_02087_ ), .B1(_02084_ ), .B2(_02086_ ), .ZN(_02089_ ) );
OR2_X4 _09610_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[3][6] ), .ZN(_02090_ ) );
OAI211_X2 _09611_ ( .A(_02090_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][6] ), .ZN(_02091_ ) );
INV_X1 _09612_ ( .A(\IF_ID_pc [11] ), .ZN(_02092_ ) );
OR2_X1 _09613_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][6] ), .ZN(_02093_ ) );
OAI211_X1 _09614_ ( .A(_02093_ ), .B(_01954_ ), .C1(_02053_ ), .C2(\myifu.myicache.tag[1][6] ), .ZN(_02094_ ) );
AND3_X1 _09615_ ( .A1(_02091_ ), .A2(_02092_ ), .A3(_02094_ ), .ZN(_02095_ ) );
AOI21_X1 _09616_ ( .A(_02092_ ), .B1(_02091_ ), .B2(_02094_ ), .ZN(_02096_ ) );
OAI22_X1 _09617_ ( .A1(_02088_ ), .A2(_02089_ ), .B1(_02095_ ), .B2(_02096_ ), .ZN(_02097_ ) );
OR2_X4 _09618_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_02098_ ) );
OAI211_X2 _09619_ ( .A(_02098_ ), .B(_01954_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_02099_ ) );
OR2_X4 _09620_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[3][25] ), .ZN(_02100_ ) );
OAI211_X4 _09621_ ( .A(_02100_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][25] ), .ZN(_02101_ ) );
NAND2_X2 _09622_ ( .A1(_02099_ ), .A2(_02101_ ), .ZN(_02102_ ) );
XOR2_X1 _09623_ ( .A(_02102_ ), .B(\IF_ID_pc [30] ), .Z(_02103_ ) );
OR2_X1 _09624_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[1][13] ), .ZN(_02104_ ) );
OAI211_X1 _09625_ ( .A(_02104_ ), .B(_01955_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][13] ), .ZN(_02105_ ) );
OR2_X2 _09626_ ( .A1(_02061_ ), .A2(\myifu.myicache.tag[3][13] ), .ZN(_02106_ ) );
OAI211_X1 _09627_ ( .A(_02106_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][13] ), .ZN(_02107_ ) );
AOI21_X1 _09628_ ( .A(\IF_ID_pc [18] ), .B1(_02105_ ), .B2(_02107_ ), .ZN(_02108_ ) );
AND3_X1 _09629_ ( .A1(_02105_ ), .A2(_02107_ ), .A3(\IF_ID_pc [18] ), .ZN(_02109_ ) );
OR4_X4 _09630_ ( .A1(_02097_ ), .A2(_02103_ ), .A3(_02108_ ), .A4(_02109_ ), .ZN(_02110_ ) );
INV_X1 _09631_ ( .A(\IF_ID_pc [26] ), .ZN(_02111_ ) );
MUX2_X1 _09632_ ( .A(\myifu.myicache.tag[2][21] ), .B(\myifu.myicache.tag[3][21] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02112_ ) );
OR2_X2 _09633_ ( .A1(_02112_ ), .A2(_01954_ ), .ZN(_02113_ ) );
MUX2_X1 _09634_ ( .A(\myifu.myicache.tag[0][21] ), .B(\myifu.myicache.tag[1][21] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02114_ ) );
OR2_X4 _09635_ ( .A1(_02114_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_02115_ ) );
AOI21_X1 _09636_ ( .A(_02111_ ), .B1(_02113_ ), .B2(_02115_ ), .ZN(_02116_ ) );
NOR2_X4 _09637_ ( .A1(_02014_ ), .A2(\IF_ID_pc [27] ), .ZN(_02117_ ) );
OR2_X4 _09638_ ( .A1(_02053_ ), .A2(\myifu.myicache.tag[1][19] ), .ZN(_02118_ ) );
OAI211_X1 _09639_ ( .A(_02118_ ), .B(_01955_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][19] ), .ZN(_02119_ ) );
OR2_X1 _09640_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][19] ), .ZN(_02120_ ) );
OAI211_X1 _09641_ ( .A(_02120_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02053_ ), .C2(\myifu.myicache.tag[3][19] ), .ZN(_02121_ ) );
AOI21_X1 _09642_ ( .A(\IF_ID_pc [24] ), .B1(_02119_ ), .B2(_02121_ ), .ZN(_02122_ ) );
AND3_X4 _09643_ ( .A1(_02113_ ), .A2(_02115_ ), .A3(_02111_ ), .ZN(_02123_ ) );
OR4_X4 _09644_ ( .A1(_02116_ ), .A2(_02117_ ), .A3(_02122_ ), .A4(_02123_ ), .ZN(_02124_ ) );
MUX2_X1 _09645_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02125_ ) );
MUX2_X1 _09646_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02126_ ) );
MUX2_X1 _09647_ ( .A(_02125_ ), .B(_02126_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02127_ ) );
NAND3_X1 _09648_ ( .A1(_02119_ ), .A2(_02121_ ), .A3(\IF_ID_pc [24] ), .ZN(_02128_ ) );
OR2_X1 _09649_ ( .A1(_02053_ ), .A2(\myifu.myicache.tag[1][1] ), .ZN(_02129_ ) );
OAI211_X1 _09650_ ( .A(_02129_ ), .B(_01955_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][1] ), .ZN(_02130_ ) );
OR2_X1 _09651_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][1] ), .ZN(_02131_ ) );
OAI211_X1 _09652_ ( .A(_02131_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02053_ ), .C2(\myifu.myicache.tag[3][1] ), .ZN(_02132_ ) );
INV_X1 _09653_ ( .A(\IF_ID_pc [6] ), .ZN(_02133_ ) );
AND3_X1 _09654_ ( .A1(_02130_ ), .A2(_02132_ ), .A3(_02133_ ), .ZN(_02134_ ) );
AOI21_X1 _09655_ ( .A(_02133_ ), .B1(_02130_ ), .B2(_02132_ ), .ZN(_02135_ ) );
OAI211_X1 _09656_ ( .A(_02127_ ), .B(_02128_ ), .C1(_02134_ ), .C2(_02135_ ), .ZN(_02136_ ) );
NOR4_X4 _09657_ ( .A1(_02082_ ), .A2(_02110_ ), .A3(_02124_ ), .A4(_02136_ ), .ZN(_02137_ ) );
AND2_X2 _09658_ ( .A1(_02052_ ), .A2(_02137_ ), .ZN(_02138_ ) );
INV_X2 _09659_ ( .A(_02138_ ), .ZN(_02139_ ) );
AND2_X4 _09660_ ( .A1(_02139_ ), .A2(\myifu.state [0] ), .ZN(_02140_ ) );
INV_X1 _09661_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_02141_ ) );
NOR2_X4 _09662_ ( .A1(_02140_ ), .A2(_02141_ ), .ZN(_02142_ ) );
NOR2_X1 _09663_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_02143_ ) );
NOR2_X4 _09664_ ( .A1(_02142_ ), .A2(_02143_ ), .ZN(_02144_ ) );
INV_X32 _09665_ ( .A(\EX_LS_flag [2] ), .ZN(_02145_ ) );
NAND4_X1 _09666_ ( .A1(_02145_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(\mylsu.state [0] ), .ZN(_02146_ ) );
INV_X1 _09667_ ( .A(EXU_valid_LSU ), .ZN(_02147_ ) );
NOR2_X1 _09668_ ( .A1(_02146_ ), .A2(_02147_ ), .ZN(_02148_ ) );
INV_X1 _09669_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_02149_ ) );
NOR2_X1 _09670_ ( .A1(_02148_ ), .A2(_02149_ ), .ZN(_02150_ ) );
NOR2_X4 _09671_ ( .A1(_02144_ ), .A2(_02150_ ), .ZN(_02151_ ) );
CLKBUF_X2 _09672_ ( .A(_02147_ ), .Z(_02152_ ) );
OR3_X1 _09673_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(_02152_ ), .ZN(_02153_ ) );
BUF_X4 _09674_ ( .A(_02148_ ), .Z(_02154_ ) );
OAI211_X1 _09675_ ( .A(_02151_ ), .B(_02153_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_02154_ ), .ZN(_02155_ ) );
BUF_X4 _09676_ ( .A(_02140_ ), .Z(_02156_ ) );
OAI221_X1 _09677_ ( .A(\IF_ID_pc [20] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02141_ ), .ZN(_02157_ ) );
AND2_X1 _09678_ ( .A1(_02155_ ), .A2(_02157_ ), .ZN(_02158_ ) );
INV_X1 _09679_ ( .A(_02158_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09680_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(_02152_ ), .ZN(_02159_ ) );
OAI211_X1 _09681_ ( .A(_02151_ ), .B(_02159_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_02148_ ), .ZN(_02160_ ) );
OAI221_X1 _09682_ ( .A(\IF_ID_pc [23] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02140_ ), .C2(_02141_ ), .ZN(_02161_ ) );
AND2_X1 _09683_ ( .A1(_02160_ ), .A2(_02161_ ), .ZN(_02162_ ) );
INV_X1 _09684_ ( .A(_02162_ ), .ZN(\io_master_araddr [23] ) );
BUF_X4 _09685_ ( .A(_02151_ ), .Z(_02163_ ) );
OR3_X1 _09686_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(_02152_ ), .ZN(_02164_ ) );
OAI211_X1 _09687_ ( .A(_02163_ ), .B(_02164_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_02154_ ), .ZN(_02165_ ) );
INV_X1 _09688_ ( .A(\IF_ID_pc [22] ), .ZN(_02166_ ) );
INV_X4 _09689_ ( .A(_02144_ ), .ZN(_02167_ ) );
OAI21_X1 _09690_ ( .A(_02165_ ), .B1(_02166_ ), .B2(_02167_ ), .ZN(\io_master_araddr [22] ) );
OR3_X1 _09691_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(_02152_ ), .ZN(_02168_ ) );
OAI211_X1 _09692_ ( .A(_02163_ ), .B(_02168_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_02154_ ), .ZN(_02169_ ) );
OAI21_X1 _09693_ ( .A(_02169_ ), .B1(_01951_ ), .B2(_02167_ ), .ZN(\io_master_araddr [21] ) );
NOR4_X2 _09694_ ( .A1(\io_master_araddr [20] ), .A2(\io_master_araddr [23] ), .A3(\io_master_araddr [22] ), .A4(\io_master_araddr [21] ), .ZN(_02170_ ) );
OR3_X1 _09695_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(_02152_ ), .ZN(_02171_ ) );
OAI211_X1 _09696_ ( .A(_02151_ ), .B(_02171_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_02154_ ), .ZN(_02172_ ) );
OAI221_X1 _09697_ ( .A(\IF_ID_pc [18] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02140_ ), .C2(_02141_ ), .ZN(_02173_ ) );
AND2_X1 _09698_ ( .A1(_02172_ ), .A2(_02173_ ), .ZN(_02174_ ) );
INV_X1 _09699_ ( .A(_02174_ ), .ZN(\io_master_araddr [18] ) );
OR3_X1 _09700_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(_02147_ ), .ZN(_02175_ ) );
OAI211_X1 _09701_ ( .A(_02151_ ), .B(_02175_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_02148_ ), .ZN(_02176_ ) );
OAI221_X1 _09702_ ( .A(\IF_ID_pc [17] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02140_ ), .C2(_02141_ ), .ZN(_02177_ ) );
AND2_X1 _09703_ ( .A1(_02176_ ), .A2(_02177_ ), .ZN(_02178_ ) );
INV_X1 _09704_ ( .A(_02178_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09705_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(_02152_ ), .ZN(_02179_ ) );
OAI211_X1 _09706_ ( .A(_02163_ ), .B(_02179_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_02154_ ), .ZN(_02180_ ) );
INV_X1 _09707_ ( .A(\IF_ID_pc [16] ), .ZN(_02181_ ) );
OAI21_X1 _09708_ ( .A(_02180_ ), .B1(_02181_ ), .B2(_02167_ ), .ZN(\io_master_araddr [16] ) );
OR3_X1 _09709_ ( .A1(_02146_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(_02152_ ), .ZN(_02182_ ) );
OAI211_X1 _09710_ ( .A(_02163_ ), .B(_02182_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_02154_ ), .ZN(_02183_ ) );
OAI21_X1 _09711_ ( .A(_02183_ ), .B1(_02064_ ), .B2(_02167_ ), .ZN(\io_master_araddr [19] ) );
NOR4_X2 _09712_ ( .A1(\io_master_araddr [18] ), .A2(\io_master_araddr [17] ), .A3(\io_master_araddr [16] ), .A4(\io_master_araddr [19] ), .ZN(_02184_ ) );
AND2_X4 _09713_ ( .A1(_02170_ ), .A2(_02184_ ), .ZN(_02185_ ) );
CLKBUF_X2 _09714_ ( .A(_02146_ ), .Z(_02186_ ) );
CLKBUF_X2 _09715_ ( .A(_02147_ ), .Z(_02187_ ) );
OR3_X1 _09716_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(_02187_ ), .ZN(_02188_ ) );
BUF_X4 _09717_ ( .A(_02154_ ), .Z(_02189_ ) );
OAI211_X1 _09718_ ( .A(_02163_ ), .B(_02188_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_02189_ ), .ZN(_02190_ ) );
BUF_X4 _09719_ ( .A(_02141_ ), .Z(_02191_ ) );
OAI221_X1 _09720_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_02192_ ) );
AND2_X1 _09721_ ( .A1(_02190_ ), .A2(_02192_ ), .ZN(_02193_ ) );
OR3_X1 _09722_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(_02187_ ), .ZN(_02194_ ) );
OAI211_X1 _09723_ ( .A(_02163_ ), .B(_02194_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_02189_ ), .ZN(_02195_ ) );
OAI221_X1 _09724_ ( .A(\IF_ID_pc [29] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_02196_ ) );
AND2_X2 _09725_ ( .A1(_02195_ ), .A2(_02196_ ), .ZN(_02197_ ) );
OR3_X1 _09726_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(_02152_ ), .ZN(_02198_ ) );
OAI211_X1 _09727_ ( .A(_02163_ ), .B(_02198_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_02154_ ), .ZN(_02199_ ) );
OAI221_X1 _09728_ ( .A(\IF_ID_pc [28] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_02200_ ) );
AND2_X2 _09729_ ( .A1(_02199_ ), .A2(_02200_ ), .ZN(_02201_ ) );
INV_X1 _09730_ ( .A(_02150_ ), .ZN(_02202_ ) );
MUX2_X1 _09731_ ( .A(\mylsu.araddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_02148_ ), .Z(_02203_ ) );
AND3_X1 _09732_ ( .A1(_02167_ ), .A2(_02202_ ), .A3(_02203_ ), .ZN(_02204_ ) );
BUF_X4 _09733_ ( .A(_02144_ ), .Z(_02205_ ) );
AOI21_X1 _09734_ ( .A(_02204_ ), .B1(\IF_ID_pc [30] ), .B2(_02205_ ), .ZN(_02206_ ) );
NAND4_X4 _09735_ ( .A1(_02193_ ), .A2(_02197_ ), .A3(_02201_ ), .A4(_02206_ ), .ZN(_02207_ ) );
OR3_X1 _09736_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(_02187_ ), .ZN(_02208_ ) );
OAI211_X1 _09737_ ( .A(_02163_ ), .B(_02208_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_02189_ ), .ZN(_02209_ ) );
OAI221_X1 _09738_ ( .A(\IF_ID_pc [24] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_02210_ ) );
AND2_X2 _09739_ ( .A1(_02209_ ), .A2(_02210_ ), .ZN(_02211_ ) );
OR3_X1 _09740_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(_02152_ ), .ZN(_02212_ ) );
OAI211_X1 _09741_ ( .A(_02163_ ), .B(_02212_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_02154_ ), .ZN(_02213_ ) );
OAI221_X1 _09742_ ( .A(\IF_ID_pc [27] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_02214_ ) );
AND2_X2 _09743_ ( .A1(_02213_ ), .A2(_02214_ ), .ZN(_02215_ ) );
OR3_X1 _09744_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(_02152_ ), .ZN(_02216_ ) );
OAI211_X1 _09745_ ( .A(_02163_ ), .B(_02216_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_02154_ ), .ZN(_02217_ ) );
OAI221_X1 _09746_ ( .A(\IF_ID_pc [26] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_02218_ ) );
AND2_X2 _09747_ ( .A1(_02217_ ), .A2(_02218_ ), .ZN(_02219_ ) );
BUF_X8 _09748_ ( .A(_02151_ ), .Z(_02220_ ) );
OR3_X1 _09749_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [25] ), .A3(_02187_ ), .ZN(_02221_ ) );
OAI211_X2 _09750_ ( .A(_02220_ ), .B(_02221_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_02189_ ), .ZN(_02222_ ) );
OAI21_X2 _09751_ ( .A(_02222_ ), .B1(_02004_ ), .B2(_02167_ ), .ZN(\io_master_araddr [25] ) );
NAND4_X4 _09752_ ( .A1(_02211_ ), .A2(_02215_ ), .A3(_02219_ ), .A4(\io_master_araddr [25] ), .ZN(_02223_ ) );
NOR2_X4 _09753_ ( .A1(_02207_ ), .A2(_02223_ ), .ZN(_02224_ ) );
AND2_X4 _09754_ ( .A1(_02185_ ), .A2(_02224_ ), .ZN(_02225_ ) );
BUF_X8 _09755_ ( .A(_02225_ ), .Z(_02226_ ) );
BUF_X2 _09756_ ( .A(_02226_ ), .Z(_02227_ ) );
BUF_X4 _09757_ ( .A(_02227_ ), .Z(_02228_ ) );
BUF_X4 _09758_ ( .A(_02228_ ), .Z(_02229_ ) );
INV_X1 _09759_ ( .A(_02229_ ), .ZN(_02230_ ) );
CLKBUF_X2 _09760_ ( .A(_02205_ ), .Z(_02231_ ) );
CLKBUF_X2 _09761_ ( .A(_02231_ ), .Z(_02232_ ) );
INV_X1 _09762_ ( .A(\EX_LS_typ [0] ), .ZN(_02233_ ) );
NOR2_X1 _09763_ ( .A1(fanout_net_6 ), .A2(\EX_LS_dest_csreg_mem [1] ), .ZN(_02234_ ) );
INV_X1 _09764_ ( .A(\EX_LS_typ [2] ), .ZN(_02235_ ) );
NOR4_X1 _09765_ ( .A1(_02234_ ), .A2(_02235_ ), .A3(\EX_LS_typ [1] ), .A4(\EX_LS_typ [3] ), .ZN(_02236_ ) );
AND2_X1 _09766_ ( .A1(fanout_net_6 ), .A2(\EX_LS_typ [1] ), .ZN(_02237_ ) );
NOR2_X1 _09767_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02238_ ) );
AND2_X1 _09768_ ( .A1(_02237_ ), .A2(_02238_ ), .ZN(_02239_ ) );
OAI21_X1 _09769_ ( .A(_02233_ ), .B1(_02236_ ), .B2(_02239_ ), .ZN(_02240_ ) );
NAND3_X1 _09770_ ( .A1(_02237_ ), .A2(_02238_ ), .A3(\EX_LS_typ [0] ), .ZN(_02241_ ) );
NAND2_X1 _09771_ ( .A1(_02240_ ), .A2(_02241_ ), .ZN(_02242_ ) );
AND2_X4 _09772_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02243_ ) );
AND2_X4 _09773_ ( .A1(_02243_ ), .A2(_02145_ ), .ZN(_02244_ ) );
INV_X1 _09774_ ( .A(\EX_LS_typ [4] ), .ZN(_02245_ ) );
AND2_X1 _09775_ ( .A1(_02244_ ), .A2(_02245_ ), .ZN(_02246_ ) );
AND2_X1 _09776_ ( .A1(_02242_ ), .A2(_02246_ ), .ZN(_02247_ ) );
OR2_X1 _09777_ ( .A1(\EX_LS_dest_csreg_mem [27] ), .A2(\EX_LS_dest_csreg_mem [25] ), .ZN(_02248_ ) );
NOR3_X1 _09778_ ( .A1(_02248_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(\EX_LS_dest_csreg_mem [24] ), .ZN(_02249_ ) );
NOR4_X1 _09779_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\EX_LS_dest_csreg_mem [29] ), .A4(\EX_LS_dest_csreg_mem [28] ), .ZN(_02250_ ) );
AND2_X1 _09780_ ( .A1(_02249_ ), .A2(_02250_ ), .ZN(_02251_ ) );
AND2_X1 _09781_ ( .A1(_02251_ ), .A2(_02244_ ), .ZN(_02252_ ) );
NOR2_X1 _09782_ ( .A1(_02247_ ), .A2(_02252_ ), .ZN(_02253_ ) );
INV_X2 _09783_ ( .A(\EX_LS_flag [1] ), .ZN(_02254_ ) );
NOR2_X1 _09784_ ( .A1(_02254_ ), .A2(\EX_LS_flag [0] ), .ZN(_02255_ ) );
AND2_X1 _09785_ ( .A1(_02255_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02256_ ) );
AND2_X1 _09786_ ( .A1(_02251_ ), .A2(_02256_ ), .ZN(_02257_ ) );
NAND3_X1 _09787_ ( .A1(_02145_ ), .A2(_02245_ ), .A3(\EX_LS_typ [0] ), .ZN(_02258_ ) );
NOR3_X1 _09788_ ( .A1(_02258_ ), .A2(_02254_ ), .A3(\EX_LS_flag [0] ), .ZN(_02259_ ) );
INV_X1 _09789_ ( .A(_02259_ ), .ZN(_02260_ ) );
INV_X1 _09790_ ( .A(_02234_ ), .ZN(_02261_ ) );
AND3_X1 _09791_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02262_ ) );
AOI22_X1 _09792_ ( .A1(_02261_ ), .A2(_02262_ ), .B1(_02237_ ), .B2(_02238_ ), .ZN(_02263_ ) );
NOR2_X1 _09793_ ( .A1(_02260_ ), .A2(_02263_ ), .ZN(_02264_ ) );
NOR2_X1 _09794_ ( .A1(_02257_ ), .A2(_02264_ ), .ZN(_02265_ ) );
AND2_X2 _09795_ ( .A1(_02253_ ), .A2(_02265_ ), .ZN(_02266_ ) );
AOI211_X1 _09796_ ( .A(_02149_ ), .B(_02232_ ), .C1(_02189_ ), .C2(_02266_ ), .ZN(_02267_ ) );
NOR2_X1 _09797_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02268_ ) );
AND3_X1 _09798_ ( .A1(_02139_ ), .A2(\myifu.state [0] ), .A3(_02268_ ), .ZN(_02269_ ) );
NOR4_X1 _09799_ ( .A1(_02142_ ), .A2(_02191_ ), .A3(_02143_ ), .A4(_02269_ ), .ZN(_02270_ ) );
OR3_X1 _09800_ ( .A1(_02230_ ), .A2(_02267_ ), .A3(_02270_ ), .ZN(_02271_ ) );
NAND2_X1 _09801_ ( .A1(_02271_ ), .A2(\myclint.rvalid ), .ZN(_02272_ ) );
AOI21_X1 _09802_ ( .A(_02232_ ), .B1(_02189_ ), .B2(_02266_ ), .ZN(_02273_ ) );
AOI211_X1 _09803_ ( .A(_02143_ ), .B(_02142_ ), .C1(\myifu.state [0] ), .C2(_02268_ ), .ZN(_02274_ ) );
OR4_X1 _09804_ ( .A1(\myclint.rvalid ), .A2(_02230_ ), .A3(_02273_ ), .A4(_02274_ ), .ZN(_02275_ ) );
AOI21_X1 _09805_ ( .A(fanout_net_2 ), .B1(_02272_ ), .B2(_02275_ ), .ZN(_00065_ ) );
INV_X1 _09806_ ( .A(\LS_WB_wdata_csreg [30] ), .ZN(_02276_ ) );
NOR2_X1 _09807_ ( .A1(_02276_ ), .A2(fanout_net_2 ), .ZN(_00066_ ) );
INV_X1 _09808_ ( .A(\LS_WB_wdata_csreg [21] ), .ZN(_02277_ ) );
NOR2_X1 _09809_ ( .A1(_02277_ ), .A2(fanout_net_2 ), .ZN(_00067_ ) );
INV_X1 _09810_ ( .A(\LS_WB_wdata_csreg [20] ), .ZN(_02278_ ) );
NOR2_X1 _09811_ ( .A1(_02278_ ), .A2(fanout_net_2 ), .ZN(_00068_ ) );
INV_X1 _09812_ ( .A(\LS_WB_wdata_csreg [19] ), .ZN(_02279_ ) );
NOR2_X1 _09813_ ( .A1(_02279_ ), .A2(fanout_net_2 ), .ZN(_00069_ ) );
INV_X1 _09814_ ( .A(\LS_WB_wdata_csreg [18] ), .ZN(_02280_ ) );
NOR2_X1 _09815_ ( .A1(_02280_ ), .A2(fanout_net_2 ), .ZN(_00070_ ) );
INV_X1 _09816_ ( .A(\LS_WB_wdata_csreg [17] ), .ZN(_02281_ ) );
NOR2_X1 _09817_ ( .A1(_02281_ ), .A2(fanout_net_2 ), .ZN(_00071_ ) );
INV_X1 _09818_ ( .A(\LS_WB_wdata_csreg [16] ), .ZN(_02282_ ) );
NOR2_X1 _09819_ ( .A1(_02282_ ), .A2(fanout_net_2 ), .ZN(_00072_ ) );
INV_X1 _09820_ ( .A(\LS_WB_wdata_csreg [15] ), .ZN(_02283_ ) );
NOR2_X1 _09821_ ( .A1(_02283_ ), .A2(fanout_net_2 ), .ZN(_00073_ ) );
INV_X1 _09822_ ( .A(\LS_WB_wdata_csreg [14] ), .ZN(_02284_ ) );
NOR2_X1 _09823_ ( .A1(_02284_ ), .A2(fanout_net_2 ), .ZN(_00074_ ) );
INV_X1 _09824_ ( .A(\LS_WB_wdata_csreg [13] ), .ZN(_02285_ ) );
NOR2_X1 _09825_ ( .A1(_02285_ ), .A2(fanout_net_2 ), .ZN(_00075_ ) );
INV_X1 _09826_ ( .A(\LS_WB_wdata_csreg [12] ), .ZN(_02286_ ) );
NOR2_X1 _09827_ ( .A1(_02286_ ), .A2(fanout_net_2 ), .ZN(_00076_ ) );
INV_X1 _09828_ ( .A(\LS_WB_wdata_csreg [29] ), .ZN(_02287_ ) );
NOR2_X1 _09829_ ( .A1(_02287_ ), .A2(fanout_net_2 ), .ZN(_00077_ ) );
INV_X1 _09830_ ( .A(\LS_WB_wdata_csreg [11] ), .ZN(_02288_ ) );
NOR2_X1 _09831_ ( .A1(_02288_ ), .A2(fanout_net_2 ), .ZN(_00078_ ) );
INV_X1 _09832_ ( .A(\LS_WB_wdata_csreg [10] ), .ZN(_02289_ ) );
NOR2_X1 _09833_ ( .A1(_02289_ ), .A2(fanout_net_2 ), .ZN(_00079_ ) );
INV_X1 _09834_ ( .A(\LS_WB_wdata_csreg [9] ), .ZN(_02290_ ) );
NOR2_X1 _09835_ ( .A1(_02290_ ), .A2(fanout_net_2 ), .ZN(_00080_ ) );
INV_X1 _09836_ ( .A(\LS_WB_wdata_csreg [8] ), .ZN(_02291_ ) );
NOR2_X1 _09837_ ( .A1(_02291_ ), .A2(fanout_net_2 ), .ZN(_00081_ ) );
INV_X1 _09838_ ( .A(\LS_WB_wdata_csreg [7] ), .ZN(_02292_ ) );
NOR2_X1 _09839_ ( .A1(_02292_ ), .A2(fanout_net_2 ), .ZN(_00082_ ) );
INV_X1 _09840_ ( .A(\LS_WB_wdata_csreg [6] ), .ZN(_02293_ ) );
NOR2_X1 _09841_ ( .A1(_02293_ ), .A2(fanout_net_2 ), .ZN(_00083_ ) );
INV_X1 _09842_ ( .A(\LS_WB_wdata_csreg [5] ), .ZN(_02294_ ) );
NOR2_X1 _09843_ ( .A1(_02294_ ), .A2(fanout_net_2 ), .ZN(_00084_ ) );
INV_X1 _09844_ ( .A(\LS_WB_wdata_csreg [4] ), .ZN(_02295_ ) );
NOR2_X1 _09845_ ( .A1(_02295_ ), .A2(fanout_net_2 ), .ZN(_00085_ ) );
INV_X1 _09846_ ( .A(\LS_WB_wdata_csreg [3] ), .ZN(_02296_ ) );
NOR2_X1 _09847_ ( .A1(_02296_ ), .A2(fanout_net_2 ), .ZN(_00086_ ) );
INV_X1 _09848_ ( .A(\LS_WB_wdata_csreg [2] ), .ZN(_02297_ ) );
NOR2_X1 _09849_ ( .A1(_02297_ ), .A2(fanout_net_2 ), .ZN(_00087_ ) );
INV_X1 _09850_ ( .A(\LS_WB_wdata_csreg [28] ), .ZN(_02298_ ) );
NOR2_X1 _09851_ ( .A1(_02298_ ), .A2(fanout_net_2 ), .ZN(_00088_ ) );
INV_X1 _09852_ ( .A(\LS_WB_wdata_csreg [1] ), .ZN(_02299_ ) );
NOR2_X1 _09853_ ( .A1(_02299_ ), .A2(fanout_net_2 ), .ZN(_00089_ ) );
INV_X1 _09854_ ( .A(\LS_WB_wdata_csreg [0] ), .ZN(_02300_ ) );
NOR2_X1 _09855_ ( .A1(_02300_ ), .A2(fanout_net_2 ), .ZN(_00090_ ) );
INV_X1 _09856_ ( .A(\LS_WB_wdata_csreg [27] ), .ZN(_02301_ ) );
NOR2_X1 _09857_ ( .A1(_02301_ ), .A2(fanout_net_3 ), .ZN(_00091_ ) );
INV_X1 _09858_ ( .A(\LS_WB_wdata_csreg [26] ), .ZN(_02302_ ) );
NOR2_X1 _09859_ ( .A1(_02302_ ), .A2(fanout_net_3 ), .ZN(_00092_ ) );
INV_X1 _09860_ ( .A(\LS_WB_wdata_csreg [25] ), .ZN(_02303_ ) );
NOR2_X1 _09861_ ( .A1(_02303_ ), .A2(fanout_net_3 ), .ZN(_00093_ ) );
INV_X1 _09862_ ( .A(\LS_WB_wdata_csreg [24] ), .ZN(_02304_ ) );
NOR2_X1 _09863_ ( .A1(_02304_ ), .A2(fanout_net_3 ), .ZN(_00094_ ) );
INV_X1 _09864_ ( .A(\LS_WB_wdata_csreg [23] ), .ZN(_02305_ ) );
NOR2_X1 _09865_ ( .A1(_02305_ ), .A2(fanout_net_3 ), .ZN(_00095_ ) );
INV_X1 _09866_ ( .A(\LS_WB_wdata_csreg [22] ), .ZN(_02306_ ) );
NOR2_X1 _09867_ ( .A1(_02306_ ), .A2(fanout_net_3 ), .ZN(_00096_ ) );
NOR3_X1 _09868_ ( .A1(_01663_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00097_ ) );
NOR3_X1 _09869_ ( .A1(_02276_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00098_ ) );
NOR3_X1 _09870_ ( .A1(_02277_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00099_ ) );
NOR3_X1 _09871_ ( .A1(_02278_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00100_ ) );
NOR3_X1 _09872_ ( .A1(_02279_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00101_ ) );
NOR3_X1 _09873_ ( .A1(_02280_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00102_ ) );
NOR3_X1 _09874_ ( .A1(_02281_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00103_ ) );
NOR3_X1 _09875_ ( .A1(_02282_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00104_ ) );
NOR3_X1 _09876_ ( .A1(_02283_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00105_ ) );
NOR3_X1 _09877_ ( .A1(_02284_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00106_ ) );
NOR3_X1 _09878_ ( .A1(_02285_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00107_ ) );
NOR3_X1 _09879_ ( .A1(_02286_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00108_ ) );
NOR3_X1 _09880_ ( .A1(_02287_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00109_ ) );
NOR3_X1 _09881_ ( .A1(_02288_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00110_ ) );
NOR3_X1 _09882_ ( .A1(_02289_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00111_ ) );
NOR3_X1 _09883_ ( .A1(_02290_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00112_ ) );
NOR3_X1 _09884_ ( .A1(_02291_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00113_ ) );
NOR3_X1 _09885_ ( .A1(_02292_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00114_ ) );
NOR3_X1 _09886_ ( .A1(_02293_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00115_ ) );
NOR3_X1 _09887_ ( .A1(_02294_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00116_ ) );
NOR3_X1 _09888_ ( .A1(_02295_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00117_ ) );
INV_X1 _09889_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02307_ ) );
NOR2_X1 _09890_ ( .A1(_02307_ ), .A2(\LS_WB_wen_csreg [3] ), .ZN(_02308_ ) );
AOI211_X1 _09891_ ( .A(fanout_net_3 ), .B(_02308_ ), .C1(_02296_ ), .C2(_02307_ ), .ZN(_00118_ ) );
NOR2_X1 _09892_ ( .A1(_02307_ ), .A2(\LS_WB_wen_csreg [2] ), .ZN(_02309_ ) );
AOI211_X1 _09893_ ( .A(fanout_net_3 ), .B(_02309_ ), .C1(_02297_ ), .C2(_02307_ ), .ZN(_00119_ ) );
NOR3_X1 _09894_ ( .A1(_02298_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00120_ ) );
NOR2_X1 _09895_ ( .A1(_02307_ ), .A2(\LS_WB_wen_csreg [1] ), .ZN(_02310_ ) );
AOI211_X1 _09896_ ( .A(fanout_net_4 ), .B(_02310_ ), .C1(_02299_ ), .C2(_02307_ ), .ZN(_00121_ ) );
NOR2_X1 _09897_ ( .A1(_02307_ ), .A2(\LS_WB_wen_csreg [0] ), .ZN(_02311_ ) );
AOI211_X1 _09898_ ( .A(fanout_net_4 ), .B(_02311_ ), .C1(_02300_ ), .C2(_02307_ ), .ZN(_00122_ ) );
NOR3_X1 _09899_ ( .A1(_02301_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00123_ ) );
NOR3_X1 _09900_ ( .A1(_02302_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00124_ ) );
NOR3_X1 _09901_ ( .A1(_02303_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00125_ ) );
NOR3_X1 _09902_ ( .A1(_02304_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00126_ ) );
NOR3_X1 _09903_ ( .A1(_02305_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00127_ ) );
NOR3_X1 _09904_ ( .A1(_02306_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00128_ ) );
AND3_X1 _09905_ ( .A1(_01813_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00129_ ) );
NOR2_X1 _09906_ ( .A1(\myec.state [1] ), .A2(\myec.state [0] ), .ZN(_02312_ ) );
AND2_X1 _09907_ ( .A1(_02312_ ), .A2(_01664_ ), .ZN(_02313_ ) );
INV_X1 _09908_ ( .A(_02313_ ), .ZN(_02314_ ) );
INV_X1 _09909_ ( .A(_02266_ ), .ZN(_02315_ ) );
INV_X1 _09910_ ( .A(exception_quest_IDU ), .ZN(_02316_ ) );
OR2_X1 _09911_ ( .A1(\myexu.pc_jump [27] ), .A2(\myexu.pc_jump [26] ), .ZN(_02317_ ) );
OR3_X1 _09912_ ( .A1(_02317_ ), .A2(\myexu.pc_jump [25] ), .A3(\myexu.pc_jump [24] ), .ZN(_02318_ ) );
OR4_X1 _09913_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02319_ ) );
NOR2_X1 _09914_ ( .A1(_02318_ ), .A2(_02319_ ), .ZN(_02320_ ) );
NOR2_X1 _09915_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02321_ ) );
INV_X1 _09916_ ( .A(_02321_ ), .ZN(_02322_ ) );
NOR2_X1 _09917_ ( .A1(_02320_ ), .A2(_02322_ ), .ZN(_02323_ ) );
AOI211_X1 _09918_ ( .A(_02314_ ), .B(_02315_ ), .C1(_02316_ ), .C2(_02323_ ), .ZN(_00130_ ) );
AOI21_X1 _09919_ ( .A(_02314_ ), .B1(_02266_ ), .B2(exception_quest_IDU ), .ZN(_00131_ ) );
INV_X1 _09920_ ( .A(fanout_net_29 ), .ZN(_02324_ ) );
BUF_X4 _09921_ ( .A(_02324_ ), .Z(_02325_ ) );
BUF_X4 _09922_ ( .A(_02325_ ), .Z(_02326_ ) );
BUF_X4 _09923_ ( .A(_02326_ ), .Z(_02327_ ) );
OR2_X1 _09924_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02328_ ) );
INV_X32 _09925_ ( .A(fanout_net_26 ), .ZN(_02329_ ) );
BUF_X4 _09926_ ( .A(_02329_ ), .Z(_02330_ ) );
BUF_X4 _09927_ ( .A(_02330_ ), .Z(_02331_ ) );
BUF_X8 _09928_ ( .A(_02331_ ), .Z(_02332_ ) );
BUF_X4 _09929_ ( .A(_02332_ ), .Z(_02333_ ) );
BUF_X4 _09930_ ( .A(_02333_ ), .Z(_02334_ ) );
BUF_X4 _09931_ ( .A(_02334_ ), .Z(_02335_ ) );
INV_X32 _09932_ ( .A(fanout_net_18 ), .ZN(_02336_ ) );
BUF_X4 _09933_ ( .A(_02336_ ), .Z(_02337_ ) );
BUF_X4 _09934_ ( .A(_02337_ ), .Z(_02338_ ) );
BUF_X8 _09935_ ( .A(_02338_ ), .Z(_02339_ ) );
BUF_X4 _09936_ ( .A(_02339_ ), .Z(_02340_ ) );
BUF_X4 _09937_ ( .A(_02340_ ), .Z(_02341_ ) );
BUF_X4 _09938_ ( .A(_02341_ ), .Z(_02342_ ) );
OAI211_X1 _09939_ ( .A(_02328_ ), .B(_02335_ ), .C1(_02342_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02343_ ) );
OR2_X1 _09940_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02344_ ) );
OAI211_X1 _09941_ ( .A(_02344_ ), .B(fanout_net_26 ), .C1(_02342_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02345_ ) );
INV_X1 _09942_ ( .A(fanout_net_28 ), .ZN(_02346_ ) );
BUF_X4 _09943_ ( .A(_02346_ ), .Z(_02347_ ) );
BUF_X4 _09944_ ( .A(_02347_ ), .Z(_02348_ ) );
BUF_X4 _09945_ ( .A(_02348_ ), .Z(_02349_ ) );
BUF_X4 _09946_ ( .A(_02349_ ), .Z(_02350_ ) );
BUF_X4 _09947_ ( .A(_02350_ ), .Z(_02351_ ) );
NAND3_X1 _09948_ ( .A1(_02343_ ), .A2(_02345_ ), .A3(_02351_ ), .ZN(_02352_ ) );
MUX2_X1 _09949_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02353_ ) );
MUX2_X1 _09950_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02354_ ) );
MUX2_X1 _09951_ ( .A(_02353_ ), .B(_02354_ ), .S(_02334_ ), .Z(_02355_ ) );
BUF_X4 _09952_ ( .A(_02350_ ), .Z(_02356_ ) );
OAI211_X1 _09953_ ( .A(_02327_ ), .B(_02352_ ), .C1(_02355_ ), .C2(_02356_ ), .ZN(_02357_ ) );
INV_X1 _09954_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02358_ ) );
INV_X1 _09955_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02359_ ) );
MUX2_X1 _09956_ ( .A(_02358_ ), .B(_02359_ ), .S(fanout_net_18 ), .Z(_02360_ ) );
AND2_X1 _09957_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02361_ ) );
BUF_X4 _09958_ ( .A(_02337_ ), .Z(_02362_ ) );
BUF_X4 _09959_ ( .A(_02362_ ), .Z(_02363_ ) );
BUF_X4 _09960_ ( .A(_02363_ ), .Z(_02364_ ) );
AOI21_X1 _09961_ ( .A(_02361_ ), .B1(_02364_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02365_ ) );
MUX2_X1 _09962_ ( .A(_02360_ ), .B(_02365_ ), .S(_02334_ ), .Z(_02366_ ) );
AND2_X1 _09963_ ( .A1(_02363_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02367_ ) );
AOI21_X1 _09964_ ( .A(_02367_ ), .B1(fanout_net_18 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02368_ ) );
NOR2_X1 _09965_ ( .A1(_02368_ ), .A2(fanout_net_26 ), .ZN(_02369_ ) );
MUX2_X1 _09966_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02370_ ) );
AOI21_X1 _09967_ ( .A(_02369_ ), .B1(fanout_net_26 ), .B2(_02370_ ), .ZN(_02371_ ) );
MUX2_X1 _09968_ ( .A(_02366_ ), .B(_02371_ ), .S(fanout_net_28 ), .Z(_02372_ ) );
OAI21_X1 _09969_ ( .A(_02357_ ), .B1(_02372_ ), .B2(_02327_ ), .ZN(_02373_ ) );
AND2_X2 _09970_ ( .A1(_02254_ ), .A2(\EX_LS_flag [0] ), .ZN(_02374_ ) );
AOI21_X4 _09971_ ( .A(_02244_ ), .B1(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .B2(_02374_ ), .ZN(_02375_ ) );
INV_X4 _09972_ ( .A(_02375_ ), .ZN(_02376_ ) );
NOR2_X1 _09973_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02377_ ) );
NOR3_X4 _09974_ ( .A1(_02243_ ), .A2(_02377_ ), .A3(_02145_ ), .ZN(_02378_ ) );
NOR2_X4 _09975_ ( .A1(_02376_ ), .A2(_02378_ ), .ZN(_02379_ ) );
XOR2_X2 _09976_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .Z(_02380_ ) );
INV_X16 _09977_ ( .A(\EX_LS_dest_reg [3] ), .ZN(_02381_ ) );
OAI21_X1 _09978_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02381_ ), .B2(\ID_EX_rs1 [3] ), .ZN(_02382_ ) );
XNOR2_X1 _09979_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .ZN(_02383_ ) );
NAND2_X1 _09980_ ( .A1(_02381_ ), .A2(\ID_EX_rs1 [3] ), .ZN(_02384_ ) );
INV_X16 _09981_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02385_ ) );
OR2_X1 _09982_ ( .A1(_02385_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02386_ ) );
NAND3_X1 _09983_ ( .A1(_02383_ ), .A2(_02384_ ), .A3(_02386_ ), .ZN(_02387_ ) );
OR4_X4 _09984_ ( .A1(_02379_ ), .A2(_02380_ ), .A3(_02382_ ), .A4(_02387_ ), .ZN(_02388_ ) );
BUF_X4 _09985_ ( .A(_02388_ ), .Z(_02389_ ) );
BUF_X2 _09986_ ( .A(_02389_ ), .Z(_02390_ ) );
XNOR2_X2 _09987_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02391_ ) );
NAND2_X1 _09988_ ( .A1(_02385_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02392_ ) );
OR3_X4 _09989_ ( .A1(\EX_LS_dest_reg [2] ), .A2(\EX_LS_dest_reg [1] ), .A3(\EX_LS_dest_reg [0] ), .ZN(_02393_ ) );
OR2_X4 _09990_ ( .A1(\EX_LS_dest_reg [4] ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02394_ ) );
OAI211_X1 _09991_ ( .A(_02391_ ), .B(_02392_ ), .C1(_02393_ ), .C2(_02394_ ), .ZN(_02395_ ) );
CLKBUF_X2 _09992_ ( .A(_02395_ ), .Z(_02396_ ) );
BUF_X2 _09993_ ( .A(_02396_ ), .Z(_02397_ ) );
NOR2_X1 _09994_ ( .A1(_02390_ ), .A2(_02397_ ), .ZN(_02398_ ) );
OR2_X2 _09995_ ( .A1(_02373_ ), .A2(_02398_ ), .ZN(_02399_ ) );
OR3_X2 _09996_ ( .A1(_02390_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02397_ ), .ZN(_02400_ ) );
AND2_X2 _09997_ ( .A1(_02399_ ), .A2(_02400_ ), .ZN(_02401_ ) );
INV_X1 _09998_ ( .A(\ID_EX_imm [30] ), .ZN(_02402_ ) );
XNOR2_X1 _09999_ ( .A(_02401_ ), .B(_02402_ ), .ZN(_02403_ ) );
OR2_X1 _10000_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02404_ ) );
BUF_X4 _10001_ ( .A(_02334_ ), .Z(_02405_ ) );
BUF_X4 _10002_ ( .A(_02341_ ), .Z(_02406_ ) );
OAI211_X1 _10003_ ( .A(_02404_ ), .B(_02405_ ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02407_ ) );
OR2_X1 _10004_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02408_ ) );
OAI211_X1 _10005_ ( .A(_02408_ ), .B(fanout_net_26 ), .C1(_02342_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02409_ ) );
NAND3_X1 _10006_ ( .A1(_02407_ ), .A2(_02409_ ), .A3(fanout_net_28 ), .ZN(_02410_ ) );
MUX2_X1 _10007_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02411_ ) );
MUX2_X1 _10008_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02412_ ) );
MUX2_X1 _10009_ ( .A(_02411_ ), .B(_02412_ ), .S(_02335_ ), .Z(_02413_ ) );
OAI211_X1 _10010_ ( .A(_02327_ ), .B(_02410_ ), .C1(_02413_ ), .C2(fanout_net_28 ), .ZN(_02414_ ) );
MUX2_X1 _10011_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02415_ ) );
AND2_X1 _10012_ ( .A1(_02415_ ), .A2(fanout_net_26 ), .ZN(_02416_ ) );
MUX2_X1 _10013_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02417_ ) );
AOI211_X1 _10014_ ( .A(fanout_net_28 ), .B(_02416_ ), .C1(_02405_ ), .C2(_02417_ ), .ZN(_02418_ ) );
MUX2_X1 _10015_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02419_ ) );
MUX2_X1 _10016_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02420_ ) );
MUX2_X1 _10017_ ( .A(_02419_ ), .B(_02420_ ), .S(fanout_net_26 ), .Z(_02421_ ) );
OAI21_X1 _10018_ ( .A(fanout_net_29 ), .B1(_02421_ ), .B2(_02351_ ), .ZN(_02422_ ) );
OAI221_X1 _10019_ ( .A(_02414_ ), .B1(_02418_ ), .B2(_02422_ ), .C1(_02390_ ), .C2(_02397_ ), .ZN(_02423_ ) );
OR3_X2 _10020_ ( .A1(_02390_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02397_ ), .ZN(_02424_ ) );
NAND2_X1 _10021_ ( .A1(_02423_ ), .A2(_02424_ ), .ZN(_02425_ ) );
INV_X1 _10022_ ( .A(\ID_EX_imm [29] ), .ZN(_02426_ ) );
XNOR2_X1 _10023_ ( .A(_02425_ ), .B(_02426_ ), .ZN(_02427_ ) );
OR3_X1 _10024_ ( .A1(_02389_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02396_ ), .ZN(_02428_ ) );
OR2_X1 _10025_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02429_ ) );
OAI211_X1 _10026_ ( .A(_02429_ ), .B(_02335_ ), .C1(_02342_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02430_ ) );
OR2_X1 _10027_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02431_ ) );
OAI211_X1 _10028_ ( .A(_02431_ ), .B(fanout_net_26 ), .C1(_02342_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02432_ ) );
NAND3_X1 _10029_ ( .A1(_02430_ ), .A2(_02432_ ), .A3(_02351_ ), .ZN(_02433_ ) );
MUX2_X1 _10030_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02434_ ) );
MUX2_X1 _10031_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02435_ ) );
MUX2_X1 _10032_ ( .A(_02434_ ), .B(_02435_ ), .S(_02334_ ), .Z(_02436_ ) );
OAI211_X1 _10033_ ( .A(_02327_ ), .B(_02433_ ), .C1(_02436_ ), .C2(_02356_ ), .ZN(_02437_ ) );
OR2_X1 _10034_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02438_ ) );
OAI211_X1 _10035_ ( .A(_02438_ ), .B(_02334_ ), .C1(_02341_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02439_ ) );
NOR2_X1 _10036_ ( .A1(_02342_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02440_ ) );
OAI21_X1 _10037_ ( .A(fanout_net_26 ), .B1(fanout_net_18 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02441_ ) );
OAI211_X1 _10038_ ( .A(_02439_ ), .B(fanout_net_28 ), .C1(_02440_ ), .C2(_02441_ ), .ZN(_02442_ ) );
MUX2_X1 _10039_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02443_ ) );
MUX2_X1 _10040_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02444_ ) );
MUX2_X1 _10041_ ( .A(_02443_ ), .B(_02444_ ), .S(fanout_net_26 ), .Z(_02445_ ) );
OAI211_X1 _10042_ ( .A(fanout_net_29 ), .B(_02442_ ), .C1(_02445_ ), .C2(fanout_net_28 ), .ZN(_02446_ ) );
OAI211_X1 _10043_ ( .A(_02437_ ), .B(_02446_ ), .C1(_02390_ ), .C2(_02397_ ), .ZN(_02447_ ) );
NAND2_X1 _10044_ ( .A1(_02428_ ), .A2(_02447_ ), .ZN(_02448_ ) );
XNOR2_X1 _10045_ ( .A(_02448_ ), .B(\ID_EX_imm [28] ), .ZN(_02449_ ) );
INV_X1 _10046_ ( .A(_02449_ ), .ZN(_02450_ ) );
OR2_X1 _10047_ ( .A1(_02381_ ), .A2(\ID_EX_rs1 [3] ), .ZN(_02451_ ) );
NAND3_X1 _10048_ ( .A1(_02383_ ), .A2(_02451_ ), .A3(_02384_ ), .ZN(_02452_ ) );
NAND3_X2 _10049_ ( .A1(_02391_ ), .A2(_02392_ ), .A3(_02386_ ), .ZN(_02453_ ) );
NOR2_X4 _10050_ ( .A1(_02393_ ), .A2(_02394_ ), .ZN(_02454_ ) );
NOR4_X4 _10051_ ( .A1(_02452_ ), .A2(_02453_ ), .A3(_02454_ ), .A4(_02380_ ), .ZN(_02455_ ) );
OAI21_X4 _10052_ ( .A(_02455_ ), .B1(_02378_ ), .B2(_02376_ ), .ZN(_02456_ ) );
INV_X1 _10053_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .ZN(_02457_ ) );
NOR2_X4 _10054_ ( .A1(_02456_ ), .A2(_02457_ ), .ZN(_02458_ ) );
BUF_X8 _10055_ ( .A(_02458_ ), .Z(_02459_ ) );
BUF_X16 _10056_ ( .A(_02459_ ), .Z(_02460_ ) );
NAND2_X1 _10057_ ( .A1(_02460_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .ZN(_02461_ ) );
OR2_X1 _10058_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02462_ ) );
OAI211_X1 _10059_ ( .A(_02462_ ), .B(_02334_ ), .C1(_02341_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02463_ ) );
INV_X1 _10060_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02464_ ) );
INV_X1 _10061_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02465_ ) );
MUX2_X1 _10062_ ( .A(_02464_ ), .B(_02465_ ), .S(fanout_net_18 ), .Z(_02466_ ) );
OAI211_X1 _10063_ ( .A(_02463_ ), .B(_02351_ ), .C1(_02466_ ), .C2(_02405_ ), .ZN(_02467_ ) );
MUX2_X1 _10064_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02468_ ) );
MUX2_X1 _10065_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02469_ ) );
MUX2_X1 _10066_ ( .A(_02468_ ), .B(_02469_ ), .S(_02334_ ), .Z(_02470_ ) );
OAI211_X1 _10067_ ( .A(fanout_net_29 ), .B(_02467_ ), .C1(_02470_ ), .C2(_02351_ ), .ZN(_02471_ ) );
OR2_X1 _10068_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02472_ ) );
OAI211_X1 _10069_ ( .A(_02472_ ), .B(_02335_ ), .C1(_02341_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02473_ ) );
OR2_X1 _10070_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02474_ ) );
OAI211_X1 _10071_ ( .A(_02474_ ), .B(fanout_net_26 ), .C1(_02341_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02475_ ) );
NAND3_X1 _10072_ ( .A1(_02473_ ), .A2(_02475_ ), .A3(_02351_ ), .ZN(_02476_ ) );
MUX2_X1 _10073_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02477_ ) );
MUX2_X1 _10074_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02478_ ) );
MUX2_X1 _10075_ ( .A(_02477_ ), .B(_02478_ ), .S(_02334_ ), .Z(_02479_ ) );
OAI211_X1 _10076_ ( .A(_02327_ ), .B(_02476_ ), .C1(_02479_ ), .C2(_02351_ ), .ZN(_02480_ ) );
NAND2_X1 _10077_ ( .A1(_02471_ ), .A2(_02480_ ), .ZN(_02481_ ) );
BUF_X16 _10078_ ( .A(_02456_ ), .Z(_02482_ ) );
BUF_X16 _10079_ ( .A(_02482_ ), .Z(_02483_ ) );
BUF_X4 _10080_ ( .A(_02457_ ), .Z(_02484_ ) );
BUF_X4 _10081_ ( .A(_02484_ ), .Z(_02485_ ) );
OAI21_X1 _10082_ ( .A(_02481_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02486_ ) );
AND2_X2 _10083_ ( .A1(_02461_ ), .A2(_02486_ ), .ZN(_02487_ ) );
INV_X1 _10084_ ( .A(\ID_EX_imm [27] ), .ZN(_02488_ ) );
XNOR2_X1 _10085_ ( .A(_02487_ ), .B(_02488_ ), .ZN(_02489_ ) );
OR3_X1 _10086_ ( .A1(_02390_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02396_ ), .ZN(_02490_ ) );
OR2_X1 _10087_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02491_ ) );
OAI211_X1 _10088_ ( .A(_02491_ ), .B(_02405_ ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02492_ ) );
OR2_X1 _10089_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02493_ ) );
OAI211_X1 _10090_ ( .A(_02493_ ), .B(fanout_net_26 ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02494_ ) );
NAND3_X1 _10091_ ( .A1(_02492_ ), .A2(_02494_ ), .A3(_02351_ ), .ZN(_02495_ ) );
MUX2_X1 _10092_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02496_ ) );
MUX2_X1 _10093_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02497_ ) );
MUX2_X1 _10094_ ( .A(_02496_ ), .B(_02497_ ), .S(_02335_ ), .Z(_02498_ ) );
OAI211_X1 _10095_ ( .A(_02327_ ), .B(_02495_ ), .C1(_02498_ ), .C2(_02356_ ), .ZN(_02499_ ) );
OR2_X1 _10096_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02500_ ) );
OAI211_X1 _10097_ ( .A(_02500_ ), .B(_02335_ ), .C1(_02342_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02501_ ) );
NOR2_X1 _10098_ ( .A1(_02406_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02502_ ) );
OAI21_X1 _10099_ ( .A(fanout_net_26 ), .B1(fanout_net_19 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02503_ ) );
OAI211_X1 _10100_ ( .A(_02501_ ), .B(fanout_net_28 ), .C1(_02502_ ), .C2(_02503_ ), .ZN(_02504_ ) );
MUX2_X1 _10101_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02505_ ) );
MUX2_X1 _10102_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02506_ ) );
MUX2_X1 _10103_ ( .A(_02505_ ), .B(_02506_ ), .S(fanout_net_26 ), .Z(_02507_ ) );
OAI211_X1 _10104_ ( .A(fanout_net_29 ), .B(_02504_ ), .C1(_02507_ ), .C2(fanout_net_28 ), .ZN(_02508_ ) );
OAI211_X1 _10105_ ( .A(_02499_ ), .B(_02508_ ), .C1(_02390_ ), .C2(_02397_ ), .ZN(_02509_ ) );
NAND2_X1 _10106_ ( .A1(_02490_ ), .A2(_02509_ ), .ZN(_02510_ ) );
INV_X1 _10107_ ( .A(\ID_EX_imm [24] ), .ZN(_02511_ ) );
XNOR2_X1 _10108_ ( .A(_02510_ ), .B(_02511_ ), .ZN(_02512_ ) );
INV_X1 _10109_ ( .A(_02512_ ), .ZN(_02513_ ) );
OR3_X1 _10110_ ( .A1(_02388_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02395_ ), .ZN(_02514_ ) );
OR2_X1 _10111_ ( .A1(_02339_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02515_ ) );
OAI211_X1 _10112_ ( .A(_02515_ ), .B(_02333_ ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02516_ ) );
BUF_X4 _10113_ ( .A(_02349_ ), .Z(_02517_ ) );
OR2_X1 _10114_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02518_ ) );
OAI211_X1 _10115_ ( .A(_02518_ ), .B(fanout_net_26 ), .C1(_02340_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02519_ ) );
NAND3_X1 _10116_ ( .A1(_02516_ ), .A2(_02517_ ), .A3(_02519_ ), .ZN(_02520_ ) );
MUX2_X1 _10117_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02521_ ) );
MUX2_X1 _10118_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02522_ ) );
MUX2_X1 _10119_ ( .A(_02521_ ), .B(_02522_ ), .S(_02333_ ), .Z(_02523_ ) );
OAI211_X1 _10120_ ( .A(fanout_net_29 ), .B(_02520_ ), .C1(_02523_ ), .C2(_02517_ ), .ZN(_02524_ ) );
OR2_X1 _10121_ ( .A1(_02339_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02525_ ) );
OAI211_X1 _10122_ ( .A(_02525_ ), .B(_02333_ ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02526_ ) );
OR2_X1 _10123_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02527_ ) );
OAI211_X1 _10124_ ( .A(_02527_ ), .B(fanout_net_26 ), .C1(_02340_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02528_ ) );
NAND3_X1 _10125_ ( .A1(_02526_ ), .A2(_02517_ ), .A3(_02528_ ), .ZN(_02529_ ) );
MUX2_X1 _10126_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02530_ ) );
MUX2_X1 _10127_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02531_ ) );
MUX2_X1 _10128_ ( .A(_02530_ ), .B(_02531_ ), .S(_02333_ ), .Z(_02532_ ) );
OAI211_X1 _10129_ ( .A(_02326_ ), .B(_02529_ ), .C1(_02532_ ), .C2(_02517_ ), .ZN(_02533_ ) );
OAI211_X4 _10130_ ( .A(_02524_ ), .B(_02533_ ), .C1(_02389_ ), .C2(_02396_ ), .ZN(_02534_ ) );
NAND2_X2 _10131_ ( .A1(_02514_ ), .A2(_02534_ ), .ZN(_02535_ ) );
INV_X1 _10132_ ( .A(\ID_EX_imm [22] ), .ZN(_02536_ ) );
XNOR2_X1 _10133_ ( .A(_02535_ ), .B(_02536_ ), .ZN(_02537_ ) );
NAND2_X1 _10134_ ( .A1(_02460_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02538_ ) );
OR2_X1 _10135_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02539_ ) );
OAI211_X1 _10136_ ( .A(_02539_ ), .B(_02333_ ), .C1(_02340_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02540_ ) );
OR2_X1 _10137_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02541_ ) );
OAI211_X1 _10138_ ( .A(_02541_ ), .B(fanout_net_26 ), .C1(_02340_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02542_ ) );
NAND3_X1 _10139_ ( .A1(_02540_ ), .A2(_02542_ ), .A3(_02349_ ), .ZN(_02543_ ) );
MUX2_X1 _10140_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02544_ ) );
MUX2_X1 _10141_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02545_ ) );
BUF_X4 _10142_ ( .A(_02330_ ), .Z(_02546_ ) );
BUF_X4 _10143_ ( .A(_02546_ ), .Z(_02547_ ) );
MUX2_X1 _10144_ ( .A(_02544_ ), .B(_02545_ ), .S(_02547_ ), .Z(_02548_ ) );
OAI211_X1 _10145_ ( .A(_02326_ ), .B(_02543_ ), .C1(_02548_ ), .C2(_02517_ ), .ZN(_02549_ ) );
OR2_X1 _10146_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02550_ ) );
OAI211_X1 _10147_ ( .A(_02550_ ), .B(fanout_net_26 ), .C1(_02340_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02551_ ) );
OR2_X1 _10148_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02552_ ) );
OAI211_X1 _10149_ ( .A(_02552_ ), .B(_02333_ ), .C1(_02340_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02553_ ) );
NAND3_X1 _10150_ ( .A1(_02551_ ), .A2(_02553_ ), .A3(fanout_net_28 ), .ZN(_02554_ ) );
MUX2_X1 _10151_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02555_ ) );
MUX2_X1 _10152_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02556_ ) );
MUX2_X1 _10153_ ( .A(_02555_ ), .B(_02556_ ), .S(fanout_net_26 ), .Z(_02557_ ) );
OAI211_X1 _10154_ ( .A(fanout_net_29 ), .B(_02554_ ), .C1(_02557_ ), .C2(fanout_net_28 ), .ZN(_02558_ ) );
NAND2_X1 _10155_ ( .A1(_02549_ ), .A2(_02558_ ), .ZN(_02559_ ) );
OAI21_X2 _10156_ ( .A(_02559_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02560_ ) );
AND2_X4 _10157_ ( .A1(_02538_ ), .A2(_02560_ ), .ZN(_02561_ ) );
INV_X1 _10158_ ( .A(\ID_EX_imm [23] ), .ZN(_02562_ ) );
XNOR2_X1 _10159_ ( .A(_02561_ ), .B(_02562_ ), .ZN(_02563_ ) );
AND2_X1 _10160_ ( .A1(_02537_ ), .A2(_02563_ ), .ZN(_02564_ ) );
NAND2_X1 _10161_ ( .A1(_02460_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02565_ ) );
OR2_X1 _10162_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02566_ ) );
OAI211_X1 _10163_ ( .A(_02566_ ), .B(_02547_ ), .C1(_02363_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02567_ ) );
OR2_X1 _10164_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02568_ ) );
OAI211_X1 _10165_ ( .A(_02568_ ), .B(fanout_net_26 ), .C1(_02363_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02569_ ) );
NAND3_X1 _10166_ ( .A1(_02567_ ), .A2(_02569_ ), .A3(_02349_ ), .ZN(_02570_ ) );
MUX2_X1 _10167_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02571_ ) );
MUX2_X1 _10168_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02572_ ) );
MUX2_X1 _10169_ ( .A(_02571_ ), .B(_02572_ ), .S(_02332_ ), .Z(_02573_ ) );
OAI211_X1 _10170_ ( .A(_02326_ ), .B(_02570_ ), .C1(_02573_ ), .C2(_02349_ ), .ZN(_02574_ ) );
OR2_X1 _10171_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02575_ ) );
OAI211_X1 _10172_ ( .A(_02575_ ), .B(fanout_net_26 ), .C1(_02363_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02576_ ) );
OR2_X1 _10173_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02577_ ) );
OAI211_X1 _10174_ ( .A(_02577_ ), .B(_02547_ ), .C1(_02339_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02578_ ) );
NAND3_X1 _10175_ ( .A1(_02576_ ), .A2(_02578_ ), .A3(fanout_net_28 ), .ZN(_02579_ ) );
MUX2_X1 _10176_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02580_ ) );
MUX2_X1 _10177_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02581_ ) );
MUX2_X1 _10178_ ( .A(_02580_ ), .B(_02581_ ), .S(fanout_net_26 ), .Z(_02582_ ) );
OAI211_X1 _10179_ ( .A(fanout_net_29 ), .B(_02579_ ), .C1(_02582_ ), .C2(fanout_net_28 ), .ZN(_02583_ ) );
NAND2_X1 _10180_ ( .A1(_02574_ ), .A2(_02583_ ), .ZN(_02584_ ) );
OAI21_X4 _10181_ ( .A(_02584_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02585_ ) );
AND3_X1 _10182_ ( .A1(_02565_ ), .A2(\ID_EX_imm [21] ), .A3(_02585_ ), .ZN(_02586_ ) );
AOI21_X1 _10183_ ( .A(\ID_EX_imm [21] ), .B1(_02565_ ), .B2(_02585_ ), .ZN(_02587_ ) );
NOR2_X1 _10184_ ( .A1(_02586_ ), .A2(_02587_ ), .ZN(_02588_ ) );
OR3_X4 _10185_ ( .A1(_02389_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02396_ ), .ZN(_02589_ ) );
OR2_X1 _10186_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02590_ ) );
BUF_X4 _10187_ ( .A(_02547_ ), .Z(_02591_ ) );
OAI211_X1 _10188_ ( .A(_02590_ ), .B(_02591_ ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02592_ ) );
OR2_X1 _10189_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02593_ ) );
OAI211_X1 _10190_ ( .A(_02593_ ), .B(fanout_net_26 ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02594_ ) );
NAND3_X1 _10191_ ( .A1(_02592_ ), .A2(_02594_ ), .A3(_02517_ ), .ZN(_02595_ ) );
MUX2_X1 _10192_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02596_ ) );
MUX2_X1 _10193_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02597_ ) );
MUX2_X1 _10194_ ( .A(_02596_ ), .B(_02597_ ), .S(_02333_ ), .Z(_02598_ ) );
OAI211_X1 _10195_ ( .A(_02326_ ), .B(_02595_ ), .C1(_02598_ ), .C2(_02350_ ), .ZN(_02599_ ) );
OR2_X1 _10196_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02600_ ) );
OAI211_X1 _10197_ ( .A(_02600_ ), .B(fanout_net_26 ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02601_ ) );
OR2_X1 _10198_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02602_ ) );
OAI211_X1 _10199_ ( .A(_02602_ ), .B(_02591_ ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02603_ ) );
NAND3_X1 _10200_ ( .A1(_02601_ ), .A2(_02603_ ), .A3(fanout_net_28 ), .ZN(_02604_ ) );
MUX2_X1 _10201_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02605_ ) );
MUX2_X1 _10202_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02606_ ) );
MUX2_X1 _10203_ ( .A(_02605_ ), .B(_02606_ ), .S(fanout_net_26 ), .Z(_02607_ ) );
OAI211_X1 _10204_ ( .A(fanout_net_29 ), .B(_02604_ ), .C1(_02607_ ), .C2(fanout_net_28 ), .ZN(_02608_ ) );
OAI211_X1 _10205_ ( .A(_02599_ ), .B(_02608_ ), .C1(_02389_ ), .C2(_02396_ ), .ZN(_02609_ ) );
NAND2_X4 _10206_ ( .A1(_02589_ ), .A2(_02609_ ), .ZN(_02610_ ) );
XOR2_X1 _10207_ ( .A(_02610_ ), .B(\ID_EX_imm [20] ), .Z(_02611_ ) );
AND3_X1 _10208_ ( .A1(_02564_ ), .A2(_02588_ ), .A3(_02611_ ), .ZN(_02612_ ) );
INV_X1 _10209_ ( .A(_02612_ ), .ZN(_02613_ ) );
OR3_X2 _10210_ ( .A1(_02389_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02396_ ), .ZN(_02614_ ) );
OR2_X1 _10211_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02615_ ) );
OAI211_X1 _10212_ ( .A(_02615_ ), .B(_02591_ ), .C1(_02341_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02616_ ) );
OR2_X1 _10213_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02617_ ) );
OAI211_X1 _10214_ ( .A(_02617_ ), .B(fanout_net_26 ), .C1(_02341_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02618_ ) );
NAND3_X1 _10215_ ( .A1(_02616_ ), .A2(_02618_ ), .A3(_02350_ ), .ZN(_02619_ ) );
MUX2_X1 _10216_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02620_ ) );
MUX2_X1 _10217_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02621_ ) );
MUX2_X1 _10218_ ( .A(_02620_ ), .B(_02621_ ), .S(_02591_ ), .Z(_02622_ ) );
OAI211_X1 _10219_ ( .A(fanout_net_29 ), .B(_02619_ ), .C1(_02622_ ), .C2(_02350_ ), .ZN(_02623_ ) );
OR2_X1 _10220_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02624_ ) );
OAI211_X1 _10221_ ( .A(_02624_ ), .B(_02591_ ), .C1(_02341_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02625_ ) );
OR2_X1 _10222_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02626_ ) );
OAI211_X1 _10223_ ( .A(_02626_ ), .B(fanout_net_26 ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02627_ ) );
NAND3_X1 _10224_ ( .A1(_02625_ ), .A2(_02627_ ), .A3(_02350_ ), .ZN(_02628_ ) );
MUX2_X1 _10225_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02629_ ) );
MUX2_X1 _10226_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02630_ ) );
MUX2_X1 _10227_ ( .A(_02629_ ), .B(_02630_ ), .S(_02591_ ), .Z(_02631_ ) );
OAI211_X1 _10228_ ( .A(_02327_ ), .B(_02628_ ), .C1(_02631_ ), .C2(_02350_ ), .ZN(_02632_ ) );
OAI211_X1 _10229_ ( .A(_02623_ ), .B(_02632_ ), .C1(_02389_ ), .C2(_02396_ ), .ZN(_02633_ ) );
NAND2_X4 _10230_ ( .A1(_02614_ ), .A2(_02633_ ), .ZN(_02634_ ) );
BUF_X4 _10231_ ( .A(_02634_ ), .Z(_02635_ ) );
INV_X1 _10232_ ( .A(\ID_EX_imm [18] ), .ZN(_02636_ ) );
XNOR2_X1 _10233_ ( .A(_02635_ ), .B(_02636_ ), .ZN(_02637_ ) );
NAND2_X1 _10234_ ( .A1(_02460_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02638_ ) );
OR2_X1 _10235_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02639_ ) );
OAI211_X1 _10236_ ( .A(_02639_ ), .B(_02547_ ), .C1(_02363_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02640_ ) );
OR2_X1 _10237_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02641_ ) );
OAI211_X1 _10238_ ( .A(_02641_ ), .B(fanout_net_26 ), .C1(_02363_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02642_ ) );
NAND3_X1 _10239_ ( .A1(_02640_ ), .A2(_02642_ ), .A3(_02349_ ), .ZN(_02643_ ) );
MUX2_X1 _10240_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02644_ ) );
MUX2_X1 _10241_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02645_ ) );
MUX2_X1 _10242_ ( .A(_02644_ ), .B(_02645_ ), .S(_02547_ ), .Z(_02646_ ) );
OAI211_X1 _10243_ ( .A(_02326_ ), .B(_02643_ ), .C1(_02646_ ), .C2(_02517_ ), .ZN(_02647_ ) );
OR2_X1 _10244_ ( .A1(_02339_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02648_ ) );
OAI211_X1 _10245_ ( .A(_02648_ ), .B(_02547_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02649_ ) );
OR2_X1 _10246_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02650_ ) );
OAI211_X1 _10247_ ( .A(_02650_ ), .B(fanout_net_26 ), .C1(_02363_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02651_ ) );
NAND3_X1 _10248_ ( .A1(_02649_ ), .A2(fanout_net_28 ), .A3(_02651_ ), .ZN(_02652_ ) );
MUX2_X1 _10249_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02653_ ) );
MUX2_X1 _10250_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02654_ ) );
MUX2_X1 _10251_ ( .A(_02653_ ), .B(_02654_ ), .S(fanout_net_26 ), .Z(_02655_ ) );
OAI211_X1 _10252_ ( .A(fanout_net_29 ), .B(_02652_ ), .C1(_02655_ ), .C2(fanout_net_28 ), .ZN(_02656_ ) );
NAND2_X1 _10253_ ( .A1(_02647_ ), .A2(_02656_ ), .ZN(_02657_ ) );
OAI21_X2 _10254_ ( .A(_02657_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02658_ ) );
AND3_X1 _10255_ ( .A1(_02638_ ), .A2(\ID_EX_imm [19] ), .A3(_02658_ ), .ZN(_02659_ ) );
AOI21_X1 _10256_ ( .A(\ID_EX_imm [19] ), .B1(_02638_ ), .B2(_02658_ ), .ZN(_02660_ ) );
NOR2_X1 _10257_ ( .A1(_02659_ ), .A2(_02660_ ), .ZN(_02661_ ) );
AND2_X1 _10258_ ( .A1(_02637_ ), .A2(_02661_ ), .ZN(_02662_ ) );
NAND2_X1 _10259_ ( .A1(_02460_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02663_ ) );
NOR2_X1 _10260_ ( .A1(_02340_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02664_ ) );
OAI21_X1 _10261_ ( .A(fanout_net_27 ), .B1(fanout_net_20 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02665_ ) );
NOR2_X1 _10262_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02666_ ) );
OAI21_X1 _10263_ ( .A(_02333_ ), .B1(_02340_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02667_ ) );
OAI221_X1 _10264_ ( .A(_02517_ ), .B1(_02664_ ), .B2(_02665_ ), .C1(_02666_ ), .C2(_02667_ ), .ZN(_02668_ ) );
MUX2_X1 _10265_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02669_ ) );
MUX2_X1 _10266_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02670_ ) );
MUX2_X1 _10267_ ( .A(_02669_ ), .B(_02670_ ), .S(fanout_net_27 ), .Z(_02671_ ) );
OAI211_X1 _10268_ ( .A(fanout_net_29 ), .B(_02668_ ), .C1(_02671_ ), .C2(_02350_ ), .ZN(_02672_ ) );
OR2_X1 _10269_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02673_ ) );
OAI211_X1 _10270_ ( .A(_02673_ ), .B(_02591_ ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02674_ ) );
OR2_X1 _10271_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02675_ ) );
OAI211_X1 _10272_ ( .A(_02675_ ), .B(fanout_net_27 ), .C1(_02340_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02676_ ) );
NAND3_X1 _10273_ ( .A1(_02674_ ), .A2(_02676_ ), .A3(fanout_net_28 ), .ZN(_02677_ ) );
MUX2_X1 _10274_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02678_ ) );
MUX2_X1 _10275_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02679_ ) );
MUX2_X1 _10276_ ( .A(_02678_ ), .B(_02679_ ), .S(_02333_ ), .Z(_02680_ ) );
OAI211_X1 _10277_ ( .A(_02326_ ), .B(_02677_ ), .C1(_02680_ ), .C2(fanout_net_28 ), .ZN(_02681_ ) );
NAND2_X1 _10278_ ( .A1(_02672_ ), .A2(_02681_ ), .ZN(_02682_ ) );
OAI21_X1 _10279_ ( .A(_02682_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02683_ ) );
AND2_X2 _10280_ ( .A1(_02663_ ), .A2(_02683_ ), .ZN(_02684_ ) );
INV_X1 _10281_ ( .A(\ID_EX_imm [17] ), .ZN(_02685_ ) );
XNOR2_X1 _10282_ ( .A(_02684_ ), .B(_02685_ ), .ZN(_02686_ ) );
NAND2_X1 _10283_ ( .A1(_02460_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02687_ ) );
OR2_X1 _10284_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02688_ ) );
OAI211_X1 _10285_ ( .A(_02688_ ), .B(_02591_ ), .C1(_02341_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02689_ ) );
OR2_X1 _10286_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02690_ ) );
OAI211_X1 _10287_ ( .A(_02690_ ), .B(fanout_net_27 ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02691_ ) );
NAND3_X1 _10288_ ( .A1(_02689_ ), .A2(_02691_ ), .A3(_02350_ ), .ZN(_02692_ ) );
MUX2_X1 _10289_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02693_ ) );
MUX2_X1 _10290_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02694_ ) );
MUX2_X1 _10291_ ( .A(_02693_ ), .B(_02694_ ), .S(_02591_ ), .Z(_02695_ ) );
OAI211_X1 _10292_ ( .A(_02326_ ), .B(_02692_ ), .C1(_02695_ ), .C2(_02350_ ), .ZN(_02696_ ) );
OR2_X1 _10293_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02697_ ) );
OAI211_X1 _10294_ ( .A(_02697_ ), .B(fanout_net_27 ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02698_ ) );
OR2_X1 _10295_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02699_ ) );
OAI211_X1 _10296_ ( .A(_02699_ ), .B(_02591_ ), .C1(_02364_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02700_ ) );
NAND3_X1 _10297_ ( .A1(_02698_ ), .A2(_02700_ ), .A3(fanout_net_28 ), .ZN(_02701_ ) );
MUX2_X1 _10298_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02702_ ) );
MUX2_X1 _10299_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02703_ ) );
MUX2_X1 _10300_ ( .A(_02702_ ), .B(_02703_ ), .S(fanout_net_27 ), .Z(_02704_ ) );
OAI211_X1 _10301_ ( .A(fanout_net_29 ), .B(_02701_ ), .C1(_02704_ ), .C2(fanout_net_28 ), .ZN(_02705_ ) );
NAND2_X1 _10302_ ( .A1(_02696_ ), .A2(_02705_ ), .ZN(_02706_ ) );
OAI21_X1 _10303_ ( .A(_02706_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02707_ ) );
AND2_X1 _10304_ ( .A1(_02687_ ), .A2(_02707_ ), .ZN(_02708_ ) );
BUF_X4 _10305_ ( .A(_02708_ ), .Z(_02709_ ) );
INV_X1 _10306_ ( .A(\ID_EX_imm [16] ), .ZN(_02710_ ) );
XNOR2_X1 _10307_ ( .A(_02709_ ), .B(_02710_ ), .ZN(_02711_ ) );
NAND3_X1 _10308_ ( .A1(_02662_ ), .A2(_02686_ ), .A3(_02711_ ), .ZN(_02712_ ) );
NAND2_X4 _10309_ ( .A1(_02460_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02713_ ) );
NOR2_X1 _10310_ ( .A1(_02362_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02714_ ) );
OAI21_X1 _10311_ ( .A(fanout_net_27 ), .B1(fanout_net_21 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02715_ ) );
NOR2_X1 _10312_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02716_ ) );
OAI21_X1 _10313_ ( .A(_02546_ ), .B1(_02362_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02717_ ) );
OAI221_X1 _10314_ ( .A(_02348_ ), .B1(_02714_ ), .B2(_02715_ ), .C1(_02716_ ), .C2(_02717_ ), .ZN(_02718_ ) );
MUX2_X1 _10315_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02719_ ) );
MUX2_X1 _10316_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02720_ ) );
MUX2_X1 _10317_ ( .A(_02719_ ), .B(_02720_ ), .S(fanout_net_27 ), .Z(_02721_ ) );
OAI211_X1 _10318_ ( .A(fanout_net_29 ), .B(_02718_ ), .C1(_02721_ ), .C2(_02348_ ), .ZN(_02722_ ) );
BUF_X2 _10319_ ( .A(_02336_ ), .Z(_02723_ ) );
OR2_X1 _10320_ ( .A1(_02723_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02724_ ) );
OAI211_X1 _10321_ ( .A(_02724_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02725_ ) );
OR2_X1 _10322_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02726_ ) );
OAI211_X1 _10323_ ( .A(_02726_ ), .B(_02546_ ), .C1(_02362_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02727_ ) );
NAND3_X1 _10324_ ( .A1(_02725_ ), .A2(fanout_net_28 ), .A3(_02727_ ), .ZN(_02728_ ) );
MUX2_X1 _10325_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02729_ ) );
MUX2_X1 _10326_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02730_ ) );
MUX2_X1 _10327_ ( .A(_02729_ ), .B(_02730_ ), .S(_02546_ ), .Z(_02731_ ) );
OAI211_X1 _10328_ ( .A(_02325_ ), .B(_02728_ ), .C1(_02731_ ), .C2(fanout_net_28 ), .ZN(_02732_ ) );
NAND2_X1 _10329_ ( .A1(_02722_ ), .A2(_02732_ ), .ZN(_02733_ ) );
OAI21_X4 _10330_ ( .A(_02733_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02734_ ) );
AND2_X4 _10331_ ( .A1(_02713_ ), .A2(_02734_ ), .ZN(_02735_ ) );
INV_X1 _10332_ ( .A(\ID_EX_imm [4] ), .ZN(_02736_ ) );
XNOR2_X1 _10333_ ( .A(_02735_ ), .B(_02736_ ), .ZN(_02737_ ) );
INV_X1 _10334_ ( .A(_02737_ ), .ZN(_02738_ ) );
NAND2_X4 _10335_ ( .A1(_02459_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02739_ ) );
OR2_X1 _10336_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02740_ ) );
OAI211_X1 _10337_ ( .A(_02740_ ), .B(fanout_net_27 ), .C1(_02338_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02741_ ) );
INV_X1 _10338_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02742_ ) );
NAND2_X1 _10339_ ( .A1(_02742_ ), .A2(fanout_net_21 ), .ZN(_02743_ ) );
BUF_X4 _10340_ ( .A(_02329_ ), .Z(_02744_ ) );
OAI211_X1 _10341_ ( .A(_02743_ ), .B(_02744_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02745_ ) );
NAND3_X1 _10342_ ( .A1(_02741_ ), .A2(_02745_ ), .A3(_02347_ ), .ZN(_02746_ ) );
MUX2_X1 _10343_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02747_ ) );
MUX2_X1 _10344_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02748_ ) );
MUX2_X1 _10345_ ( .A(_02747_ ), .B(_02748_ ), .S(_02744_ ), .Z(_02749_ ) );
BUF_X4 _10346_ ( .A(_02346_ ), .Z(_02750_ ) );
OAI211_X1 _10347_ ( .A(_02325_ ), .B(_02746_ ), .C1(_02749_ ), .C2(_02750_ ), .ZN(_02751_ ) );
OR2_X1 _10348_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02752_ ) );
OAI211_X1 _10349_ ( .A(_02752_ ), .B(_02744_ ), .C1(_02338_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02753_ ) );
OR2_X1 _10350_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02754_ ) );
OAI211_X1 _10351_ ( .A(_02754_ ), .B(fanout_net_27 ), .C1(_02338_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02755_ ) );
NAND3_X1 _10352_ ( .A1(_02753_ ), .A2(_02755_ ), .A3(fanout_net_28 ), .ZN(_02756_ ) );
MUX2_X1 _10353_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02757_ ) );
MUX2_X1 _10354_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02758_ ) );
MUX2_X1 _10355_ ( .A(_02757_ ), .B(_02758_ ), .S(fanout_net_27 ), .Z(_02759_ ) );
OAI211_X1 _10356_ ( .A(fanout_net_29 ), .B(_02756_ ), .C1(_02759_ ), .C2(fanout_net_28 ), .ZN(_02760_ ) );
NAND2_X1 _10357_ ( .A1(_02751_ ), .A2(_02760_ ), .ZN(_02761_ ) );
OAI21_X1 _10358_ ( .A(_02761_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_02762_ ) );
AND2_X2 _10359_ ( .A1(_02739_ ), .A2(_02762_ ), .ZN(_02763_ ) );
BUF_X8 _10360_ ( .A(_02763_ ), .Z(_02764_ ) );
XNOR2_X2 _10361_ ( .A(_02764_ ), .B(\ID_EX_imm [5] ), .ZN(_02765_ ) );
NOR2_X1 _10362_ ( .A1(_02738_ ), .A2(_02765_ ), .ZN(_02766_ ) );
OR2_X1 _10363_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02767_ ) );
OAI211_X1 _10364_ ( .A(_02767_ ), .B(_02547_ ), .C1(_02363_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02768_ ) );
OR2_X1 _10365_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02769_ ) );
OAI211_X1 _10366_ ( .A(_02769_ ), .B(fanout_net_27 ), .C1(_02363_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02770_ ) );
NAND3_X1 _10367_ ( .A1(_02768_ ), .A2(_02770_ ), .A3(_02349_ ), .ZN(_02771_ ) );
MUX2_X1 _10368_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02772_ ) );
MUX2_X1 _10369_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02773_ ) );
MUX2_X1 _10370_ ( .A(_02772_ ), .B(_02773_ ), .S(_02332_ ), .Z(_02774_ ) );
OAI211_X1 _10371_ ( .A(fanout_net_29 ), .B(_02771_ ), .C1(_02774_ ), .C2(_02517_ ), .ZN(_02775_ ) );
MUX2_X1 _10372_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02776_ ) );
AND2_X1 _10373_ ( .A1(_02776_ ), .A2(_02547_ ), .ZN(_02777_ ) );
MUX2_X1 _10374_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02778_ ) );
AOI211_X1 _10375_ ( .A(fanout_net_28 ), .B(_02777_ ), .C1(fanout_net_27 ), .C2(_02778_ ), .ZN(_02779_ ) );
MUX2_X1 _10376_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02780_ ) );
MUX2_X1 _10377_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02781_ ) );
MUX2_X1 _10378_ ( .A(_02780_ ), .B(_02781_ ), .S(_02332_ ), .Z(_02782_ ) );
OAI21_X1 _10379_ ( .A(_02326_ ), .B1(_02782_ ), .B2(_02517_ ), .ZN(_02783_ ) );
OAI21_X1 _10380_ ( .A(_02775_ ), .B1(_02779_ ), .B2(_02783_ ), .ZN(_02784_ ) );
OAI21_X1 _10381_ ( .A(_02784_ ), .B1(_02485_ ), .B2(_02483_ ), .ZN(_02785_ ) );
NAND2_X1 _10382_ ( .A1(_02460_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02786_ ) );
AND2_X2 _10383_ ( .A1(_02785_ ), .A2(_02786_ ), .ZN(_02787_ ) );
BUF_X4 _10384_ ( .A(_02787_ ), .Z(_02788_ ) );
XOR2_X2 _10385_ ( .A(_02788_ ), .B(\ID_EX_imm [6] ), .Z(_02789_ ) );
NAND2_X1 _10386_ ( .A1(_02460_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02790_ ) );
OR2_X1 _10387_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02791_ ) );
OAI211_X1 _10388_ ( .A(_02791_ ), .B(_02547_ ), .C1(_02339_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02792_ ) );
OR2_X1 _10389_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02793_ ) );
OAI211_X1 _10390_ ( .A(_02793_ ), .B(fanout_net_27 ), .C1(_02339_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02794_ ) );
NAND3_X1 _10391_ ( .A1(_02792_ ), .A2(_02794_ ), .A3(_02349_ ), .ZN(_02795_ ) );
MUX2_X1 _10392_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02796_ ) );
MUX2_X1 _10393_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02797_ ) );
MUX2_X1 _10394_ ( .A(_02796_ ), .B(_02797_ ), .S(_02332_ ), .Z(_02798_ ) );
OAI211_X1 _10395_ ( .A(_02326_ ), .B(_02795_ ), .C1(_02798_ ), .C2(_02349_ ), .ZN(_02799_ ) );
OR2_X1 _10396_ ( .A1(_02362_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02800_ ) );
OAI211_X1 _10397_ ( .A(_02800_ ), .B(fanout_net_27 ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02801_ ) );
OR2_X1 _10398_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02802_ ) );
OAI211_X1 _10399_ ( .A(_02802_ ), .B(_02332_ ), .C1(_02339_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02803_ ) );
NAND3_X1 _10400_ ( .A1(_02801_ ), .A2(fanout_net_28 ), .A3(_02803_ ), .ZN(_02804_ ) );
MUX2_X1 _10401_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02805_ ) );
MUX2_X1 _10402_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02806_ ) );
MUX2_X1 _10403_ ( .A(_02805_ ), .B(_02806_ ), .S(fanout_net_27 ), .Z(_02807_ ) );
OAI211_X1 _10404_ ( .A(fanout_net_29 ), .B(_02804_ ), .C1(_02807_ ), .C2(fanout_net_28 ), .ZN(_02808_ ) );
NAND2_X1 _10405_ ( .A1(_02799_ ), .A2(_02808_ ), .ZN(_02809_ ) );
OAI21_X1 _10406_ ( .A(_02809_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02810_ ) );
AND2_X2 _10407_ ( .A1(_02790_ ), .A2(_02810_ ), .ZN(_02811_ ) );
BUF_X4 _10408_ ( .A(_02811_ ), .Z(_02812_ ) );
XOR2_X1 _10409_ ( .A(_02812_ ), .B(\ID_EX_imm [7] ), .Z(_02813_ ) );
AND2_X1 _10410_ ( .A1(_02789_ ), .A2(_02813_ ), .ZN(_02814_ ) );
OR3_X4 _10411_ ( .A1(_02388_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02395_ ), .ZN(_02815_ ) );
OR2_X1 _10412_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02816_ ) );
OAI211_X1 _10413_ ( .A(_02816_ ), .B(_02332_ ), .C1(_02339_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02817_ ) );
OR2_X1 _10414_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02818_ ) );
OAI211_X1 _10415_ ( .A(_02818_ ), .B(fanout_net_27 ), .C1(_02362_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02819_ ) );
NAND3_X1 _10416_ ( .A1(_02817_ ), .A2(_02819_ ), .A3(_02348_ ), .ZN(_02820_ ) );
MUX2_X1 _10417_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02821_ ) );
MUX2_X1 _10418_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02822_ ) );
MUX2_X1 _10419_ ( .A(_02821_ ), .B(_02822_ ), .S(_02332_ ), .Z(_02823_ ) );
OAI211_X1 _10420_ ( .A(_02325_ ), .B(_02820_ ), .C1(_02823_ ), .C2(_02349_ ), .ZN(_02824_ ) );
OR2_X1 _10421_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02825_ ) );
OAI211_X1 _10422_ ( .A(_02825_ ), .B(fanout_net_27 ), .C1(_02339_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02826_ ) );
OR2_X1 _10423_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02827_ ) );
OAI211_X1 _10424_ ( .A(_02827_ ), .B(_02332_ ), .C1(_02362_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02828_ ) );
NAND3_X1 _10425_ ( .A1(_02826_ ), .A2(_02828_ ), .A3(fanout_net_28 ), .ZN(_02829_ ) );
MUX2_X1 _10426_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02830_ ) );
MUX2_X1 _10427_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02831_ ) );
MUX2_X1 _10428_ ( .A(_02830_ ), .B(_02831_ ), .S(fanout_net_27 ), .Z(_02832_ ) );
OAI211_X1 _10429_ ( .A(fanout_net_29 ), .B(_02829_ ), .C1(_02832_ ), .C2(fanout_net_28 ), .ZN(_02833_ ) );
OAI211_X2 _10430_ ( .A(_02824_ ), .B(_02833_ ), .C1(_02388_ ), .C2(_02395_ ), .ZN(_02834_ ) );
NAND2_X4 _10431_ ( .A1(_02815_ ), .A2(_02834_ ), .ZN(_02835_ ) );
INV_X1 _10432_ ( .A(\ID_EX_imm [1] ), .ZN(_02836_ ) );
XNOR2_X2 _10433_ ( .A(_02835_ ), .B(_02836_ ), .ZN(_02837_ ) );
NAND2_X1 _10434_ ( .A1(_02460_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_02838_ ) );
OR2_X1 _10435_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(fanout_net_22 ), .ZN(_02839_ ) );
BUF_X4 _10436_ ( .A(_02337_ ), .Z(_02840_ ) );
OAI211_X1 _10437_ ( .A(_02839_ ), .B(_02546_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_02840_ ), .ZN(_02841_ ) );
NOR2_X1 _10438_ ( .A1(_02362_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02842_ ) );
OAI21_X1 _10439_ ( .A(fanout_net_27 ), .B1(fanout_net_22 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02843_ ) );
OAI211_X1 _10440_ ( .A(_02841_ ), .B(_02750_ ), .C1(_02842_ ), .C2(_02843_ ), .ZN(_02844_ ) );
MUX2_X1 _10441_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02845_ ) );
MUX2_X1 _10442_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02846_ ) );
MUX2_X1 _10443_ ( .A(_02845_ ), .B(_02846_ ), .S(_02546_ ), .Z(_02847_ ) );
OAI211_X1 _10444_ ( .A(_02325_ ), .B(_02844_ ), .C1(_02847_ ), .C2(_02348_ ), .ZN(_02848_ ) );
OR2_X1 _10445_ ( .A1(fanout_net_23 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02849_ ) );
OAI211_X1 _10446_ ( .A(_02849_ ), .B(_02546_ ), .C1(_02362_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02850_ ) );
OR2_X1 _10447_ ( .A1(fanout_net_23 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02851_ ) );
OAI211_X1 _10448_ ( .A(_02851_ ), .B(fanout_net_27 ), .C1(_02362_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02852_ ) );
NAND3_X1 _10449_ ( .A1(_02850_ ), .A2(_02852_ ), .A3(_02348_ ), .ZN(_02853_ ) );
MUX2_X1 _10450_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02854_ ) );
MUX2_X1 _10451_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02855_ ) );
MUX2_X1 _10452_ ( .A(_02854_ ), .B(_02855_ ), .S(_02546_ ), .Z(_02856_ ) );
OAI211_X1 _10453_ ( .A(fanout_net_29 ), .B(_02853_ ), .C1(_02856_ ), .C2(_02348_ ), .ZN(_02857_ ) );
NAND2_X1 _10454_ ( .A1(_02848_ ), .A2(_02857_ ), .ZN(_02858_ ) );
OAI21_X4 _10455_ ( .A(_02858_ ), .B1(_02483_ ), .B2(_02485_ ), .ZN(_02859_ ) );
AND3_X1 _10456_ ( .A1(_02838_ ), .A2(\ID_EX_imm [0] ), .A3(_02859_ ), .ZN(_02860_ ) );
NAND2_X1 _10457_ ( .A1(_02837_ ), .A2(_02860_ ), .ZN(_02861_ ) );
INV_X1 _10458_ ( .A(_02835_ ), .ZN(_02862_ ) );
OAI21_X1 _10459_ ( .A(_02861_ ), .B1(_02836_ ), .B2(_02862_ ), .ZN(_02863_ ) );
NAND2_X4 _10460_ ( .A1(_02459_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02864_ ) );
OR2_X1 _10461_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02865_ ) );
OAI211_X1 _10462_ ( .A(_02865_ ), .B(_02744_ ), .C1(_02338_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02866_ ) );
OR2_X1 _10463_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02867_ ) );
OAI211_X1 _10464_ ( .A(_02867_ ), .B(fanout_net_27 ), .C1(_02723_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02868_ ) );
NAND3_X1 _10465_ ( .A1(_02866_ ), .A2(_02868_ ), .A3(_02347_ ), .ZN(_02869_ ) );
MUX2_X1 _10466_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02870_ ) );
MUX2_X1 _10467_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02871_ ) );
MUX2_X1 _10468_ ( .A(_02870_ ), .B(_02871_ ), .S(_02330_ ), .Z(_02872_ ) );
OAI211_X1 _10469_ ( .A(_02324_ ), .B(_02869_ ), .C1(_02872_ ), .C2(_02750_ ), .ZN(_02873_ ) );
OR2_X1 _10470_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02874_ ) );
OAI211_X1 _10471_ ( .A(_02874_ ), .B(fanout_net_27 ), .C1(_02723_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02875_ ) );
OR2_X1 _10472_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02876_ ) );
OAI211_X1 _10473_ ( .A(_02876_ ), .B(_02744_ ), .C1(_02723_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02877_ ) );
NAND3_X1 _10474_ ( .A1(_02875_ ), .A2(_02877_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02878_ ) );
MUX2_X1 _10475_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02879_ ) );
MUX2_X1 _10476_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02880_ ) );
MUX2_X1 _10477_ ( .A(_02879_ ), .B(_02880_ ), .S(fanout_net_27 ), .Z(_02881_ ) );
OAI211_X1 _10478_ ( .A(fanout_net_29 ), .B(_02878_ ), .C1(_02881_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02882_ ) );
NAND2_X1 _10479_ ( .A1(_02873_ ), .A2(_02882_ ), .ZN(_02883_ ) );
OAI21_X4 _10480_ ( .A(_02883_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_02884_ ) );
AND2_X4 _10481_ ( .A1(_02864_ ), .A2(_02884_ ), .ZN(_02885_ ) );
BUF_X8 _10482_ ( .A(_02885_ ), .Z(_02886_ ) );
XOR2_X1 _10483_ ( .A(_02886_ ), .B(\ID_EX_imm [2] ), .Z(_02887_ ) );
AND2_X1 _10484_ ( .A1(_02863_ ), .A2(_02887_ ), .ZN(_02888_ ) );
AND3_X1 _10485_ ( .A1(_02864_ ), .A2(\ID_EX_imm [2] ), .A3(_02884_ ), .ZN(_02889_ ) );
OR2_X2 _10486_ ( .A1(_02888_ ), .A2(_02889_ ), .ZN(_02890_ ) );
OR2_X1 _10487_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02891_ ) );
OAI211_X1 _10488_ ( .A(_02891_ ), .B(_02331_ ), .C1(_02840_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02892_ ) );
OR2_X1 _10489_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02893_ ) );
OAI211_X1 _10490_ ( .A(_02893_ ), .B(fanout_net_27 ), .C1(_02840_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02894_ ) );
NAND3_X1 _10491_ ( .A1(_02892_ ), .A2(_02894_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02895_ ) );
MUX2_X1 _10492_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02896_ ) );
MUX2_X1 _10493_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02897_ ) );
MUX2_X1 _10494_ ( .A(_02896_ ), .B(_02897_ ), .S(_02331_ ), .Z(_02898_ ) );
OAI211_X1 _10495_ ( .A(_02325_ ), .B(_02895_ ), .C1(_02898_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02899_ ) );
MUX2_X1 _10496_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02900_ ) );
AND2_X1 _10497_ ( .A1(_02900_ ), .A2(fanout_net_27 ), .ZN(_02901_ ) );
MUX2_X1 _10498_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02902_ ) );
AOI211_X1 _10499_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_02901_ ), .C1(_02332_ ), .C2(_02902_ ), .ZN(_02903_ ) );
MUX2_X1 _10500_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02904_ ) );
MUX2_X1 _10501_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02905_ ) );
MUX2_X1 _10502_ ( .A(_02904_ ), .B(_02905_ ), .S(fanout_net_27 ), .Z(_02906_ ) );
OAI21_X1 _10503_ ( .A(fanout_net_29 ), .B1(_02906_ ), .B2(_02750_ ), .ZN(_02907_ ) );
OAI221_X2 _10504_ ( .A(_02899_ ), .B1(_02903_ ), .B2(_02907_ ), .C1(_02388_ ), .C2(_02395_ ), .ZN(_02908_ ) );
OR3_X4 _10505_ ( .A1(_02388_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02395_ ), .ZN(_02909_ ) );
NAND2_X4 _10506_ ( .A1(_02908_ ), .A2(_02909_ ), .ZN(_02910_ ) );
INV_X1 _10507_ ( .A(\ID_EX_imm [3] ), .ZN(_02911_ ) );
XNOR2_X1 _10508_ ( .A(_02910_ ), .B(_02911_ ), .ZN(_02912_ ) );
AND2_X1 _10509_ ( .A1(_02890_ ), .A2(_02912_ ), .ZN(_02913_ ) );
AOI21_X1 _10510_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B1(_02908_ ), .B2(_02909_ ), .ZN(_02914_ ) );
OAI211_X1 _10511_ ( .A(_02766_ ), .B(_02814_ ), .C1(_02913_ ), .C2(_02914_ ), .ZN(_02915_ ) );
XNOR2_X1 _10512_ ( .A(_02812_ ), .B(\ID_EX_imm [7] ), .ZN(_02916_ ) );
NAND2_X1 _10513_ ( .A1(_02788_ ), .A2(\ID_EX_imm [6] ), .ZN(_02917_ ) );
NOR2_X1 _10514_ ( .A1(_02916_ ), .A2(_02917_ ), .ZN(_02918_ ) );
INV_X2 _10515_ ( .A(_02735_ ), .ZN(_02919_ ) );
NOR3_X1 _10516_ ( .A1(_02765_ ), .A2(_02736_ ), .A3(_02919_ ), .ZN(_02920_ ) );
INV_X1 _10517_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02921_ ) );
AOI21_X1 _10518_ ( .A(_02920_ ), .B1(_02921_ ), .B2(_02764_ ), .ZN(_02922_ ) );
INV_X1 _10519_ ( .A(_02922_ ), .ZN(_02923_ ) );
AOI221_X4 _10520_ ( .A(_02918_ ), .B1(\ID_EX_imm [7] ), .B2(_02812_ ), .C1(_02923_ ), .C2(_02814_ ), .ZN(_02924_ ) );
NAND2_X2 _10521_ ( .A1(_02915_ ), .A2(_02924_ ), .ZN(_02925_ ) );
NAND2_X1 _10522_ ( .A1(_02459_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02926_ ) );
OR2_X1 _10523_ ( .A1(_02337_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02927_ ) );
OAI211_X1 _10524_ ( .A(_02927_ ), .B(fanout_net_27 ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02928_ ) );
OR2_X1 _10525_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02929_ ) );
OAI211_X1 _10526_ ( .A(_02929_ ), .B(_02331_ ), .C1(_02338_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02930_ ) );
NAND3_X1 _10527_ ( .A1(_02928_ ), .A2(_02750_ ), .A3(_02930_ ), .ZN(_02931_ ) );
MUX2_X1 _10528_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02932_ ) );
MUX2_X1 _10529_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02933_ ) );
MUX2_X1 _10530_ ( .A(_02932_ ), .B(_02933_ ), .S(_02744_ ), .Z(_02934_ ) );
OAI211_X1 _10531_ ( .A(_02325_ ), .B(_02931_ ), .C1(_02934_ ), .C2(_02348_ ), .ZN(_02935_ ) );
OR2_X1 _10532_ ( .A1(_02337_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02936_ ) );
OAI211_X1 _10533_ ( .A(_02936_ ), .B(fanout_net_27 ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02937_ ) );
OR2_X1 _10534_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02938_ ) );
OAI211_X1 _10535_ ( .A(_02938_ ), .B(_02331_ ), .C1(_02338_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02939_ ) );
NAND3_X1 _10536_ ( .A1(_02937_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02939_ ), .ZN(_02940_ ) );
MUX2_X1 _10537_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02941_ ) );
MUX2_X1 _10538_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02942_ ) );
MUX2_X1 _10539_ ( .A(_02941_ ), .B(_02942_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02943_ ) );
OAI211_X1 _10540_ ( .A(fanout_net_29 ), .B(_02940_ ), .C1(_02943_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02944_ ) );
NAND2_X1 _10541_ ( .A1(_02935_ ), .A2(_02944_ ), .ZN(_02945_ ) );
OAI21_X2 _10542_ ( .A(_02945_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_02946_ ) );
AND2_X4 _10543_ ( .A1(_02926_ ), .A2(_02946_ ), .ZN(_02947_ ) );
BUF_X8 _10544_ ( .A(_02947_ ), .Z(_02948_ ) );
XOR2_X1 _10545_ ( .A(_02948_ ), .B(\ID_EX_imm [12] ), .Z(_02949_ ) );
NAND2_X1 _10546_ ( .A1(_02459_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02950_ ) );
OR2_X1 _10547_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02951_ ) );
OAI211_X1 _10548_ ( .A(_02951_ ), .B(_02331_ ), .C1(_02338_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02952_ ) );
OR2_X1 _10549_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02953_ ) );
OAI211_X1 _10550_ ( .A(_02953_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02338_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02954_ ) );
NAND3_X1 _10551_ ( .A1(_02952_ ), .A2(_02954_ ), .A3(_02347_ ), .ZN(_02955_ ) );
MUX2_X1 _10552_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02956_ ) );
MUX2_X1 _10553_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02957_ ) );
MUX2_X1 _10554_ ( .A(_02956_ ), .B(_02957_ ), .S(_02744_ ), .Z(_02958_ ) );
OAI211_X1 _10555_ ( .A(_02325_ ), .B(_02955_ ), .C1(_02958_ ), .C2(_02750_ ), .ZN(_02959_ ) );
OR2_X1 _10556_ ( .A1(_02336_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02960_ ) );
OAI211_X1 _10557_ ( .A(_02960_ ), .B(_02744_ ), .C1(fanout_net_24 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02961_ ) );
OR2_X1 _10558_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02962_ ) );
OAI211_X1 _10559_ ( .A(_02962_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02723_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02963_ ) );
NAND3_X1 _10560_ ( .A1(_02961_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02963_ ), .ZN(_02964_ ) );
MUX2_X1 _10561_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02965_ ) );
MUX2_X1 _10562_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02966_ ) );
MUX2_X1 _10563_ ( .A(_02965_ ), .B(_02966_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02967_ ) );
OAI211_X1 _10564_ ( .A(fanout_net_29 ), .B(_02964_ ), .C1(_02967_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02968_ ) );
NAND2_X1 _10565_ ( .A1(_02959_ ), .A2(_02968_ ), .ZN(_02969_ ) );
OAI21_X2 _10566_ ( .A(_02969_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_02970_ ) );
AOI21_X1 _10567_ ( .A(\ID_EX_imm [13] ), .B1(_02950_ ), .B2(_02970_ ), .ZN(_02971_ ) );
INV_X1 _10568_ ( .A(_02971_ ), .ZN(_02972_ ) );
NAND3_X1 _10569_ ( .A1(_02950_ ), .A2(\ID_EX_imm [13] ), .A3(_02970_ ), .ZN(_02973_ ) );
AND3_X1 _10570_ ( .A1(_02949_ ), .A2(_02972_ ), .A3(_02973_ ), .ZN(_02974_ ) );
NAND2_X1 _10571_ ( .A1(_02459_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02975_ ) );
NOR2_X1 _10572_ ( .A1(_02338_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02976_ ) );
OAI21_X1 _10573_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_24 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02977_ ) );
NOR2_X1 _10574_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02978_ ) );
OAI21_X1 _10575_ ( .A(_02331_ ), .B1(_02840_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02979_ ) );
OAI221_X1 _10576_ ( .A(_02750_ ), .B1(_02976_ ), .B2(_02977_ ), .C1(_02978_ ), .C2(_02979_ ), .ZN(_02980_ ) );
MUX2_X1 _10577_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02981_ ) );
MUX2_X1 _10578_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02982_ ) );
MUX2_X1 _10579_ ( .A(_02981_ ), .B(_02982_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02983_ ) );
OAI211_X1 _10580_ ( .A(fanout_net_29 ), .B(_02980_ ), .C1(_02983_ ), .C2(_02348_ ), .ZN(_02984_ ) );
OR2_X1 _10581_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02985_ ) );
OAI211_X1 _10582_ ( .A(_02985_ ), .B(_02546_ ), .C1(_02840_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02986_ ) );
OR2_X1 _10583_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02987_ ) );
OAI211_X1 _10584_ ( .A(_02987_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02840_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02988_ ) );
NAND3_X1 _10585_ ( .A1(_02986_ ), .A2(_02988_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02989_ ) );
MUX2_X1 _10586_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02990_ ) );
MUX2_X1 _10587_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02991_ ) );
MUX2_X1 _10588_ ( .A(_02990_ ), .B(_02991_ ), .S(_02331_ ), .Z(_02992_ ) );
OAI211_X1 _10589_ ( .A(_02325_ ), .B(_02989_ ), .C1(_02992_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02993_ ) );
NAND2_X1 _10590_ ( .A1(_02984_ ), .A2(_02993_ ), .ZN(_02994_ ) );
OAI21_X2 _10591_ ( .A(_02994_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_02995_ ) );
AND2_X4 _10592_ ( .A1(_02975_ ), .A2(_02995_ ), .ZN(_02996_ ) );
XOR2_X1 _10593_ ( .A(_02996_ ), .B(\ID_EX_imm [15] ), .Z(_02997_ ) );
NAND2_X1 _10594_ ( .A1(_02459_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02998_ ) );
OR2_X1 _10595_ ( .A1(_02336_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02999_ ) );
OAI211_X1 _10596_ ( .A(_02999_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_24 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03000_ ) );
OR2_X1 _10597_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03001_ ) );
OAI211_X1 _10598_ ( .A(_03001_ ), .B(_02744_ ), .C1(_02723_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03002_ ) );
NAND3_X1 _10599_ ( .A1(_03000_ ), .A2(_02347_ ), .A3(_03002_ ), .ZN(_03003_ ) );
MUX2_X1 _10600_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03004_ ) );
MUX2_X1 _10601_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03005_ ) );
MUX2_X1 _10602_ ( .A(_03004_ ), .B(_03005_ ), .S(_02330_ ), .Z(_03006_ ) );
OAI211_X1 _10603_ ( .A(_02324_ ), .B(_03003_ ), .C1(_03006_ ), .C2(_02750_ ), .ZN(_03007_ ) );
OR2_X1 _10604_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03008_ ) );
OAI211_X1 _10605_ ( .A(_03008_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02723_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03009_ ) );
OR2_X1 _10606_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03010_ ) );
OAI211_X1 _10607_ ( .A(_03010_ ), .B(_02330_ ), .C1(_02723_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03011_ ) );
NAND3_X1 _10608_ ( .A1(_03009_ ), .A2(_03011_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03012_ ) );
MUX2_X1 _10609_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03013_ ) );
MUX2_X1 _10610_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03014_ ) );
MUX2_X1 _10611_ ( .A(_03013_ ), .B(_03014_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03015_ ) );
OAI211_X1 _10612_ ( .A(fanout_net_29 ), .B(_03012_ ), .C1(_03015_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03016_ ) );
NAND2_X1 _10613_ ( .A1(_03007_ ), .A2(_03016_ ), .ZN(_03017_ ) );
OAI21_X4 _10614_ ( .A(_03017_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_03018_ ) );
AND2_X4 _10615_ ( .A1(_02998_ ), .A2(_03018_ ), .ZN(_03019_ ) );
BUF_X8 _10616_ ( .A(_03019_ ), .Z(_03020_ ) );
XOR2_X1 _10617_ ( .A(_03020_ ), .B(\ID_EX_imm [14] ), .Z(_03021_ ) );
AND3_X1 _10618_ ( .A1(_02974_ ), .A2(_02997_ ), .A3(_03021_ ), .ZN(_03022_ ) );
NAND2_X1 _10619_ ( .A1(_02459_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03023_ ) );
NOR2_X1 _10620_ ( .A1(_02840_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03024_ ) );
OAI21_X1 _10621_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_24 ), .B2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03025_ ) );
NOR2_X1 _10622_ ( .A1(fanout_net_24 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03026_ ) );
OAI21_X1 _10623_ ( .A(_02331_ ), .B1(_02840_ ), .B2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03027_ ) );
OAI221_X1 _10624_ ( .A(_02750_ ), .B1(_03024_ ), .B2(_03025_ ), .C1(_03026_ ), .C2(_03027_ ), .ZN(_03028_ ) );
MUX2_X1 _10625_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03029_ ) );
MUX2_X1 _10626_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03030_ ) );
MUX2_X1 _10627_ ( .A(_03029_ ), .B(_03030_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03031_ ) );
OAI211_X1 _10628_ ( .A(fanout_net_29 ), .B(_03028_ ), .C1(_03031_ ), .C2(_02348_ ), .ZN(_03032_ ) );
OR2_X1 _10629_ ( .A1(fanout_net_24 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03033_ ) );
OAI211_X1 _10630_ ( .A(_03033_ ), .B(_02546_ ), .C1(_02840_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03034_ ) );
OR2_X1 _10631_ ( .A1(fanout_net_24 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03035_ ) );
OAI211_X1 _10632_ ( .A(_03035_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02840_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03036_ ) );
NAND3_X1 _10633_ ( .A1(_03034_ ), .A2(_03036_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03037_ ) );
MUX2_X1 _10634_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03038_ ) );
MUX2_X1 _10635_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03039_ ) );
MUX2_X1 _10636_ ( .A(_03038_ ), .B(_03039_ ), .S(_02331_ ), .Z(_03040_ ) );
OAI211_X1 _10637_ ( .A(_02325_ ), .B(_03037_ ), .C1(_03040_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03041_ ) );
NAND2_X1 _10638_ ( .A1(_03032_ ), .A2(_03041_ ), .ZN(_03042_ ) );
OAI21_X1 _10639_ ( .A(_03042_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_03043_ ) );
AND2_X1 _10640_ ( .A1(_03023_ ), .A2(_03043_ ), .ZN(_03044_ ) );
BUF_X4 _10641_ ( .A(_03044_ ), .Z(_03045_ ) );
XOR2_X1 _10642_ ( .A(_03045_ ), .B(\ID_EX_imm [8] ), .Z(_03046_ ) );
NAND2_X1 _10643_ ( .A1(_02459_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03047_ ) );
OR2_X1 _10644_ ( .A1(_02336_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03048_ ) );
OAI211_X1 _10645_ ( .A(_03048_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_25 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03049_ ) );
OR2_X1 _10646_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03050_ ) );
OAI211_X1 _10647_ ( .A(_03050_ ), .B(_02329_ ), .C1(_02336_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03051_ ) );
NAND3_X1 _10648_ ( .A1(_03049_ ), .A2(_02346_ ), .A3(_03051_ ), .ZN(_03052_ ) );
MUX2_X1 _10649_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03053_ ) );
MUX2_X1 _10650_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03054_ ) );
MUX2_X1 _10651_ ( .A(_03053_ ), .B(_03054_ ), .S(_02329_ ), .Z(_03055_ ) );
OAI211_X1 _10652_ ( .A(fanout_net_29 ), .B(_03052_ ), .C1(_03055_ ), .C2(_02347_ ), .ZN(_03056_ ) );
OR2_X1 _10653_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03057_ ) );
OAI211_X1 _10654_ ( .A(_03057_ ), .B(_02330_ ), .C1(_02337_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03058_ ) );
OR2_X1 _10655_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03059_ ) );
OAI211_X1 _10656_ ( .A(_03059_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02336_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03060_ ) );
NAND3_X1 _10657_ ( .A1(_03058_ ), .A2(_03060_ ), .A3(_02346_ ), .ZN(_03061_ ) );
MUX2_X1 _10658_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03062_ ) );
MUX2_X1 _10659_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03063_ ) );
MUX2_X1 _10660_ ( .A(_03062_ ), .B(_03063_ ), .S(_02329_ ), .Z(_03064_ ) );
OAI211_X1 _10661_ ( .A(_02324_ ), .B(_03061_ ), .C1(_03064_ ), .C2(_02347_ ), .ZN(_03065_ ) );
NAND2_X1 _10662_ ( .A1(_03056_ ), .A2(_03065_ ), .ZN(_03066_ ) );
OAI21_X2 _10663_ ( .A(_03066_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_03067_ ) );
AND2_X4 _10664_ ( .A1(_03047_ ), .A2(_03067_ ), .ZN(_03068_ ) );
AND2_X1 _10665_ ( .A1(_03068_ ), .A2(\ID_EX_imm [9] ), .ZN(_03069_ ) );
INV_X1 _10666_ ( .A(_03069_ ), .ZN(_03070_ ) );
OR2_X1 _10667_ ( .A1(_03068_ ), .A2(\ID_EX_imm [9] ), .ZN(_03071_ ) );
AND3_X1 _10668_ ( .A1(_03046_ ), .A2(_03070_ ), .A3(_03071_ ), .ZN(_03072_ ) );
NAND2_X1 _10669_ ( .A1(_02459_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_03073_ ) );
NOR2_X1 _10670_ ( .A1(_02337_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03074_ ) );
OAI21_X1 _10671_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_25 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03075_ ) );
NOR2_X1 _10672_ ( .A1(fanout_net_25 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03076_ ) );
OAI21_X1 _10673_ ( .A(_02330_ ), .B1(_02337_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03077_ ) );
OAI221_X1 _10674_ ( .A(_02347_ ), .B1(_03074_ ), .B2(_03075_ ), .C1(_03076_ ), .C2(_03077_ ), .ZN(_03078_ ) );
MUX2_X1 _10675_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03079_ ) );
MUX2_X1 _10676_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03080_ ) );
MUX2_X1 _10677_ ( .A(_03079_ ), .B(_03080_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03081_ ) );
OAI211_X1 _10678_ ( .A(fanout_net_29 ), .B(_03078_ ), .C1(_03081_ ), .C2(_02750_ ), .ZN(_03082_ ) );
OR2_X1 _10679_ ( .A1(fanout_net_25 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03083_ ) );
OAI211_X1 _10680_ ( .A(_03083_ ), .B(_02744_ ), .C1(_02723_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03084_ ) );
OR2_X1 _10681_ ( .A1(fanout_net_25 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03085_ ) );
OAI211_X1 _10682_ ( .A(_03085_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02723_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03086_ ) );
NAND3_X1 _10683_ ( .A1(_03084_ ), .A2(_03086_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03087_ ) );
MUX2_X1 _10684_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03088_ ) );
MUX2_X1 _10685_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03089_ ) );
MUX2_X1 _10686_ ( .A(_03088_ ), .B(_03089_ ), .S(_02330_ ), .Z(_03090_ ) );
OAI211_X1 _10687_ ( .A(_02324_ ), .B(_03087_ ), .C1(_03090_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03091_ ) );
NAND2_X1 _10688_ ( .A1(_03082_ ), .A2(_03091_ ), .ZN(_03092_ ) );
OAI21_X4 _10689_ ( .A(_03092_ ), .B1(_02482_ ), .B2(_02484_ ), .ZN(_03093_ ) );
AND2_X2 _10690_ ( .A1(_03073_ ), .A2(_03093_ ), .ZN(_03094_ ) );
BUF_X8 _10691_ ( .A(_03094_ ), .Z(_03095_ ) );
INV_X1 _10692_ ( .A(\ID_EX_imm [10] ), .ZN(_03096_ ) );
XNOR2_X1 _10693_ ( .A(_03095_ ), .B(_03096_ ), .ZN(_03097_ ) );
NAND2_X1 _10694_ ( .A1(_02458_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03098_ ) );
OR2_X1 _10695_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03099_ ) );
OAI211_X1 _10696_ ( .A(_03099_ ), .B(_02330_ ), .C1(_02337_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03100_ ) );
OR2_X1 _10697_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03101_ ) );
OAI211_X1 _10698_ ( .A(_03101_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02336_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03102_ ) );
NAND3_X1 _10699_ ( .A1(_03100_ ), .A2(_03102_ ), .A3(_02346_ ), .ZN(_03103_ ) );
MUX2_X1 _10700_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03104_ ) );
MUX2_X1 _10701_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03105_ ) );
MUX2_X1 _10702_ ( .A(_03104_ ), .B(_03105_ ), .S(_02329_ ), .Z(_03106_ ) );
OAI211_X1 _10703_ ( .A(fanout_net_29 ), .B(_03103_ ), .C1(_03106_ ), .C2(_02347_ ), .ZN(_03107_ ) );
OR2_X1 _10704_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03108_ ) );
OAI211_X1 _10705_ ( .A(_03108_ ), .B(_02330_ ), .C1(_02337_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03109_ ) );
OR2_X1 _10706_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03110_ ) );
OAI211_X1 _10707_ ( .A(_03110_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02336_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03111_ ) );
NAND3_X1 _10708_ ( .A1(_03109_ ), .A2(_03111_ ), .A3(_02346_ ), .ZN(_03112_ ) );
MUX2_X1 _10709_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03113_ ) );
MUX2_X1 _10710_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03114_ ) );
MUX2_X1 _10711_ ( .A(_03113_ ), .B(_03114_ ), .S(_02329_ ), .Z(_03115_ ) );
OAI211_X1 _10712_ ( .A(_02324_ ), .B(_03112_ ), .C1(_03115_ ), .C2(_02347_ ), .ZN(_03116_ ) );
NAND2_X1 _10713_ ( .A1(_03107_ ), .A2(_03116_ ), .ZN(_03117_ ) );
OAI21_X1 _10714_ ( .A(_03117_ ), .B1(_02456_ ), .B2(_02457_ ), .ZN(_03118_ ) );
AND3_X1 _10715_ ( .A1(_03098_ ), .A2(\ID_EX_imm [11] ), .A3(_03118_ ), .ZN(_03119_ ) );
AOI21_X1 _10716_ ( .A(\ID_EX_imm [11] ), .B1(_03098_ ), .B2(_03118_ ), .ZN(_03120_ ) );
NOR2_X1 _10717_ ( .A1(_03119_ ), .A2(_03120_ ), .ZN(_03121_ ) );
AND2_X1 _10718_ ( .A1(_03097_ ), .A2(_03121_ ), .ZN(_03122_ ) );
AND2_X1 _10719_ ( .A1(_03072_ ), .A2(_03122_ ), .ZN(_03123_ ) );
AND3_X1 _10720_ ( .A1(_02925_ ), .A2(_03022_ ), .A3(_03123_ ), .ZN(_03124_ ) );
INV_X2 _10721_ ( .A(_03124_ ), .ZN(_03125_ ) );
XNOR2_X1 _10722_ ( .A(_03068_ ), .B(\ID_EX_imm [9] ), .ZN(_03126_ ) );
NAND3_X1 _10723_ ( .A1(_03023_ ), .A2(\ID_EX_imm [8] ), .A3(_03043_ ), .ZN(_03127_ ) );
OAI21_X1 _10724_ ( .A(_03070_ ), .B1(_03126_ ), .B2(_03127_ ), .ZN(_03128_ ) );
NAND2_X1 _10725_ ( .A1(_03122_ ), .A2(_03128_ ), .ZN(_03129_ ) );
AND2_X1 _10726_ ( .A1(_03095_ ), .A2(\ID_EX_imm [10] ), .ZN(_03130_ ) );
AOI21_X1 _10727_ ( .A(_03119_ ), .B1(_03130_ ), .B2(_03121_ ), .ZN(_03131_ ) );
AND2_X1 _10728_ ( .A1(_03129_ ), .A2(_03131_ ), .ZN(_03132_ ) );
INV_X1 _10729_ ( .A(_03132_ ), .ZN(_03133_ ) );
AND2_X1 _10730_ ( .A1(_03133_ ), .A2(_03022_ ), .ZN(_03134_ ) );
AND2_X1 _10731_ ( .A1(_02996_ ), .A2(\ID_EX_imm [15] ), .ZN(_03135_ ) );
NAND2_X1 _10732_ ( .A1(_02948_ ), .A2(\ID_EX_imm [12] ), .ZN(_03136_ ) );
AOI21_X1 _10733_ ( .A(_02971_ ), .B1(_03136_ ), .B2(_02973_ ), .ZN(_03137_ ) );
AND3_X1 _10734_ ( .A1(_02997_ ), .A2(_03021_ ), .A3(_03137_ ), .ZN(_03138_ ) );
AND2_X1 _10735_ ( .A1(_03020_ ), .A2(\ID_EX_imm [14] ), .ZN(_03139_ ) );
AND2_X1 _10736_ ( .A1(_02997_ ), .A2(_03139_ ), .ZN(_03140_ ) );
NOR4_X1 _10737_ ( .A1(_03134_ ), .A2(_03135_ ), .A3(_03138_ ), .A4(_03140_ ), .ZN(_03141_ ) );
AOI211_X1 _10738_ ( .A(_02613_ ), .B(_02712_ ), .C1(_03125_ ), .C2(_03141_ ), .ZN(_03142_ ) );
INV_X1 _10739_ ( .A(_03142_ ), .ZN(_03143_ ) );
AND2_X1 _10740_ ( .A1(_02709_ ), .A2(\ID_EX_imm [16] ), .ZN(_03144_ ) );
AND2_X1 _10741_ ( .A1(_02686_ ), .A2(_03144_ ), .ZN(_03145_ ) );
AOI21_X1 _10742_ ( .A(_03145_ ), .B1(\ID_EX_imm [17] ), .B2(_02684_ ), .ZN(_03146_ ) );
INV_X1 _10743_ ( .A(_02637_ ), .ZN(_03147_ ) );
NOR4_X1 _10744_ ( .A1(_03146_ ), .A2(_02659_ ), .A3(_02660_ ), .A4(_03147_ ), .ZN(_03148_ ) );
AND3_X1 _10745_ ( .A1(_02661_ ), .A2(\ID_EX_imm [18] ), .A3(_02635_ ), .ZN(_03149_ ) );
NOR3_X1 _10746_ ( .A1(_03148_ ), .A2(_02659_ ), .A3(_03149_ ), .ZN(_03150_ ) );
NOR2_X1 _10747_ ( .A1(_03150_ ), .A2(_02613_ ), .ZN(_03151_ ) );
AND2_X1 _10748_ ( .A1(_02561_ ), .A2(\ID_EX_imm [23] ), .ZN(_03152_ ) );
NAND2_X1 _10749_ ( .A1(_02610_ ), .A2(\ID_EX_imm [20] ), .ZN(_03153_ ) );
INV_X1 _10750_ ( .A(_02586_ ), .ZN(_03154_ ) );
AOI21_X1 _10751_ ( .A(_02587_ ), .B1(_03153_ ), .B2(_03154_ ), .ZN(_03155_ ) );
AND3_X1 _10752_ ( .A1(_02537_ ), .A2(_03155_ ), .A3(_02563_ ), .ZN(_03156_ ) );
AND2_X1 _10753_ ( .A1(_02535_ ), .A2(\ID_EX_imm [22] ), .ZN(_03157_ ) );
AND2_X1 _10754_ ( .A1(_02563_ ), .A2(_03157_ ), .ZN(_03158_ ) );
NOR4_X1 _10755_ ( .A1(_03151_ ), .A2(_03152_ ), .A3(_03156_ ), .A4(_03158_ ), .ZN(_03159_ ) );
AOI21_X2 _10756_ ( .A(_02513_ ), .B1(_03143_ ), .B2(_03159_ ), .ZN(_03160_ ) );
AOI21_X1 _10757_ ( .A(_02511_ ), .B1(_02490_ ), .B2(_02509_ ), .ZN(_03161_ ) );
NOR2_X1 _10758_ ( .A1(_03160_ ), .A2(_03161_ ), .ZN(_03162_ ) );
OR3_X1 _10759_ ( .A1(_02389_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02396_ ), .ZN(_03163_ ) );
OR2_X1 _10760_ ( .A1(fanout_net_25 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03164_ ) );
OAI211_X1 _10761_ ( .A(_03164_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02342_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03165_ ) );
INV_X1 _10762_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03166_ ) );
NAND2_X1 _10763_ ( .A1(_03166_ ), .A2(fanout_net_25 ), .ZN(_03167_ ) );
OAI211_X1 _10764_ ( .A(_03167_ ), .B(_02335_ ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03168_ ) );
NAND3_X1 _10765_ ( .A1(_03165_ ), .A2(_03168_ ), .A3(_02351_ ), .ZN(_03169_ ) );
MUX2_X1 _10766_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03170_ ) );
MUX2_X1 _10767_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03171_ ) );
MUX2_X1 _10768_ ( .A(_03170_ ), .B(_03171_ ), .S(_02335_ ), .Z(_03172_ ) );
OAI211_X1 _10769_ ( .A(fanout_net_29 ), .B(_03169_ ), .C1(_03172_ ), .C2(_02356_ ), .ZN(_03173_ ) );
OR2_X1 _10770_ ( .A1(fanout_net_25 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03174_ ) );
OAI211_X1 _10771_ ( .A(_03174_ ), .B(_02335_ ), .C1(_02342_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03175_ ) );
OR2_X1 _10772_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03176_ ) );
OAI211_X1 _10773_ ( .A(_03176_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02342_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03177_ ) );
NAND3_X1 _10774_ ( .A1(_03175_ ), .A2(_03177_ ), .A3(_02351_ ), .ZN(_03178_ ) );
MUX2_X1 _10775_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03179_ ) );
MUX2_X1 _10776_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03180_ ) );
MUX2_X1 _10777_ ( .A(_03179_ ), .B(_03180_ ), .S(_02334_ ), .Z(_03181_ ) );
OAI211_X1 _10778_ ( .A(_02327_ ), .B(_03178_ ), .C1(_03181_ ), .C2(_02356_ ), .ZN(_03182_ ) );
OAI211_X1 _10779_ ( .A(_03173_ ), .B(_03182_ ), .C1(_02389_ ), .C2(_02397_ ), .ZN(_03183_ ) );
NAND2_X1 _10780_ ( .A1(_03163_ ), .A2(_03183_ ), .ZN(_03184_ ) );
NAND2_X1 _10781_ ( .A1(_03184_ ), .A2(\ID_EX_imm [25] ), .ZN(_03185_ ) );
NAND2_X1 _10782_ ( .A1(_03162_ ), .A2(_03185_ ), .ZN(_03186_ ) );
OR3_X1 _10783_ ( .A1(_02390_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02397_ ), .ZN(_03187_ ) );
OR2_X1 _10784_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03188_ ) );
OAI211_X1 _10785_ ( .A(_03188_ ), .B(_02405_ ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03189_ ) );
OR2_X1 _10786_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03190_ ) );
OAI211_X1 _10787_ ( .A(_03190_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03191_ ) );
NAND3_X1 _10788_ ( .A1(_03189_ ), .A2(_03191_ ), .A3(_02356_ ), .ZN(_03192_ ) );
MUX2_X1 _10789_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03193_ ) );
MUX2_X1 _10790_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03194_ ) );
MUX2_X1 _10791_ ( .A(_03193_ ), .B(_03194_ ), .S(_02405_ ), .Z(_03195_ ) );
OAI211_X1 _10792_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03192_ ), .C1(_03195_ ), .C2(_02356_ ), .ZN(_03196_ ) );
OR2_X1 _10793_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03197_ ) );
OAI211_X1 _10794_ ( .A(_03197_ ), .B(_02405_ ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03198_ ) );
OR2_X1 _10795_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03199_ ) );
OAI211_X1 _10796_ ( .A(_03199_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03200_ ) );
NAND3_X1 _10797_ ( .A1(_03198_ ), .A2(_03200_ ), .A3(_02356_ ), .ZN(_03201_ ) );
MUX2_X1 _10798_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03202_ ) );
MUX2_X1 _10799_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03203_ ) );
MUX2_X1 _10800_ ( .A(_03202_ ), .B(_03203_ ), .S(_02405_ ), .Z(_03204_ ) );
OAI211_X1 _10801_ ( .A(_02327_ ), .B(_03201_ ), .C1(_03204_ ), .C2(_02356_ ), .ZN(_03205_ ) );
OAI211_X1 _10802_ ( .A(_03196_ ), .B(_03205_ ), .C1(_02390_ ), .C2(_02397_ ), .ZN(_03206_ ) );
NAND2_X2 _10803_ ( .A1(_03187_ ), .A2(_03206_ ), .ZN(_03207_ ) );
INV_X1 _10804_ ( .A(\ID_EX_imm [26] ), .ZN(_03208_ ) );
XNOR2_X1 _10805_ ( .A(_03207_ ), .B(_03208_ ), .ZN(_03209_ ) );
INV_X1 _10806_ ( .A(\ID_EX_imm [25] ), .ZN(_03210_ ) );
NAND3_X1 _10807_ ( .A1(_03163_ ), .A2(_03210_ ), .A3(_03183_ ), .ZN(_03211_ ) );
AND4_X2 _10808_ ( .A1(_02489_ ), .A2(_03186_ ), .A3(_03209_ ), .A4(_03211_ ), .ZN(_03212_ ) );
AND2_X1 _10809_ ( .A1(_03207_ ), .A2(\ID_EX_imm [26] ), .ZN(_03213_ ) );
AND2_X1 _10810_ ( .A1(_03213_ ), .A2(_02489_ ), .ZN(_03214_ ) );
AOI21_X1 _10811_ ( .A(_03214_ ), .B1(\ID_EX_imm [27] ), .B2(_02487_ ), .ZN(_03215_ ) );
INV_X1 _10812_ ( .A(_03215_ ), .ZN(_03216_ ) );
OAI211_X1 _10813_ ( .A(_02427_ ), .B(_02450_ ), .C1(_03212_ ), .C2(_03216_ ), .ZN(_03217_ ) );
AOI21_X1 _10814_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02428_ ), .B2(_02447_ ), .ZN(_03218_ ) );
INV_X1 _10815_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03219_ ) );
AOI22_X1 _10816_ ( .A1(_02427_ ), .A2(_03218_ ), .B1(_03219_ ), .B2(_02425_ ), .ZN(_03220_ ) );
AOI21_X2 _10817_ ( .A(_02403_ ), .B1(_03217_ ), .B2(_03220_ ), .ZN(_03221_ ) );
AOI21_X1 _10818_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02399_ ), .B2(_02400_ ), .ZN(_03222_ ) );
NOR2_X1 _10819_ ( .A1(_03221_ ), .A2(_03222_ ), .ZN(_03223_ ) );
OR2_X1 _10820_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03224_ ) );
OAI211_X1 _10821_ ( .A(_03224_ ), .B(_02405_ ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03225_ ) );
OR2_X1 _10822_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03226_ ) );
OAI211_X1 _10823_ ( .A(_03226_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02406_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03227_ ) );
NAND3_X1 _10824_ ( .A1(_03225_ ), .A2(_03227_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03228_ ) );
MUX2_X1 _10825_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03229_ ) );
MUX2_X1 _10826_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03230_ ) );
MUX2_X1 _10827_ ( .A(_03229_ ), .B(_03230_ ), .S(_02335_ ), .Z(_03231_ ) );
OAI211_X1 _10828_ ( .A(_02327_ ), .B(_03228_ ), .C1(_03231_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03232_ ) );
MUX2_X1 _10829_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03233_ ) );
AND2_X1 _10830_ ( .A1(_03233_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_03234_ ) );
MUX2_X1 _10831_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03235_ ) );
AOI211_X1 _10832_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_03234_ ), .C1(_02405_ ), .C2(_03235_ ), .ZN(_03236_ ) );
MUX2_X1 _10833_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03237_ ) );
MUX2_X1 _10834_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03238_ ) );
MUX2_X1 _10835_ ( .A(_03237_ ), .B(_03238_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03239_ ) );
OAI21_X1 _10836_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B1(_03239_ ), .B2(_02356_ ), .ZN(_03240_ ) );
OAI221_X1 _10837_ ( .A(_03232_ ), .B1(_03236_ ), .B2(_03240_ ), .C1(_02390_ ), .C2(_02397_ ), .ZN(_03241_ ) );
OR3_X1 _10838_ ( .A1(_02389_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02396_ ), .ZN(_03242_ ) );
NAND2_X1 _10839_ ( .A1(_03241_ ), .A2(_03242_ ), .ZN(_03243_ ) );
XNOR2_X1 _10840_ ( .A(_03243_ ), .B(\ID_EX_imm [31] ), .ZN(_03244_ ) );
XNOR2_X1 _10841_ ( .A(_03223_ ), .B(_03244_ ), .ZN(_03245_ ) );
AND2_X2 _10842_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_03246_ ) );
BUF_X4 _10843_ ( .A(_03246_ ), .Z(_03247_ ) );
BUF_X4 _10844_ ( .A(_03247_ ), .Z(_03248_ ) );
NOR2_X1 _10845_ ( .A1(_03245_ ), .A2(_03248_ ), .ZN(_00133_ ) );
AND3_X1 _10846_ ( .A1(_03217_ ), .A2(_03220_ ), .A3(_02403_ ), .ZN(_03249_ ) );
NOR3_X1 _10847_ ( .A1(_03249_ ), .A2(_03221_ ), .A3(_03247_ ), .ZN(_00134_ ) );
AOI21_X1 _10848_ ( .A(_02712_ ), .B1(_03125_ ), .B2(_03141_ ), .ZN(_03250_ ) );
INV_X1 _10849_ ( .A(_03150_ ), .ZN(_03251_ ) );
OAI21_X1 _10850_ ( .A(_02611_ ), .B1(_03250_ ), .B2(_03251_ ), .ZN(_03252_ ) );
NAND2_X1 _10851_ ( .A1(_03252_ ), .A2(_03153_ ), .ZN(_03253_ ) );
XNOR2_X1 _10852_ ( .A(_03253_ ), .B(_02588_ ), .ZN(_03254_ ) );
NOR2_X1 _10853_ ( .A1(_03254_ ), .A2(_03248_ ), .ZN(_00135_ ) );
OR3_X1 _10854_ ( .A1(_03250_ ), .A2(_02611_ ), .A3(_03251_ ), .ZN(_03255_ ) );
INV_X1 _10855_ ( .A(_03246_ ), .ZN(_03256_ ) );
BUF_X2 _10856_ ( .A(_03256_ ), .Z(_03257_ ) );
AND3_X1 _10857_ ( .A1(_03255_ ), .A2(_03257_ ), .A3(_03252_ ), .ZN(_00136_ ) );
INV_X1 _10858_ ( .A(_02711_ ), .ZN(_03258_ ) );
AOI21_X1 _10859_ ( .A(_03258_ ), .B1(_03125_ ), .B2(_03141_ ), .ZN(_03259_ ) );
AND2_X1 _10860_ ( .A1(_03259_ ), .A2(_02686_ ), .ZN(_03260_ ) );
INV_X1 _10861_ ( .A(_03260_ ), .ZN(_03261_ ) );
AOI21_X1 _10862_ ( .A(_03147_ ), .B1(_03261_ ), .B2(_03146_ ), .ZN(_03262_ ) );
AND2_X1 _10863_ ( .A1(_02635_ ), .A2(\ID_EX_imm [18] ), .ZN(_03263_ ) );
OR2_X1 _10864_ ( .A1(_03262_ ), .A2(_03263_ ), .ZN(_03264_ ) );
XNOR2_X1 _10865_ ( .A(_03264_ ), .B(_02661_ ), .ZN(_03265_ ) );
NOR2_X1 _10866_ ( .A1(_03265_ ), .A2(_03248_ ), .ZN(_00137_ ) );
AND3_X1 _10867_ ( .A1(_03261_ ), .A2(_03147_ ), .A3(_03146_ ), .ZN(_03266_ ) );
NOR3_X1 _10868_ ( .A1(_03266_ ), .A2(_03262_ ), .A3(_03247_ ), .ZN(_00138_ ) );
OR2_X1 _10869_ ( .A1(_03259_ ), .A2(_03144_ ), .ZN(_03267_ ) );
XNOR2_X1 _10870_ ( .A(_03267_ ), .B(_02686_ ), .ZN(_03268_ ) );
NOR2_X1 _10871_ ( .A1(_03268_ ), .A2(_03248_ ), .ZN(_00139_ ) );
AND3_X1 _10872_ ( .A1(_03125_ ), .A2(_03141_ ), .A3(_03258_ ), .ZN(_03269_ ) );
NOR3_X1 _10873_ ( .A1(_03269_ ), .A2(_03259_ ), .A3(_03247_ ), .ZN(_00140_ ) );
NAND2_X1 _10874_ ( .A1(_02972_ ), .A2(_02973_ ), .ZN(_03270_ ) );
INV_X1 _10875_ ( .A(_02949_ ), .ZN(_03271_ ) );
NAND2_X1 _10876_ ( .A1(_02925_ ), .A2(_03123_ ), .ZN(_03272_ ) );
AOI211_X1 _10877_ ( .A(_03270_ ), .B(_03271_ ), .C1(_03272_ ), .C2(_03132_ ), .ZN(_03273_ ) );
OR2_X1 _10878_ ( .A1(_03273_ ), .A2(_03137_ ), .ZN(_03274_ ) );
AND2_X1 _10879_ ( .A1(_03274_ ), .A2(_03021_ ), .ZN(_03275_ ) );
OR2_X1 _10880_ ( .A1(_03275_ ), .A2(_03139_ ), .ZN(_03276_ ) );
XNOR2_X1 _10881_ ( .A(_03276_ ), .B(_02997_ ), .ZN(_03277_ ) );
NOR2_X1 _10882_ ( .A1(_03277_ ), .A2(_03248_ ), .ZN(_00141_ ) );
XOR2_X1 _10883_ ( .A(_03274_ ), .B(_03021_ ), .Z(_03278_ ) );
AND2_X1 _10884_ ( .A1(_03278_ ), .A2(_03257_ ), .ZN(_00142_ ) );
NAND2_X1 _10885_ ( .A1(_03272_ ), .A2(_03132_ ), .ZN(_03279_ ) );
NAND2_X1 _10886_ ( .A1(_03279_ ), .A2(_02949_ ), .ZN(_03280_ ) );
AND2_X1 _10887_ ( .A1(_03280_ ), .A2(_03136_ ), .ZN(_03281_ ) );
XNOR2_X1 _10888_ ( .A(_03281_ ), .B(_03270_ ), .ZN(_03282_ ) );
NOR2_X1 _10889_ ( .A1(_03282_ ), .A2(_03248_ ), .ZN(_00143_ ) );
XNOR2_X1 _10890_ ( .A(_03279_ ), .B(_03271_ ), .ZN(_03283_ ) );
AND2_X1 _10891_ ( .A1(_03283_ ), .A2(_03257_ ), .ZN(_00144_ ) );
NOR2_X1 _10892_ ( .A1(_03212_ ), .A2(_03216_ ), .ZN(_03284_ ) );
NOR2_X1 _10893_ ( .A1(_03284_ ), .A2(_02449_ ), .ZN(_03285_ ) );
OR2_X2 _10894_ ( .A1(_03285_ ), .A2(_03218_ ), .ZN(_03286_ ) );
XNOR2_X1 _10895_ ( .A(_03286_ ), .B(_02427_ ), .ZN(_03287_ ) );
NOR2_X1 _10896_ ( .A1(_03287_ ), .A2(_03248_ ), .ZN(_00145_ ) );
XNOR2_X1 _10897_ ( .A(_03284_ ), .B(_02450_ ), .ZN(_03288_ ) );
AND2_X1 _10898_ ( .A1(_03288_ ), .A2(_03257_ ), .ZN(_00146_ ) );
AND3_X1 _10899_ ( .A1(_03186_ ), .A2(_03209_ ), .A3(_03211_ ), .ZN(_03289_ ) );
OR2_X1 _10900_ ( .A1(_03289_ ), .A2(_03213_ ), .ZN(_03290_ ) );
XNOR2_X1 _10901_ ( .A(_03290_ ), .B(_02489_ ), .ZN(_03291_ ) );
NOR2_X1 _10902_ ( .A1(_03291_ ), .A2(_03248_ ), .ZN(_00147_ ) );
AOI21_X1 _10903_ ( .A(_03209_ ), .B1(_03186_ ), .B2(_03211_ ), .ZN(_03292_ ) );
NOR3_X1 _10904_ ( .A1(_03289_ ), .A2(_03292_ ), .A3(_03247_ ), .ZN(_00148_ ) );
NAND2_X1 _10905_ ( .A1(_03185_ ), .A2(_03211_ ), .ZN(_03293_ ) );
XNOR2_X1 _10906_ ( .A(_03162_ ), .B(_03293_ ), .ZN(_03294_ ) );
NOR2_X1 _10907_ ( .A1(_03294_ ), .A2(_03248_ ), .ZN(_00149_ ) );
AND3_X1 _10908_ ( .A1(_03143_ ), .A2(_03159_ ), .A3(_02513_ ), .ZN(_03295_ ) );
NOR3_X1 _10909_ ( .A1(_03295_ ), .A2(_03160_ ), .A3(_03247_ ), .ZN(_00150_ ) );
AND2_X1 _10910_ ( .A1(_02611_ ), .A2(_02588_ ), .ZN(_03296_ ) );
OAI21_X1 _10911_ ( .A(_03296_ ), .B1(_03250_ ), .B2(_03251_ ), .ZN(_03297_ ) );
INV_X1 _10912_ ( .A(_03297_ ), .ZN(_03298_ ) );
OR2_X1 _10913_ ( .A1(_03298_ ), .A2(_03155_ ), .ZN(_03299_ ) );
AND2_X1 _10914_ ( .A1(_03299_ ), .A2(_02537_ ), .ZN(_03300_ ) );
OR2_X1 _10915_ ( .A1(_03300_ ), .A2(_03157_ ), .ZN(_03301_ ) );
XNOR2_X1 _10916_ ( .A(_03301_ ), .B(_02563_ ), .ZN(_03302_ ) );
NOR2_X1 _10917_ ( .A1(_03302_ ), .A2(_03248_ ), .ZN(_00151_ ) );
XOR2_X1 _10918_ ( .A(_03299_ ), .B(_02537_ ), .Z(_03303_ ) );
AND2_X1 _10919_ ( .A1(_03303_ ), .A2(_03257_ ), .ZN(_00152_ ) );
INV_X1 _10920_ ( .A(\IF_ID_inst [6] ), .ZN(_03304_ ) );
NOR2_X1 _10921_ ( .A1(_03304_ ), .A2(\IF_ID_inst [12] ), .ZN(_03305_ ) );
AND2_X1 _10922_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03306_ ) );
BUF_X2 _10923_ ( .A(_03306_ ), .Z(_03307_ ) );
AND3_X1 _10924_ ( .A1(_03305_ ), .A2(\IF_ID_inst [13] ), .A3(_03307_ ), .ZN(_03308_ ) );
AND2_X2 _10925_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_03309_ ) );
NOR2_X1 _10926_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_03310_ ) );
AND2_X1 _10927_ ( .A1(_03309_ ), .A2(_03310_ ), .ZN(_03311_ ) );
BUF_X2 _10928_ ( .A(_03311_ ), .Z(_03312_ ) );
CLKBUF_X2 _10929_ ( .A(_03312_ ), .Z(_03313_ ) );
AND2_X1 _10930_ ( .A1(_03308_ ), .A2(_03313_ ), .ZN(_03314_ ) );
AND4_X1 _10931_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03315_ ) );
AND2_X1 _10932_ ( .A1(_03313_ ), .A2(_03315_ ), .ZN(_03316_ ) );
NOR2_X2 _10933_ ( .A1(_03314_ ), .A2(_03316_ ), .ZN(_03317_ ) );
BUF_X4 _10934_ ( .A(_03317_ ), .Z(_03318_ ) );
INV_X1 _10935_ ( .A(\IF_ID_inst [31] ), .ZN(_03319_ ) );
NOR2_X1 _10936_ ( .A1(fanout_net_4 ), .A2(fanout_net_17 ), .ZN(_03320_ ) );
AND2_X2 _10937_ ( .A1(_02312_ ), .A2(_03320_ ), .ZN(_03321_ ) );
INV_X2 _10938_ ( .A(_03321_ ), .ZN(_03322_ ) );
BUF_X4 _10939_ ( .A(_03322_ ), .Z(_03323_ ) );
NOR3_X1 _10940_ ( .A1(_03318_ ), .A2(_03319_ ), .A3(_03323_ ), .ZN(_00231_ ) );
INV_X1 _10941_ ( .A(\IF_ID_inst [30] ), .ZN(_03324_ ) );
NOR3_X1 _10942_ ( .A1(_03318_ ), .A2(_03324_ ), .A3(_03323_ ), .ZN(_00232_ ) );
INV_X1 _10943_ ( .A(\IF_ID_inst [21] ), .ZN(_03325_ ) );
NOR3_X1 _10944_ ( .A1(_03318_ ), .A2(_03325_ ), .A3(_03323_ ), .ZN(_00233_ ) );
BUF_X4 _10945_ ( .A(_03322_ ), .Z(_03326_ ) );
INV_X1 _10946_ ( .A(_03317_ ), .ZN(_03327_ ) );
INV_X1 _10947_ ( .A(\IF_ID_inst [20] ), .ZN(_03328_ ) );
AOI21_X1 _10948_ ( .A(_03326_ ), .B1(_03327_ ), .B2(_03328_ ), .ZN(_00234_ ) );
INV_X1 _10949_ ( .A(\IF_ID_inst [29] ), .ZN(_03329_ ) );
AOI21_X1 _10950_ ( .A(_03326_ ), .B1(_03327_ ), .B2(_03329_ ), .ZN(_00235_ ) );
INV_X1 _10951_ ( .A(\IF_ID_inst [28] ), .ZN(_03330_ ) );
AOI21_X1 _10952_ ( .A(_03326_ ), .B1(_03327_ ), .B2(_03330_ ), .ZN(_00236_ ) );
INV_X1 _10953_ ( .A(\IF_ID_inst [27] ), .ZN(_03331_ ) );
NOR3_X1 _10954_ ( .A1(_03318_ ), .A2(_03331_ ), .A3(_03323_ ), .ZN(_00237_ ) );
INV_X1 _10955_ ( .A(\IF_ID_inst [26] ), .ZN(_03332_ ) );
AOI21_X1 _10956_ ( .A(_03326_ ), .B1(_03327_ ), .B2(_03332_ ), .ZN(_00238_ ) );
INV_X1 _10957_ ( .A(\IF_ID_inst [25] ), .ZN(_03333_ ) );
BUF_X4 _10958_ ( .A(_03322_ ), .Z(_03334_ ) );
NOR3_X1 _10959_ ( .A1(_03318_ ), .A2(_03333_ ), .A3(_03334_ ), .ZN(_00239_ ) );
INV_X1 _10960_ ( .A(\IF_ID_inst [24] ), .ZN(_03335_ ) );
NOR3_X1 _10961_ ( .A1(_03318_ ), .A2(_03335_ ), .A3(_03334_ ), .ZN(_00240_ ) );
INV_X1 _10962_ ( .A(\IF_ID_inst [23] ), .ZN(_03336_ ) );
NOR3_X1 _10963_ ( .A1(_03318_ ), .A2(_03336_ ), .A3(_03334_ ), .ZN(_00241_ ) );
INV_X1 _10964_ ( .A(\IF_ID_inst [22] ), .ZN(_03337_ ) );
NOR3_X1 _10965_ ( .A1(_03318_ ), .A2(_03337_ ), .A3(_03334_ ), .ZN(_00242_ ) );
BUF_X2 _10966_ ( .A(_03320_ ), .Z(_03338_ ) );
AND3_X1 _10967_ ( .A1(_02312_ ), .A2(_03338_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00243_ ) );
AND3_X1 _10968_ ( .A1(_02312_ ), .A2(_03338_ ), .A3(\myidu.state [2] ), .ZN(_00244_ ) );
INV_X1 _10969_ ( .A(\IF_ID_inst [5] ), .ZN(_03339_ ) );
NOR2_X2 _10970_ ( .A1(_03339_ ), .A2(\IF_ID_inst [4] ), .ZN(_03340_ ) );
NOR2_X1 _10971_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03341_ ) );
AND3_X1 _10972_ ( .A1(_03312_ ), .A2(_03340_ ), .A3(_03341_ ), .ZN(_03342_ ) );
NOR2_X1 _10973_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03343_ ) );
BUF_X2 _10974_ ( .A(_03343_ ), .Z(_03344_ ) );
AND2_X1 _10975_ ( .A1(_03342_ ), .A2(_03344_ ), .ZN(_03345_ ) );
INV_X1 _10976_ ( .A(\IF_ID_inst [12] ), .ZN(_03346_ ) );
NOR2_X1 _10977_ ( .A1(_03346_ ), .A2(\IF_ID_inst [6] ), .ZN(_03347_ ) );
AND3_X1 _10978_ ( .A1(_03313_ ), .A2(_03340_ ), .A3(_03347_ ), .ZN(_03348_ ) );
AND2_X1 _10979_ ( .A1(_03348_ ), .A2(_03344_ ), .ZN(_03349_ ) );
NOR2_X1 _10980_ ( .A1(_03345_ ), .A2(_03349_ ), .ZN(_03350_ ) );
AND2_X1 _10981_ ( .A1(_03305_ ), .A2(_03340_ ), .ZN(_03351_ ) );
AND2_X1 _10982_ ( .A1(_03351_ ), .A2(_03313_ ), .ZN(_03352_ ) );
INV_X1 _10983_ ( .A(\IF_ID_inst [13] ), .ZN(_03353_ ) );
NOR2_X1 _10984_ ( .A1(_03353_ ), .A2(\IF_ID_inst [14] ), .ZN(_03354_ ) );
AOI22_X1 _10985_ ( .A1(_03344_ ), .A2(_03352_ ), .B1(_03342_ ), .B2(_03354_ ), .ZN(_03355_ ) );
NAND2_X1 _10986_ ( .A1(_03350_ ), .A2(_03355_ ), .ZN(_03356_ ) );
INV_X1 _10987_ ( .A(\IF_ID_inst [4] ), .ZN(_03357_ ) );
AND4_X1 _10988_ ( .A1(_03357_ ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03358_ ) );
AND2_X1 _10989_ ( .A1(_03313_ ), .A2(_03358_ ), .ZN(_03359_ ) );
AOI221_X4 _10990_ ( .A(_03356_ ), .B1(\IF_ID_inst [14] ), .B2(_03352_ ), .C1(_03353_ ), .C2(_03359_ ), .ZN(_03360_ ) );
BUF_X2 _10991_ ( .A(_03321_ ), .Z(_03361_ ) );
INV_X1 _10992_ ( .A(\IF_ID_inst [7] ), .ZN(_03362_ ) );
AND4_X1 _10993_ ( .A1(\IF_ID_inst [6] ), .A2(_03313_ ), .A3(_03362_ ), .A4(_03306_ ), .ZN(_03363_ ) );
OR3_X1 _10994_ ( .A1(\IF_ID_inst [11] ), .A2(\IF_ID_inst [10] ), .A3(\IF_ID_inst [9] ), .ZN(_03364_ ) );
NOR2_X1 _10995_ ( .A1(_03364_ ), .A2(\IF_ID_inst [8] ), .ZN(_03365_ ) );
NOR4_X1 _10996_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_03366_ ) );
AND3_X1 _10997_ ( .A1(_03363_ ), .A2(_03365_ ), .A3(_03366_ ), .ZN(_03367_ ) );
NAND2_X1 _10998_ ( .A1(\IF_ID_inst [29] ), .A2(\IF_ID_inst [28] ), .ZN(_03368_ ) );
NOR3_X1 _10999_ ( .A1(_03368_ ), .A2(\IF_ID_inst [30] ), .A3(\IF_ID_inst [31] ), .ZN(_03369_ ) );
NOR3_X1 _11000_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .A3(\IF_ID_inst [24] ), .ZN(_03370_ ) );
AND3_X1 _11001_ ( .A1(_03369_ ), .A2(_03331_ ), .A3(_03370_ ), .ZN(_03371_ ) );
NOR2_X1 _11002_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [18] ), .ZN(_03372_ ) );
NOR2_X1 _11003_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_03373_ ) );
AND2_X1 _11004_ ( .A1(_03372_ ), .A2(_03373_ ), .ZN(_03374_ ) );
NOR2_X1 _11005_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_03375_ ) );
AND3_X1 _11006_ ( .A1(_03375_ ), .A2(\IF_ID_inst [21] ), .A3(_03328_ ), .ZN(_03376_ ) );
AND3_X1 _11007_ ( .A1(_03371_ ), .A2(_03374_ ), .A3(_03376_ ), .ZN(_03377_ ) );
AND2_X1 _11008_ ( .A1(_03367_ ), .A2(_03377_ ), .ZN(_03378_ ) );
NAND2_X1 _11009_ ( .A1(_03370_ ), .A2(_03331_ ), .ZN(_03379_ ) );
NAND4_X1 _11010_ ( .A1(_03324_ ), .A2(_03329_ ), .A3(_03330_ ), .A4(_03319_ ), .ZN(_03380_ ) );
NOR2_X1 _11011_ ( .A1(_03379_ ), .A2(_03380_ ), .ZN(_03381_ ) );
AND3_X1 _11012_ ( .A1(_03372_ ), .A2(_03373_ ), .A3(_03375_ ), .ZN(_03382_ ) );
AND4_X1 _11013_ ( .A1(_03325_ ), .A2(_03381_ ), .A3(\IF_ID_inst [20] ), .A4(_03382_ ), .ZN(_03383_ ) );
AND2_X1 _11014_ ( .A1(_03367_ ), .A2(_03383_ ), .ZN(_03384_ ) );
AND2_X2 _11015_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03385_ ) );
AND2_X1 _11016_ ( .A1(_03359_ ), .A2(_03385_ ), .ZN(_03386_ ) );
AND3_X1 _11017_ ( .A1(_03309_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_03387_ ) );
NOR2_X1 _11018_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03388_ ) );
AND3_X1 _11019_ ( .A1(_03388_ ), .A2(\IF_ID_inst [12] ), .A3(_03304_ ), .ZN(_03389_ ) );
NAND2_X1 _11020_ ( .A1(_03387_ ), .A2(_03389_ ), .ZN(_03390_ ) );
INV_X1 _11021_ ( .A(_03344_ ), .ZN(_03391_ ) );
NOR2_X1 _11022_ ( .A1(_03390_ ), .A2(_03391_ ), .ZN(_03392_ ) );
NOR4_X1 _11023_ ( .A1(_03378_ ), .A2(_03384_ ), .A3(_03386_ ), .A4(_03392_ ), .ZN(_03393_ ) );
AND4_X1 _11024_ ( .A1(\IF_ID_inst [11] ), .A2(_03360_ ), .A3(_03361_ ), .A4(_03393_ ), .ZN(_00245_ ) );
AND4_X1 _11025_ ( .A1(\IF_ID_inst [10] ), .A2(_03360_ ), .A3(_03361_ ), .A4(_03393_ ), .ZN(_00246_ ) );
AND4_X1 _11026_ ( .A1(\IF_ID_inst [9] ), .A2(_03360_ ), .A3(_03321_ ), .A4(_03393_ ), .ZN(_00247_ ) );
AND4_X1 _11027_ ( .A1(\IF_ID_inst [8] ), .A2(_03360_ ), .A3(_03321_ ), .A4(_03393_ ), .ZN(_00248_ ) );
AND4_X1 _11028_ ( .A1(\IF_ID_inst [7] ), .A2(_03360_ ), .A3(_03321_ ), .A4(_03393_ ), .ZN(_00249_ ) );
OR2_X2 _11029_ ( .A1(_03384_ ), .A2(_03392_ ), .ZN(_03394_ ) );
INV_X1 _11030_ ( .A(\IF_ID_inst [19] ), .ZN(_03395_ ) );
INV_X1 _11031_ ( .A(\IF_ID_inst [2] ), .ZN(_03396_ ) );
NOR2_X1 _11032_ ( .A1(_03396_ ), .A2(\IF_ID_inst [3] ), .ZN(_03397_ ) );
AND2_X1 _11033_ ( .A1(_03397_ ), .A2(_03309_ ), .ZN(_03398_ ) );
NOR2_X1 _11034_ ( .A1(_03357_ ), .A2(\IF_ID_inst [6] ), .ZN(_03399_ ) );
AND2_X1 _11035_ ( .A1(_03398_ ), .A2(_03399_ ), .ZN(_03400_ ) );
INV_X1 _11036_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03401_ ) );
AND2_X1 _11037_ ( .A1(_03340_ ), .A2(_03401_ ), .ZN(_03402_ ) );
AND2_X4 _11038_ ( .A1(_03402_ ), .A2(_03387_ ), .ZN(_03403_ ) );
CLKBUF_X2 _11039_ ( .A(_03403_ ), .Z(_03404_ ) );
BUF_X2 _11040_ ( .A(_03404_ ), .Z(_03405_ ) );
NOR2_X1 _11041_ ( .A1(_03400_ ), .A2(_03405_ ), .ZN(_03406_ ) );
NAND3_X1 _11042_ ( .A1(_03376_ ), .A2(_03374_ ), .A3(_03369_ ), .ZN(_03407_ ) );
NOR2_X1 _11043_ ( .A1(_03407_ ), .A2(_03379_ ), .ZN(_03408_ ) );
INV_X1 _11044_ ( .A(_03408_ ), .ZN(_03409_ ) );
INV_X1 _11045_ ( .A(\IF_ID_inst [15] ), .ZN(_03410_ ) );
AND4_X1 _11046_ ( .A1(\IF_ID_inst [4] ), .A2(_03362_ ), .A3(_03410_ ), .A4(\IF_ID_inst [5] ), .ZN(_03411_ ) );
AND3_X1 _11047_ ( .A1(_03411_ ), .A2(_03305_ ), .A3(_03343_ ), .ZN(_03412_ ) );
BUF_X2 _11048_ ( .A(_03313_ ), .Z(_03413_ ) );
NAND3_X1 _11049_ ( .A1(_03412_ ), .A2(_03413_ ), .A3(_03365_ ), .ZN(_03414_ ) );
OAI21_X1 _11050_ ( .A(_03406_ ), .B1(_03409_ ), .B2(_03414_ ), .ZN(_03415_ ) );
NOR4_X1 _11051_ ( .A1(_03394_ ), .A2(_03395_ ), .A3(_03334_ ), .A4(_03415_ ), .ZN(_00250_ ) );
INV_X1 _11052_ ( .A(\IF_ID_inst [18] ), .ZN(_03416_ ) );
NOR4_X1 _11053_ ( .A1(_03394_ ), .A2(_03416_ ), .A3(_03334_ ), .A4(_03415_ ), .ZN(_00251_ ) );
INV_X1 _11054_ ( .A(\IF_ID_inst [17] ), .ZN(_03417_ ) );
NOR4_X1 _11055_ ( .A1(_03394_ ), .A2(_03417_ ), .A3(_03334_ ), .A4(_03415_ ), .ZN(_00252_ ) );
NOR2_X1 _11056_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_03418_ ) );
AND3_X1 _11057_ ( .A1(_03385_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_03418_ ), .ZN(_03419_ ) );
NOR3_X1 _11058_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_03420_ ) );
AND3_X1 _11059_ ( .A1(_03419_ ), .A2(_03331_ ), .A3(_03420_ ), .ZN(_03421_ ) );
AND2_X1 _11060_ ( .A1(_03312_ ), .A2(_03341_ ), .ZN(_03422_ ) );
BUF_X2 _11061_ ( .A(_03422_ ), .Z(_03423_ ) );
NAND3_X1 _11062_ ( .A1(_03421_ ), .A2(_03307_ ), .A3(_03423_ ), .ZN(_03424_ ) );
AND3_X1 _11063_ ( .A1(_03309_ ), .A2(\IF_ID_inst [12] ), .A3(_03310_ ), .ZN(_03425_ ) );
AND3_X1 _11064_ ( .A1(_03304_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_03426_ ) );
AND2_X1 _11065_ ( .A1(_03425_ ), .A2(_03426_ ), .ZN(_03427_ ) );
NAND2_X1 _11066_ ( .A1(_03421_ ), .A2(_03427_ ), .ZN(_03428_ ) );
NAND2_X1 _11067_ ( .A1(_03424_ ), .A2(_03428_ ), .ZN(_03429_ ) );
AND3_X1 _11068_ ( .A1(_03420_ ), .A2(_03331_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03430_ ) );
INV_X1 _11069_ ( .A(\IF_ID_inst [14] ), .ZN(_03431_ ) );
NOR2_X1 _11070_ ( .A1(_03431_ ), .A2(\IF_ID_inst [13] ), .ZN(_03432_ ) );
AND2_X1 _11071_ ( .A1(_03432_ ), .A2(_03418_ ), .ZN(_03433_ ) );
AND2_X1 _11072_ ( .A1(_03430_ ), .A2(_03433_ ), .ZN(_03434_ ) );
AND3_X1 _11073_ ( .A1(_03434_ ), .A2(_03307_ ), .A3(_03422_ ), .ZN(_03435_ ) );
AND2_X2 _11074_ ( .A1(_03343_ ), .A2(_03418_ ), .ZN(_03436_ ) );
AND4_X1 _11075_ ( .A1(_03307_ ), .A2(_03422_ ), .A3(_03430_ ), .A4(_03436_ ), .ZN(_03437_ ) );
NOR3_X1 _11076_ ( .A1(_03429_ ), .A2(_03435_ ), .A3(_03437_ ), .ZN(_03438_ ) );
INV_X1 _11077_ ( .A(_03438_ ), .ZN(_03439_ ) );
AND2_X2 _11078_ ( .A1(_03420_ ), .A2(_03331_ ), .ZN(_03440_ ) );
AND4_X1 _11079_ ( .A1(_03431_ ), .A2(_03418_ ), .A3(\IF_ID_inst [13] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03441_ ) );
AND2_X1 _11080_ ( .A1(_03440_ ), .A2(_03441_ ), .ZN(_03442_ ) );
AND3_X1 _11081_ ( .A1(_03343_ ), .A2(_03418_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03443_ ) );
AND2_X1 _11082_ ( .A1(_03440_ ), .A2(_03443_ ), .ZN(_03444_ ) );
AND4_X1 _11083_ ( .A1(\IF_ID_inst [14] ), .A2(_03418_ ), .A3(_03353_ ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03445_ ) );
AND2_X1 _11084_ ( .A1(_03440_ ), .A2(_03445_ ), .ZN(_03446_ ) );
NOR3_X1 _11085_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(_03446_ ), .ZN(_03447_ ) );
INV_X1 _11086_ ( .A(_03447_ ), .ZN(_03448_ ) );
AND2_X1 _11087_ ( .A1(_03448_ ), .A2(_03427_ ), .ZN(_03449_ ) );
NOR2_X1 _11088_ ( .A1(_03324_ ), .A2(\IF_ID_inst [29] ), .ZN(_03450_ ) );
NOR2_X1 _11089_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_03451_ ) );
AND3_X1 _11090_ ( .A1(_03450_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_03451_ ), .ZN(_03452_ ) );
AND2_X1 _11091_ ( .A1(_03452_ ), .A2(_03433_ ), .ZN(_03453_ ) );
AND2_X1 _11092_ ( .A1(_03453_ ), .A2(_03427_ ), .ZN(_03454_ ) );
NOR3_X1 _11093_ ( .A1(_03439_ ), .A2(_03449_ ), .A3(_03454_ ), .ZN(_03455_ ) );
NOR2_X1 _11094_ ( .A1(_03357_ ), .A2(\IF_ID_inst [5] ), .ZN(_03456_ ) );
AND2_X1 _11095_ ( .A1(_03422_ ), .A2(_03456_ ), .ZN(_03457_ ) );
INV_X1 _11096_ ( .A(_03354_ ), .ZN(_03458_ ) );
NAND2_X1 _11097_ ( .A1(_03457_ ), .A2(_03458_ ), .ZN(_03459_ ) );
AND4_X2 _11098_ ( .A1(\IF_ID_inst [4] ), .A2(_03339_ ), .A3(_03304_ ), .A4(\IF_ID_inst [12] ), .ZN(_03460_ ) );
AND2_X2 _11099_ ( .A1(_03312_ ), .A2(_03460_ ), .ZN(_03461_ ) );
AND2_X1 _11100_ ( .A1(_03461_ ), .A2(_03354_ ), .ZN(_03462_ ) );
INV_X1 _11101_ ( .A(_03462_ ), .ZN(_03463_ ) );
INV_X1 _11102_ ( .A(_03385_ ), .ZN(_03464_ ) );
NAND3_X1 _11103_ ( .A1(_03422_ ), .A2(_03464_ ), .A3(_03388_ ), .ZN(_03465_ ) );
NAND3_X1 _11104_ ( .A1(_03461_ ), .A2(\IF_ID_inst [14] ), .A3(\IF_ID_inst [13] ), .ZN(_03466_ ) );
NAND4_X1 _11105_ ( .A1(_03459_ ), .A2(_03463_ ), .A3(_03465_ ), .A4(_03466_ ), .ZN(_03467_ ) );
NAND2_X1 _11106_ ( .A1(_03457_ ), .A2(_03354_ ), .ZN(_03468_ ) );
AND3_X1 _11107_ ( .A1(_03305_ ), .A2(_03340_ ), .A3(_03343_ ), .ZN(_03469_ ) );
AND2_X1 _11108_ ( .A1(_03469_ ), .A2(_03398_ ), .ZN(_03470_ ) );
INV_X1 _11109_ ( .A(_03470_ ), .ZN(_03471_ ) );
AND2_X1 _11110_ ( .A1(_03389_ ), .A2(_03313_ ), .ZN(_03472_ ) );
NAND2_X1 _11111_ ( .A1(_03472_ ), .A2(_03353_ ), .ZN(_03473_ ) );
NAND3_X1 _11112_ ( .A1(_03468_ ), .A2(_03471_ ), .A3(_03473_ ), .ZN(_03474_ ) );
NOR2_X2 _11113_ ( .A1(_03467_ ), .A2(_03474_ ), .ZN(_03475_ ) );
AND2_X1 _11114_ ( .A1(_03475_ ), .A2(_03317_ ), .ZN(_03476_ ) );
AND2_X1 _11115_ ( .A1(_03342_ ), .A2(_03354_ ), .ZN(_03477_ ) );
INV_X1 _11116_ ( .A(_03477_ ), .ZN(_03478_ ) );
OAI21_X1 _11117_ ( .A(_03343_ ), .B1(_03342_ ), .B2(_03348_ ), .ZN(_03479_ ) );
AND2_X1 _11118_ ( .A1(_03478_ ), .A2(_03479_ ), .ZN(_03480_ ) );
INV_X2 _11119_ ( .A(_03480_ ), .ZN(_03481_ ) );
OR2_X1 _11120_ ( .A1(_03352_ ), .A2(_03359_ ), .ZN(_03482_ ) );
AND2_X1 _11121_ ( .A1(_03482_ ), .A2(_03458_ ), .ZN(_03483_ ) );
OAI21_X1 _11122_ ( .A(_03461_ ), .B1(_03434_ ), .B2(_03453_ ), .ZN(_03484_ ) );
NAND3_X1 _11123_ ( .A1(_03442_ ), .A2(_03307_ ), .A3(_03423_ ), .ZN(_03485_ ) );
NAND4_X1 _11124_ ( .A1(_03423_ ), .A2(_03307_ ), .A3(_03452_ ), .A4(_03436_ ), .ZN(_03486_ ) );
NAND3_X1 _11125_ ( .A1(_03461_ ), .A2(_03430_ ), .A3(_03436_ ), .ZN(_03487_ ) );
NAND4_X1 _11126_ ( .A1(_03484_ ), .A2(_03485_ ), .A3(_03486_ ), .A4(_03487_ ), .ZN(_03488_ ) );
NOR3_X1 _11127_ ( .A1(_03481_ ), .A2(_03483_ ), .A3(_03488_ ), .ZN(_03489_ ) );
AND3_X1 _11128_ ( .A1(_03455_ ), .A2(_03476_ ), .A3(_03489_ ), .ZN(_03490_ ) );
NOR2_X1 _11129_ ( .A1(_03394_ ), .A2(_03415_ ), .ZN(_03491_ ) );
AND2_X1 _11130_ ( .A1(_03490_ ), .A2(_03491_ ), .ZN(_03492_ ) );
INV_X1 _11131_ ( .A(_03492_ ), .ZN(_03493_ ) );
XNOR2_X1 _11132_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_03494_ ) );
XNOR2_X1 _11133_ ( .A(\myexu.pc_jump [2] ), .B(\IF_ID_pc [2] ), .ZN(_03495_ ) );
XNOR2_X1 _11134_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_03496_ ) );
XNOR2_X1 _11135_ ( .A(fanout_net_9 ), .B(\myexu.pc_jump [3] ), .ZN(_03497_ ) );
AND4_X1 _11136_ ( .A1(_03494_ ), .A2(_03495_ ), .A3(_03496_ ), .A4(_03497_ ), .ZN(_03498_ ) );
XNOR2_X1 _11137_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_03499_ ) );
XNOR2_X1 _11138_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_03500_ ) );
XNOR2_X1 _11139_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_03501_ ) );
XNOR2_X1 _11140_ ( .A(fanout_net_13 ), .B(\myexu.pc_jump [4] ), .ZN(_03502_ ) );
AND4_X1 _11141_ ( .A1(_03499_ ), .A2(_03500_ ), .A3(_03501_ ), .A4(_03502_ ), .ZN(_03503_ ) );
XNOR2_X1 _11142_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_03504_ ) );
XNOR2_X1 _11143_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_03505_ ) );
XNOR2_X1 _11144_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_03506_ ) );
XNOR2_X1 _11145_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_03507_ ) );
AND4_X1 _11146_ ( .A1(_03504_ ), .A2(_03505_ ), .A3(_03506_ ), .A4(_03507_ ), .ZN(_03508_ ) );
XNOR2_X1 _11147_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_03509_ ) );
XNOR2_X1 _11148_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_03510_ ) );
XNOR2_X1 _11149_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_03511_ ) );
XNOR2_X1 _11150_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_03512_ ) );
AND4_X1 _11151_ ( .A1(_03509_ ), .A2(_03510_ ), .A3(_03511_ ), .A4(_03512_ ), .ZN(_03513_ ) );
AND4_X1 _11152_ ( .A1(_03498_ ), .A2(_03503_ ), .A3(_03508_ ), .A4(_03513_ ), .ZN(_03514_ ) );
XNOR2_X1 _11153_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_03515_ ) );
XNOR2_X1 _11154_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_03516_ ) );
XNOR2_X1 _11155_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_03517_ ) );
XNOR2_X1 _11156_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_03518_ ) );
AND4_X1 _11157_ ( .A1(_03515_ ), .A2(_03516_ ), .A3(_03517_ ), .A4(_03518_ ), .ZN(_03519_ ) );
XNOR2_X1 _11158_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_03520_ ) );
XNOR2_X1 _11159_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_03521_ ) );
XNOR2_X1 _11160_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_03522_ ) );
XNOR2_X1 _11161_ ( .A(\IF_ID_pc [25] ), .B(\myexu.pc_jump [25] ), .ZN(_03523_ ) );
AND4_X1 _11162_ ( .A1(_03520_ ), .A2(_03521_ ), .A3(_03522_ ), .A4(_03523_ ), .ZN(_03524_ ) );
XNOR2_X1 _11163_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_03525_ ) );
XNOR2_X1 _11164_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_03526_ ) );
XNOR2_X1 _11165_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_03527_ ) );
XNOR2_X1 _11166_ ( .A(\IF_ID_pc [21] ), .B(\myexu.pc_jump [21] ), .ZN(_03528_ ) );
AND4_X1 _11167_ ( .A1(_03525_ ), .A2(_03526_ ), .A3(_03527_ ), .A4(_03528_ ), .ZN(_03529_ ) );
XNOR2_X1 _11168_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_03530_ ) );
XNOR2_X1 _11169_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_03531_ ) );
XNOR2_X1 _11170_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_03532_ ) );
XNOR2_X1 _11171_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_03533_ ) );
AND4_X1 _11172_ ( .A1(_03530_ ), .A2(_03531_ ), .A3(_03532_ ), .A4(_03533_ ), .ZN(_03534_ ) );
AND4_X1 _11173_ ( .A1(_03519_ ), .A2(_03524_ ), .A3(_03529_ ), .A4(_03534_ ), .ZN(_03535_ ) );
AND2_X1 _11174_ ( .A1(_03514_ ), .A2(_03535_ ), .ZN(_03536_ ) );
INV_X1 _11175_ ( .A(check_quest ), .ZN(_03537_ ) );
NOR2_X1 _11176_ ( .A1(_03536_ ), .A2(_03537_ ), .ZN(_03538_ ) );
INV_X1 _11177_ ( .A(\myifu.state [1] ), .ZN(_03539_ ) );
NOR2_X1 _11178_ ( .A1(_03539_ ), .A2(\myifu.to_reset ), .ZN(_03540_ ) );
INV_X1 _11179_ ( .A(_03540_ ), .ZN(_03541_ ) );
NOR2_X1 _11180_ ( .A1(_03538_ ), .A2(_03541_ ), .ZN(_03542_ ) );
AND2_X1 _11181_ ( .A1(_03542_ ), .A2(IDU_ready_IFU ), .ZN(_03543_ ) );
NAND4_X1 _11182_ ( .A1(_03493_ ), .A2(\IF_ID_inst [18] ), .A3(_03491_ ), .A4(_03543_ ), .ZN(_03544_ ) );
BUF_X4 _11183_ ( .A(_03492_ ), .Z(_03545_ ) );
INV_X1 _11184_ ( .A(_03543_ ), .ZN(_03546_ ) );
BUF_X4 _11185_ ( .A(_03546_ ), .Z(_03547_ ) );
OAI21_X1 _11186_ ( .A(\ID_EX_rs1 [3] ), .B1(_03545_ ), .B2(_03547_ ), .ZN(_03548_ ) );
AOI21_X1 _11187_ ( .A(_03326_ ), .B1(_03544_ ), .B2(_03548_ ), .ZN(_00253_ ) );
INV_X1 _11188_ ( .A(\IF_ID_inst [16] ), .ZN(_03549_ ) );
NOR4_X1 _11189_ ( .A1(_03394_ ), .A2(_03549_ ), .A3(_03334_ ), .A4(_03415_ ), .ZN(_00254_ ) );
NAND4_X1 _11190_ ( .A1(_03493_ ), .A2(\IF_ID_inst [17] ), .A3(_03491_ ), .A4(_03543_ ), .ZN(_03550_ ) );
OAI21_X1 _11191_ ( .A(\ID_EX_rs1 [2] ), .B1(_03545_ ), .B2(_03547_ ), .ZN(_03551_ ) );
AOI21_X1 _11192_ ( .A(_03326_ ), .B1(_03550_ ), .B2(_03551_ ), .ZN(_00255_ ) );
NOR4_X1 _11193_ ( .A1(_03394_ ), .A2(_03410_ ), .A3(_03334_ ), .A4(_03415_ ), .ZN(_00256_ ) );
NOR2_X1 _11194_ ( .A1(_03492_ ), .A2(_03546_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OAI21_X1 _11195_ ( .A(_03321_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [1] ), .ZN(_03552_ ) );
OR3_X1 _11196_ ( .A1(_03394_ ), .A2(_03549_ ), .A3(_03415_ ), .ZN(_03553_ ) );
AOI21_X1 _11197_ ( .A(_03552_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(_03553_ ), .ZN(_00257_ ) );
AND4_X1 _11198_ ( .A1(_03313_ ), .A2(_03440_ ), .A3(_03433_ ), .A4(_03460_ ), .ZN(_03554_ ) );
NAND2_X1 _11199_ ( .A1(_03554_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03555_ ) );
AND4_X1 _11200_ ( .A1(_03313_ ), .A2(_03440_ ), .A3(_03436_ ), .A4(_03460_ ), .ZN(_03556_ ) );
NAND2_X1 _11201_ ( .A1(_03556_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03557_ ) );
NAND3_X1 _11202_ ( .A1(_03423_ ), .A2(_03432_ ), .A3(_03456_ ), .ZN(_03558_ ) );
NAND4_X1 _11203_ ( .A1(_03463_ ), .A2(_03555_ ), .A3(_03557_ ), .A4(_03558_ ), .ZN(_03559_ ) );
NAND3_X1 _11204_ ( .A1(_03423_ ), .A2(_03385_ ), .A3(_03456_ ), .ZN(_03560_ ) );
NAND3_X1 _11205_ ( .A1(_03413_ ), .A2(_03460_ ), .A3(_03385_ ), .ZN(_03561_ ) );
NAND2_X1 _11206_ ( .A1(_03560_ ), .A2(_03561_ ), .ZN(_03562_ ) );
AND2_X1 _11207_ ( .A1(_03457_ ), .A2(_03344_ ), .ZN(_03563_ ) );
OR4_X1 _11208_ ( .A1(_03405_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03563_ ), .ZN(_03564_ ) );
NAND3_X1 _11209_ ( .A1(_03423_ ), .A2(_03353_ ), .A3(_03388_ ), .ZN(_03565_ ) );
NAND2_X1 _11210_ ( .A1(_03565_ ), .A2(_03473_ ), .ZN(_03566_ ) );
AND4_X1 _11211_ ( .A1(_03433_ ), .A2(_03461_ ), .A3(_03450_ ), .A4(_03451_ ), .ZN(_03567_ ) );
NAND2_X1 _11212_ ( .A1(_03567_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03568_ ) );
NAND2_X1 _11213_ ( .A1(_03568_ ), .A2(_03468_ ), .ZN(_03569_ ) );
OR4_X2 _11214_ ( .A1(_03400_ ), .A2(_03564_ ), .A3(_03566_ ), .A4(_03569_ ), .ZN(_03570_ ) );
AND2_X1 _11215_ ( .A1(_03423_ ), .A2(_03388_ ), .ZN(_03571_ ) );
AND2_X1 _11216_ ( .A1(_03571_ ), .A2(_03354_ ), .ZN(_03572_ ) );
NAND4_X1 _11217_ ( .A1(_03305_ ), .A2(_03340_ ), .A3(_03397_ ), .A4(_03309_ ), .ZN(_03573_ ) );
NOR2_X1 _11218_ ( .A1(_03573_ ), .A2(_03391_ ), .ZN(_03574_ ) );
NOR4_X1 _11219_ ( .A1(_03378_ ), .A2(_03572_ ), .A3(_03392_ ), .A4(_03574_ ), .ZN(_03575_ ) );
INV_X1 _11220_ ( .A(_03314_ ), .ZN(_03576_ ) );
NAND3_X1 _11221_ ( .A1(_03413_ ), .A2(_03353_ ), .A3(_03315_ ), .ZN(_03577_ ) );
INV_X1 _11222_ ( .A(_03384_ ), .ZN(_03578_ ) );
NAND4_X1 _11223_ ( .A1(_03315_ ), .A2(_03309_ ), .A3(_03310_ ), .A4(_03354_ ), .ZN(_03579_ ) );
NAND3_X1 _11224_ ( .A1(_03413_ ), .A2(_03315_ ), .A3(_03385_ ), .ZN(_03580_ ) );
AND3_X1 _11225_ ( .A1(_03578_ ), .A2(_03579_ ), .A3(_03580_ ), .ZN(_03581_ ) );
NAND4_X1 _11226_ ( .A1(_03575_ ), .A2(_03576_ ), .A3(_03577_ ), .A4(_03581_ ), .ZN(_03582_ ) );
NOR4_X1 _11227_ ( .A1(_03570_ ), .A2(_03335_ ), .A3(_03334_ ), .A4(_03582_ ), .ZN(_00258_ ) );
AOI211_X1 _11228_ ( .A(_03547_ ), .B(_03545_ ), .C1(\IF_ID_inst [15] ), .C2(_03491_ ), .ZN(_03583_ ) );
AOI21_X1 _11229_ ( .A(\ID_EX_rs1 [0] ), .B1(_03493_ ), .B2(_03543_ ), .ZN(_03584_ ) );
NOR3_X1 _11230_ ( .A1(_03583_ ), .A2(_03326_ ), .A3(_03584_ ), .ZN(_00259_ ) );
NOR4_X1 _11231_ ( .A1(_03570_ ), .A2(_03336_ ), .A3(_03322_ ), .A4(_03582_ ), .ZN(_00260_ ) );
NOR4_X1 _11232_ ( .A1(_03570_ ), .A2(_03337_ ), .A3(_03322_ ), .A4(_03582_ ), .ZN(_00261_ ) );
NOR2_X1 _11233_ ( .A1(_03570_ ), .A2(_03582_ ), .ZN(_03585_ ) );
AOI211_X1 _11234_ ( .A(_03545_ ), .B(_03547_ ), .C1(_03585_ ), .C2(\IF_ID_inst [23] ), .ZN(_03586_ ) );
OAI21_X1 _11235_ ( .A(_03361_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs2 [3] ), .ZN(_03587_ ) );
NOR2_X1 _11236_ ( .A1(_03586_ ), .A2(_03587_ ), .ZN(_00262_ ) );
NOR4_X1 _11237_ ( .A1(_03570_ ), .A2(_03325_ ), .A3(_03322_ ), .A4(_03582_ ), .ZN(_00263_ ) );
AOI211_X1 _11238_ ( .A(_03545_ ), .B(_03547_ ), .C1(_03585_ ), .C2(\IF_ID_inst [22] ), .ZN(_03588_ ) );
AOI21_X1 _11239_ ( .A(\ID_EX_rs2 [2] ), .B1(_03493_ ), .B2(_03543_ ), .ZN(_03589_ ) );
NOR3_X1 _11240_ ( .A1(_03588_ ), .A2(_03326_ ), .A3(_03589_ ), .ZN(_00264_ ) );
NOR4_X1 _11241_ ( .A1(_03570_ ), .A2(_03328_ ), .A3(_03322_ ), .A4(_03582_ ), .ZN(_00265_ ) );
AOI211_X1 _11242_ ( .A(_03545_ ), .B(_03547_ ), .C1(_03585_ ), .C2(\IF_ID_inst [21] ), .ZN(_03590_ ) );
OAI21_X1 _11243_ ( .A(_03361_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs2 [1] ), .ZN(_03591_ ) );
NOR2_X1 _11244_ ( .A1(_03590_ ), .A2(_03591_ ), .ZN(_00266_ ) );
INV_X1 _11245_ ( .A(IDU_valid_EXU ), .ZN(_03592_ ) );
AND4_X1 _11246_ ( .A1(\IF_ID_inst [12] ), .A2(_03344_ ), .A3(_03388_ ), .A4(_03304_ ), .ZN(_03593_ ) );
AND4_X1 _11247_ ( .A1(_03592_ ), .A2(_03593_ ), .A3(_03321_ ), .A4(_03387_ ), .ZN(_00267_ ) );
AOI211_X1 _11248_ ( .A(_03545_ ), .B(_03547_ ), .C1(_03585_ ), .C2(\IF_ID_inst [20] ), .ZN(_03594_ ) );
OAI21_X1 _11249_ ( .A(_03361_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs2 [0] ), .ZN(_03595_ ) );
NOR2_X1 _11250_ ( .A1(_03594_ ), .A2(_03595_ ), .ZN(_00268_ ) );
INV_X1 _11251_ ( .A(_03475_ ), .ZN(_03596_ ) );
XNOR2_X1 _11252_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_03597_ ) );
XNOR2_X1 _11253_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_03598_ ) );
XNOR2_X1 _11254_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_03599_ ) );
XNOR2_X1 _11255_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_03600_ ) );
AND4_X1 _11256_ ( .A1(_03597_ ), .A2(_03598_ ), .A3(_03599_ ), .A4(_03600_ ), .ZN(_03601_ ) );
XNOR2_X1 _11257_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_03602_ ) );
AND2_X1 _11258_ ( .A1(_03601_ ), .A2(_03602_ ), .ZN(_03603_ ) );
AND2_X1 _11259_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03604_ ) );
INV_X1 _11260_ ( .A(\ID_EX_typ [7] ), .ZN(_03605_ ) );
AND2_X1 _11261_ ( .A1(_03604_ ), .A2(_03605_ ), .ZN(_03606_ ) );
AND2_X1 _11262_ ( .A1(_03603_ ), .A2(_03606_ ), .ZN(_03607_ ) );
XNOR2_X1 _11263_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_03608_ ) );
XNOR2_X1 _11264_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_03609_ ) );
XNOR2_X1 _11265_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_03610_ ) );
NAND4_X1 _11266_ ( .A1(_03606_ ), .A2(_03608_ ), .A3(_03609_ ), .A4(_03610_ ), .ZN(_03611_ ) );
XOR2_X1 _11267_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .Z(_03612_ ) );
XOR2_X1 _11268_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .Z(_03613_ ) );
NOR3_X1 _11269_ ( .A1(_03611_ ), .A2(_03612_ ), .A3(_03613_ ), .ZN(_03614_ ) );
OR2_X1 _11270_ ( .A1(_03607_ ), .A2(_03614_ ), .ZN(_03615_ ) );
AOI211_X1 _11271_ ( .A(_03327_ ), .B(_03596_ ), .C1(_03491_ ), .C2(_03615_ ), .ZN(_03616_ ) );
INV_X1 _11272_ ( .A(IDU_ready_IFU ), .ZN(_03617_ ) );
AOI21_X1 _11273_ ( .A(_03607_ ), .B1(_03475_ ), .B2(_03317_ ), .ZN(_03618_ ) );
NOR4_X1 _11274_ ( .A1(_03616_ ), .A2(_03617_ ), .A3(_03322_ ), .A4(_03618_ ), .ZN(_00269_ ) );
BUF_X4 _11275_ ( .A(_03483_ ), .Z(_03619_ ) );
NAND4_X1 _11276_ ( .A1(_03412_ ), .A2(_03328_ ), .A3(_03413_ ), .A4(_03365_ ), .ZN(_03620_ ) );
NAND3_X1 _11277_ ( .A1(_03381_ ), .A2(_03325_ ), .A3(_03382_ ), .ZN(_03621_ ) );
NOR2_X1 _11278_ ( .A1(_03620_ ), .A2(_03621_ ), .ZN(_03622_ ) );
NOR2_X1 _11279_ ( .A1(_03405_ ), .A2(_03574_ ), .ZN(_03623_ ) );
INV_X1 _11280_ ( .A(_03623_ ), .ZN(_03624_ ) );
NOR4_X1 _11281_ ( .A1(_03619_ ), .A2(_03327_ ), .A3(_03622_ ), .A4(_03624_ ), .ZN(_03625_ ) );
AND2_X1 _11282_ ( .A1(_03593_ ), .A2(_03387_ ), .ZN(_03626_ ) );
INV_X1 _11283_ ( .A(_03414_ ), .ZN(_03627_ ) );
AOI21_X1 _11284_ ( .A(_03626_ ), .B1(_03627_ ), .B2(_03408_ ), .ZN(_03628_ ) );
AOI21_X1 _11285_ ( .A(_03326_ ), .B1(_03625_ ), .B2(_03628_ ), .ZN(_00270_ ) );
NAND2_X1 _11286_ ( .A1(_03472_ ), .A2(_03432_ ), .ZN(_03629_ ) );
NAND2_X1 _11287_ ( .A1(_03472_ ), .A2(_03344_ ), .ZN(_03630_ ) );
AND4_X1 _11288_ ( .A1(_03480_ ), .A2(_03629_ ), .A3(_03630_ ), .A4(_03465_ ), .ZN(_03631_ ) );
NOR2_X1 _11289_ ( .A1(_03622_ ), .A2(_03327_ ), .ZN(_03632_ ) );
AOI21_X1 _11290_ ( .A(_03326_ ), .B1(_03631_ ), .B2(_03632_ ), .ZN(_00271_ ) );
NAND3_X1 _11291_ ( .A1(_03446_ ), .A2(_03307_ ), .A3(_03423_ ), .ZN(_03633_ ) );
NAND4_X1 _11292_ ( .A1(_03423_ ), .A2(_03307_ ), .A3(_03440_ ), .A4(_03443_ ), .ZN(_03634_ ) );
NAND2_X1 _11293_ ( .A1(_03633_ ), .A2(_03634_ ), .ZN(_03635_ ) );
AND3_X1 _11294_ ( .A1(_03307_ ), .A2(_03309_ ), .A3(_03310_ ), .ZN(_03636_ ) );
AND2_X1 _11295_ ( .A1(_03636_ ), .A2(_03347_ ), .ZN(_03637_ ) );
AOI21_X1 _11296_ ( .A(_03635_ ), .B1(_03448_ ), .B2(_03637_ ), .ZN(_03638_ ) );
AND4_X1 _11297_ ( .A1(_03331_ ), .A2(_03420_ ), .A3(_03385_ ), .A4(_03418_ ), .ZN(_03639_ ) );
AND2_X1 _11298_ ( .A1(_03423_ ), .A2(_03307_ ), .ZN(_03640_ ) );
OAI211_X1 _11299_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B(_03639_ ), .C1(_03640_ ), .C2(_03637_ ), .ZN(_03641_ ) );
AND3_X1 _11300_ ( .A1(_03456_ ), .A2(_03309_ ), .A3(_03310_ ), .ZN(_03642_ ) );
NAND3_X1 _11301_ ( .A1(_03642_ ), .A2(\IF_ID_inst [13] ), .A3(_03347_ ), .ZN(_03643_ ) );
NAND4_X1 _11302_ ( .A1(_03638_ ), .A2(_03641_ ), .A3(_03459_ ), .A4(_03643_ ), .ZN(_03644_ ) );
NAND4_X1 _11303_ ( .A1(_03413_ ), .A2(_03411_ ), .A3(_03305_ ), .A4(_03344_ ), .ZN(_03645_ ) );
NOR4_X1 _11304_ ( .A1(_03645_ ), .A2(\IF_ID_inst [20] ), .A3(\IF_ID_inst [8] ), .A4(_03364_ ), .ZN(_03646_ ) );
AND3_X1 _11305_ ( .A1(_03381_ ), .A2(_03325_ ), .A3(_03382_ ), .ZN(_03647_ ) );
NAND2_X1 _11306_ ( .A1(_03646_ ), .A2(_03647_ ), .ZN(_03648_ ) );
AND2_X1 _11307_ ( .A1(_03453_ ), .A2(_03637_ ), .ZN(_03649_ ) );
INV_X1 _11308_ ( .A(_03649_ ), .ZN(_03650_ ) );
NAND2_X1 _11309_ ( .A1(_03648_ ), .A2(_03650_ ), .ZN(_03651_ ) );
AND2_X1 _11310_ ( .A1(_03452_ ), .A2(_03436_ ), .ZN(_03652_ ) );
OR2_X1 _11311_ ( .A1(_03652_ ), .A2(_03442_ ), .ZN(_03653_ ) );
AND2_X1 _11312_ ( .A1(_03653_ ), .A2(_03640_ ), .ZN(_03654_ ) );
OR3_X1 _11313_ ( .A1(_03654_ ), .A2(_03572_ ), .A3(_03624_ ), .ZN(_03655_ ) );
NOR4_X1 _11314_ ( .A1(_03644_ ), .A2(_03566_ ), .A3(_03651_ ), .A4(_03655_ ), .ZN(_03656_ ) );
NAND4_X1 _11315_ ( .A1(_03440_ ), .A2(_03433_ ), .A3(_03413_ ), .A4(_03460_ ), .ZN(_03657_ ) );
INV_X1 _11316_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03658_ ) );
NOR2_X1 _11317_ ( .A1(_03657_ ), .A2(_03658_ ), .ZN(_03659_ ) );
NAND4_X1 _11318_ ( .A1(_03440_ ), .A2(_03413_ ), .A3(_03436_ ), .A4(_03460_ ), .ZN(_03660_ ) );
NOR2_X1 _11319_ ( .A1(_03660_ ), .A2(_03658_ ), .ZN(_03661_ ) );
NOR2_X1 _11320_ ( .A1(_03659_ ), .A2(_03661_ ), .ZN(_03662_ ) );
NAND3_X1 _11321_ ( .A1(_03568_ ), .A2(_03662_ ), .A3(_03468_ ), .ZN(_03663_ ) );
NOR2_X1 _11322_ ( .A1(_03663_ ), .A2(_03400_ ), .ZN(_03664_ ) );
AOI21_X1 _11323_ ( .A(_03323_ ), .B1(_03656_ ), .B2(_03664_ ), .ZN(_00272_ ) );
AOI221_X4 _11324_ ( .A(_03626_ ), .B1(\IF_ID_inst [13] ), .B2(_03461_ ), .C1(_03457_ ), .C2(_03458_ ), .ZN(_03665_ ) );
AOI21_X1 _11325_ ( .A(_03323_ ), .B1(_03664_ ), .B2(_03665_ ), .ZN(_00273_ ) );
AOI22_X1 _11326_ ( .A1(_03653_ ), .A2(_03640_ ), .B1(_03627_ ), .B2(_03408_ ), .ZN(_03666_ ) );
INV_X1 _11327_ ( .A(_03400_ ), .ZN(_03667_ ) );
AND3_X1 _11328_ ( .A1(_03666_ ), .A2(_03667_ ), .A3(_03468_ ), .ZN(_03668_ ) );
AOI21_X1 _11329_ ( .A(_03323_ ), .B1(_03668_ ), .B2(_03478_ ), .ZN(_00274_ ) );
AOI21_X1 _11330_ ( .A(_03649_ ), .B1(_03448_ ), .B2(_03637_ ), .ZN(_03669_ ) );
AND3_X1 _11331_ ( .A1(_03642_ ), .A2(_03354_ ), .A3(_03347_ ), .ZN(_03670_ ) );
AOI21_X1 _11332_ ( .A(_03670_ ), .B1(_03571_ ), .B2(_03354_ ), .ZN(_03671_ ) );
AND4_X1 _11333_ ( .A1(_03478_ ), .A2(_03669_ ), .A3(_03667_ ), .A4(_03671_ ), .ZN(_03672_ ) );
NAND3_X1 _11334_ ( .A1(_03453_ ), .A2(_03347_ ), .A3(_03642_ ), .ZN(_03673_ ) );
NAND3_X1 _11335_ ( .A1(_03444_ ), .A2(_03347_ ), .A3(_03642_ ), .ZN(_03674_ ) );
NAND4_X1 _11336_ ( .A1(_03642_ ), .A2(_03440_ ), .A3(_03445_ ), .A4(_03347_ ), .ZN(_03675_ ) );
NAND3_X1 _11337_ ( .A1(_03673_ ), .A2(_03674_ ), .A3(_03675_ ), .ZN(_03676_ ) );
AOI221_X4 _11338_ ( .A(_03676_ ), .B1(\IF_ID_inst [14] ), .B2(_03359_ ), .C1(\IF_ID_inst [13] ), .C2(_03316_ ), .ZN(_03677_ ) );
AOI21_X1 _11339_ ( .A(_03323_ ), .B1(_03672_ ), .B2(_03677_ ), .ZN(_00275_ ) );
INV_X1 _11340_ ( .A(_03349_ ), .ZN(_03678_ ) );
AOI221_X4 _11341_ ( .A(_03314_ ), .B1(_03342_ ), .B2(_03354_ ), .C1(\IF_ID_inst [14] ), .C2(_03352_ ), .ZN(_03679_ ) );
INV_X1 _11342_ ( .A(_03435_ ), .ZN(_03680_ ) );
AOI22_X1 _11343_ ( .A1(_03472_ ), .A2(_03344_ ), .B1(_03398_ ), .B2(_03426_ ), .ZN(_03681_ ) );
AND4_X1 _11344_ ( .A1(_03678_ ), .A2(_03679_ ), .A3(_03680_ ), .A4(_03681_ ), .ZN(_03682_ ) );
AND2_X1 _11345_ ( .A1(_03457_ ), .A2(\IF_ID_inst [14] ), .ZN(_03683_ ) );
INV_X1 _11346_ ( .A(_03683_ ), .ZN(_03684_ ) );
OAI22_X1 _11347_ ( .A1(_03434_ ), .A2(_03453_ ), .B1(_03427_ ), .B2(_03461_ ), .ZN(_03685_ ) );
AOI22_X1 _11348_ ( .A1(_03640_ ), .A2(_03421_ ), .B1(_03432_ ), .B2(_03472_ ), .ZN(_03686_ ) );
AND3_X1 _11349_ ( .A1(_03684_ ), .A2(_03685_ ), .A3(_03686_ ), .ZN(_03687_ ) );
AOI21_X1 _11350_ ( .A(_03323_ ), .B1(_03682_ ), .B2(_03687_ ), .ZN(_00276_ ) );
AND3_X1 _11351_ ( .A1(_03412_ ), .A2(_03413_ ), .A3(_03365_ ), .ZN(_03688_ ) );
AND2_X1 _11352_ ( .A1(_03688_ ), .A2(_03381_ ), .ZN(_03689_ ) );
AND3_X1 _11353_ ( .A1(_03382_ ), .A2(_03325_ ), .A3(\IF_ID_inst [20] ), .ZN(_03690_ ) );
NAND2_X1 _11354_ ( .A1(_03689_ ), .A2(_03690_ ), .ZN(_03691_ ) );
NAND3_X1 _11355_ ( .A1(_03691_ ), .A2(_03478_ ), .A3(_03471_ ), .ZN(_03692_ ) );
AOI21_X1 _11356_ ( .A(_03431_ ), .B1(_03576_ ), .B2(_03577_ ), .ZN(_03693_ ) );
NAND3_X1 _11357_ ( .A1(_03457_ ), .A2(\IF_ID_inst [14] ), .A3(_03353_ ), .ZN(_03694_ ) );
AND2_X1 _11358_ ( .A1(_03430_ ), .A2(_03436_ ), .ZN(_03695_ ) );
AOI22_X1 _11359_ ( .A1(_03695_ ), .A2(_03427_ ), .B1(_03344_ ), .B2(_03359_ ), .ZN(_03696_ ) );
NAND3_X1 _11360_ ( .A1(_03680_ ), .A2(_03694_ ), .A3(_03696_ ), .ZN(_03697_ ) );
NAND2_X1 _11361_ ( .A1(_03479_ ), .A2(_03487_ ), .ZN(_03698_ ) );
NOR4_X1 _11362_ ( .A1(_03692_ ), .A2(_03693_ ), .A3(_03697_ ), .A4(_03698_ ), .ZN(_03699_ ) );
INV_X1 _11363_ ( .A(_03386_ ), .ZN(_03700_ ) );
INV_X1 _11364_ ( .A(_03454_ ), .ZN(_03701_ ) );
AND4_X1 _11365_ ( .A1(_03701_ ), .A2(_03428_ ), .A3(_03485_ ), .A4(_03466_ ), .ZN(_03702_ ) );
NAND4_X1 _11366_ ( .A1(_03452_ ), .A2(_03433_ ), .A3(_03413_ ), .A4(_03460_ ), .ZN(_03703_ ) );
NAND2_X1 _11367_ ( .A1(_03629_ ), .A2(_03703_ ), .ZN(_03704_ ) );
AOI21_X1 _11368_ ( .A(_03704_ ), .B1(_03432_ ), .B2(_03571_ ), .ZN(_03705_ ) );
OAI21_X1 _11369_ ( .A(_03385_ ), .B1(_03352_ ), .B2(_03316_ ), .ZN(_03706_ ) );
AND4_X1 _11370_ ( .A1(_03700_ ), .A2(_03702_ ), .A3(_03705_ ), .A4(_03706_ ), .ZN(_03707_ ) );
AOI21_X1 _11371_ ( .A(_03323_ ), .B1(_03699_ ), .B2(_03707_ ), .ZN(_00277_ ) );
INV_X1 _11372_ ( .A(_03536_ ), .ZN(_03708_ ) );
INV_X1 _11373_ ( .A(\myifu.to_reset ), .ZN(_03709_ ) );
BUF_X4 _11374_ ( .A(_03709_ ), .Z(_03710_ ) );
NAND4_X1 _11375_ ( .A1(_03708_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_03710_ ), .ZN(_03711_ ) );
NAND2_X1 _11376_ ( .A1(\mtvec [0] ), .A2(\myifu.to_reset ), .ZN(_03712_ ) );
AOI21_X1 _11377_ ( .A(fanout_net_4 ), .B1(_03711_ ), .B2(_03712_ ), .ZN(_00281_ ) );
AND4_X1 _11378_ ( .A1(\IF_ID_inst [31] ), .A2(_03357_ ), .A3(_03401_ ), .A4(\IF_ID_inst [5] ), .ZN(_03713_ ) );
AND2_X2 _11379_ ( .A1(_03312_ ), .A2(_03713_ ), .ZN(_03714_ ) );
AOI21_X1 _11380_ ( .A(_03714_ ), .B1(_03405_ ), .B2(\IF_ID_inst [31] ), .ZN(_03715_ ) );
AND2_X1 _11381_ ( .A1(_03714_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03716_ ) );
NOR2_X1 _11382_ ( .A1(_03715_ ), .A2(_03716_ ), .ZN(_03717_ ) );
BUF_X4 _11383_ ( .A(_03717_ ), .Z(_03718_ ) );
XNOR2_X1 _11384_ ( .A(_03718_ ), .B(_02004_ ), .ZN(_03719_ ) );
XOR2_X1 _11385_ ( .A(_03718_ ), .B(\IF_ID_pc [24] ), .Z(_03720_ ) );
XOR2_X1 _11386_ ( .A(_03717_ ), .B(\IF_ID_pc [20] ), .Z(_03721_ ) );
NAND4_X1 _11387_ ( .A1(_03340_ ), .A2(_03401_ ), .A3(_03309_ ), .A4(_03310_ ), .ZN(_03722_ ) );
NOR2_X1 _11388_ ( .A1(_03722_ ), .A2(_03319_ ), .ZN(_03723_ ) );
AND2_X1 _11389_ ( .A1(_03723_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03724_ ) );
INV_X1 _11390_ ( .A(_03724_ ), .ZN(_03725_ ) );
AND2_X1 _11391_ ( .A1(_03405_ ), .A2(\IF_ID_inst [19] ), .ZN(_03726_ ) );
OAI21_X1 _11392_ ( .A(_03725_ ), .B1(_03726_ ), .B2(_03723_ ), .ZN(_03727_ ) );
XNOR2_X1 _11393_ ( .A(_03727_ ), .B(\IF_ID_pc [19] ), .ZN(_03728_ ) );
AND2_X1 _11394_ ( .A1(_03721_ ), .A2(_03728_ ), .ZN(_03729_ ) );
AND2_X1 _11395_ ( .A1(_03405_ ), .A2(\IF_ID_inst [17] ), .ZN(_03730_ ) );
INV_X1 _11396_ ( .A(_03714_ ), .ZN(_03731_ ) );
MUX2_X1 _11397_ ( .A(_03658_ ), .B(_03730_ ), .S(_03731_ ), .Z(_03732_ ) );
XOR2_X1 _11398_ ( .A(_03732_ ), .B(\IF_ID_pc [17] ), .Z(_03733_ ) );
AND2_X1 _11399_ ( .A1(_03404_ ), .A2(\IF_ID_inst [18] ), .ZN(_03734_ ) );
INV_X1 _11400_ ( .A(_03734_ ), .ZN(_03735_ ) );
INV_X1 _11401_ ( .A(_03723_ ), .ZN(_03736_ ) );
AOI21_X1 _11402_ ( .A(_03724_ ), .B1(_03735_ ), .B2(_03736_ ), .ZN(_03737_ ) );
XOR2_X1 _11403_ ( .A(_03737_ ), .B(\IF_ID_pc [18] ), .Z(_03738_ ) );
AND2_X1 _11404_ ( .A1(_03733_ ), .A2(_03738_ ), .ZN(_03739_ ) );
AND2_X1 _11405_ ( .A1(_03404_ ), .A2(\IF_ID_inst [13] ), .ZN(_03740_ ) );
INV_X1 _11406_ ( .A(_03740_ ), .ZN(_03741_ ) );
AOI21_X1 _11407_ ( .A(_03724_ ), .B1(_03741_ ), .B2(_03736_ ), .ZN(_03742_ ) );
INV_X1 _11408_ ( .A(\IF_ID_pc [13] ), .ZN(_03743_ ) );
XNOR2_X1 _11409_ ( .A(_03742_ ), .B(_03743_ ), .ZN(_03744_ ) );
AOI21_X1 _11410_ ( .A(_03714_ ), .B1(_03404_ ), .B2(\IF_ID_inst [14] ), .ZN(_03745_ ) );
NOR2_X1 _11411_ ( .A1(_03745_ ), .A2(_03716_ ), .ZN(_03746_ ) );
XNOR2_X1 _11412_ ( .A(_03746_ ), .B(_02024_ ), .ZN(_03747_ ) );
AND2_X1 _11413_ ( .A1(_03744_ ), .A2(_03747_ ), .ZN(_03748_ ) );
AND2_X1 _11414_ ( .A1(_03404_ ), .A2(\IF_ID_inst [16] ), .ZN(_03749_ ) );
OAI21_X1 _11415_ ( .A(_03725_ ), .B1(_03749_ ), .B2(_03723_ ), .ZN(_03750_ ) );
XNOR2_X1 _11416_ ( .A(_03750_ ), .B(\IF_ID_pc [16] ), .ZN(_03751_ ) );
INV_X1 _11417_ ( .A(_03751_ ), .ZN(_03752_ ) );
AND2_X1 _11418_ ( .A1(_03404_ ), .A2(\IF_ID_inst [15] ), .ZN(_03753_ ) );
OAI21_X1 _11419_ ( .A(_03725_ ), .B1(_03753_ ), .B2(_03723_ ), .ZN(_03754_ ) );
XNOR2_X1 _11420_ ( .A(_03754_ ), .B(_01993_ ), .ZN(_03755_ ) );
NOR2_X1 _11421_ ( .A1(_03752_ ), .A2(_03755_ ), .ZN(_03756_ ) );
NAND2_X1 _11422_ ( .A1(_03748_ ), .A2(_03756_ ), .ZN(_03757_ ) );
AND2_X1 _11423_ ( .A1(_03404_ ), .A2(\IF_ID_inst [20] ), .ZN(_03758_ ) );
INV_X1 _11424_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03759_ ) );
AOI21_X1 _11425_ ( .A(_03758_ ), .B1(_03759_ ), .B2(_03714_ ), .ZN(_03760_ ) );
XNOR2_X1 _11426_ ( .A(_03760_ ), .B(\IF_ID_pc [11] ), .ZN(_03761_ ) );
AOI21_X1 _11427_ ( .A(_03714_ ), .B1(_03404_ ), .B2(\IF_ID_inst [12] ), .ZN(_03762_ ) );
NOR2_X1 _11428_ ( .A1(_03762_ ), .A2(_03716_ ), .ZN(_03763_ ) );
XNOR2_X1 _11429_ ( .A(_03763_ ), .B(_01975_ ), .ZN(_03764_ ) );
AND2_X1 _11430_ ( .A1(_03761_ ), .A2(_03764_ ), .ZN(_03765_ ) );
AND2_X1 _11431_ ( .A1(_03405_ ), .A2(\IF_ID_inst [29] ), .ZN(_03766_ ) );
INV_X1 _11432_ ( .A(_03766_ ), .ZN(_03767_ ) );
INV_X1 _11433_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03768_ ) );
NAND4_X1 _11434_ ( .A1(_03402_ ), .A2(\IF_ID_inst [31] ), .A3(_03312_ ), .A4(_03768_ ), .ZN(_03769_ ) );
AND3_X1 _11435_ ( .A1(_03767_ ), .A2(_01960_ ), .A3(_03769_ ), .ZN(_03770_ ) );
AOI21_X1 _11436_ ( .A(_01960_ ), .B1(_03767_ ), .B2(_03769_ ), .ZN(_03771_ ) );
NOR2_X1 _11437_ ( .A1(_03770_ ), .A2(_03771_ ), .ZN(_03772_ ) );
AND2_X1 _11438_ ( .A1(_03404_ ), .A2(\IF_ID_inst [30] ), .ZN(_03773_ ) );
INV_X1 _11439_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03774_ ) );
AOI21_X1 _11440_ ( .A(_03773_ ), .B1(_03774_ ), .B2(_03714_ ), .ZN(_03775_ ) );
XNOR2_X1 _11441_ ( .A(_03775_ ), .B(\IF_ID_pc [10] ), .ZN(_03776_ ) );
NAND3_X1 _11442_ ( .A1(_03765_ ), .A2(_03772_ ), .A3(_03776_ ), .ZN(_03777_ ) );
AND2_X1 _11443_ ( .A1(_03403_ ), .A2(\IF_ID_inst [25] ), .ZN(_03778_ ) );
INV_X1 _11444_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03779_ ) );
AND3_X1 _11445_ ( .A1(_03311_ ), .A2(_03713_ ), .A3(_03779_ ), .ZN(_03780_ ) );
NOR2_X1 _11446_ ( .A1(_03778_ ), .A2(_03780_ ), .ZN(_03781_ ) );
INV_X1 _11447_ ( .A(\IF_ID_pc [5] ), .ZN(_03782_ ) );
XNOR2_X1 _11448_ ( .A(_03781_ ), .B(_03782_ ), .ZN(_03783_ ) );
NAND4_X1 _11449_ ( .A1(_03402_ ), .A2(\IF_ID_inst [31] ), .A3(_03311_ ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03784_ ) );
NAND3_X1 _11450_ ( .A1(_03402_ ), .A2(_03387_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_03785_ ) );
AND2_X1 _11451_ ( .A1(_03784_ ), .A2(_03785_ ), .ZN(_03786_ ) );
XOR2_X1 _11452_ ( .A(_03786_ ), .B(\IF_ID_pc [2] ), .Z(_03787_ ) );
INV_X1 _11453_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03788_ ) );
AND3_X1 _11454_ ( .A1(_03311_ ), .A2(_03713_ ), .A3(_03788_ ), .ZN(_03789_ ) );
AOI21_X1 _11455_ ( .A(_03789_ ), .B1(\IF_ID_inst [21] ), .B2(_03403_ ), .ZN(_03790_ ) );
INV_X1 _11456_ ( .A(\IF_ID_pc [1] ), .ZN(_03791_ ) );
NOR2_X2 _11457_ ( .A1(_03790_ ), .A2(_03791_ ), .ZN(_03792_ ) );
AND2_X1 _11458_ ( .A1(_03787_ ), .A2(_03792_ ), .ZN(_03793_ ) );
AND2_X1 _11459_ ( .A1(_03786_ ), .A2(\IF_ID_pc [2] ), .ZN(_03794_ ) );
NOR2_X1 _11460_ ( .A1(_03793_ ), .A2(_03794_ ), .ZN(_03795_ ) );
AND2_X1 _11461_ ( .A1(_03403_ ), .A2(\IF_ID_inst [23] ), .ZN(_03796_ ) );
INV_X1 _11462_ ( .A(_03796_ ), .ZN(_03797_ ) );
MUX2_X1 _11463_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .B(_03797_ ), .S(_03736_ ), .Z(_03798_ ) );
INV_X1 _11464_ ( .A(fanout_net_9 ), .ZN(_03799_ ) );
XNOR2_X1 _11465_ ( .A(_03798_ ), .B(_03799_ ), .ZN(_03800_ ) );
OR2_X1 _11466_ ( .A1(_03795_ ), .A2(_03800_ ), .ZN(_03801_ ) );
OR2_X2 _11467_ ( .A1(_03798_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03802_ ) );
NAND2_X1 _11468_ ( .A1(_03801_ ), .A2(_03802_ ), .ZN(_03803_ ) );
INV_X1 _11469_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03804_ ) );
NAND3_X1 _11470_ ( .A1(_03312_ ), .A2(_03713_ ), .A3(_03804_ ), .ZN(_03805_ ) );
INV_X1 _11471_ ( .A(_03403_ ), .ZN(_03806_ ) );
OAI21_X1 _11472_ ( .A(_03805_ ), .B1(_03806_ ), .B2(_03335_ ), .ZN(_03807_ ) );
OAI21_X1 _11473_ ( .A(_03803_ ), .B1(fanout_net_13 ), .B2(_03807_ ), .ZN(_03808_ ) );
NAND2_X1 _11474_ ( .A1(_03807_ ), .A2(fanout_net_13 ), .ZN(_03809_ ) );
AOI21_X2 _11475_ ( .A(_03783_ ), .B1(_03808_ ), .B2(_03809_ ), .ZN(_03810_ ) );
INV_X1 _11476_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03811_ ) );
AND3_X1 _11477_ ( .A1(_03312_ ), .A2(_03713_ ), .A3(_03811_ ), .ZN(_03812_ ) );
AOI21_X1 _11478_ ( .A(_03812_ ), .B1(\IF_ID_inst [26] ), .B2(_03404_ ), .ZN(_03813_ ) );
NOR2_X1 _11479_ ( .A1(_03813_ ), .A2(_02133_ ), .ZN(_03814_ ) );
NOR2_X1 _11480_ ( .A1(_03781_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03815_ ) );
OR3_X1 _11481_ ( .A1(_03810_ ), .A2(_03814_ ), .A3(_03815_ ), .ZN(_03816_ ) );
INV_X1 _11482_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03817_ ) );
AND3_X1 _11483_ ( .A1(_03312_ ), .A2(_03713_ ), .A3(_03817_ ), .ZN(_03818_ ) );
AOI21_X1 _11484_ ( .A(_03818_ ), .B1(\IF_ID_inst [27] ), .B2(_03405_ ), .ZN(_03819_ ) );
XNOR2_X1 _11485_ ( .A(_03819_ ), .B(\IF_ID_pc [7] ), .ZN(_03820_ ) );
NAND2_X1 _11486_ ( .A1(_03813_ ), .A2(_02133_ ), .ZN(_03821_ ) );
AND3_X2 _11487_ ( .A1(_03816_ ), .A2(_03820_ ), .A3(_03821_ ), .ZN(_03822_ ) );
INV_X1 _11488_ ( .A(_03819_ ), .ZN(_03823_ ) );
AND2_X1 _11489_ ( .A1(_03823_ ), .A2(\IF_ID_pc [7] ), .ZN(_03824_ ) );
INV_X1 _11490_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03825_ ) );
AND3_X1 _11491_ ( .A1(_03312_ ), .A2(_03713_ ), .A3(_03825_ ), .ZN(_03826_ ) );
AOI21_X1 _11492_ ( .A(_03826_ ), .B1(\IF_ID_inst [28] ), .B2(_03405_ ), .ZN(_03827_ ) );
INV_X1 _11493_ ( .A(_03827_ ), .ZN(_03828_ ) );
OAI22_X1 _11494_ ( .A1(_03822_ ), .A2(_03824_ ), .B1(\IF_ID_pc [8] ), .B2(_03828_ ), .ZN(_03829_ ) );
NOR2_X1 _11495_ ( .A1(_03827_ ), .A2(_01983_ ), .ZN(_03830_ ) );
INV_X1 _11496_ ( .A(_03830_ ), .ZN(_03831_ ) );
AOI211_X2 _11497_ ( .A(_03757_ ), .B(_03777_ ), .C1(_03829_ ), .C2(_03831_ ), .ZN(_03832_ ) );
NOR2_X1 _11498_ ( .A1(_03775_ ), .A2(_02022_ ), .ZN(_03833_ ) );
AND2_X1 _11499_ ( .A1(_03776_ ), .A2(_03771_ ), .ZN(_03834_ ) );
OAI21_X1 _11500_ ( .A(_03765_ ), .B1(_03833_ ), .B2(_03834_ ), .ZN(_03835_ ) );
NOR3_X1 _11501_ ( .A1(_03762_ ), .A2(_03724_ ), .A3(_01975_ ), .ZN(_03836_ ) );
NOR2_X1 _11502_ ( .A1(_03760_ ), .A2(_02092_ ), .ZN(_03837_ ) );
AOI21_X1 _11503_ ( .A(_03836_ ), .B1(_03764_ ), .B2(_03837_ ), .ZN(_03838_ ) );
AOI21_X1 _11504_ ( .A(_03757_ ), .B1(_03835_ ), .B2(_03838_ ), .ZN(_03839_ ) );
AND3_X1 _11505_ ( .A1(_03747_ ), .A2(\IF_ID_pc [13] ), .A3(_03742_ ), .ZN(_03840_ ) );
AND2_X1 _11506_ ( .A1(_03746_ ), .A2(\IF_ID_pc [14] ), .ZN(_03841_ ) );
OR2_X1 _11507_ ( .A1(_03840_ ), .A2(_03841_ ), .ZN(_03842_ ) );
AND2_X1 _11508_ ( .A1(_03842_ ), .A2(_03756_ ), .ZN(_03843_ ) );
NOR2_X1 _11509_ ( .A1(_03754_ ), .A2(_01993_ ), .ZN(_03844_ ) );
NAND2_X1 _11510_ ( .A1(_03751_ ), .A2(_03844_ ), .ZN(_03845_ ) );
OAI21_X1 _11511_ ( .A(_03845_ ), .B1(_02181_ ), .B2(_03750_ ), .ZN(_03846_ ) );
OR3_X1 _11512_ ( .A1(_03839_ ), .A2(_03843_ ), .A3(_03846_ ), .ZN(_03847_ ) );
OAI211_X1 _11513_ ( .A(_03729_ ), .B(_03739_ ), .C1(_03832_ ), .C2(_03847_ ), .ZN(_03848_ ) );
AND2_X1 _11514_ ( .A1(_03732_ ), .A2(\IF_ID_pc [17] ), .ZN(_03849_ ) );
AND2_X1 _11515_ ( .A1(_03738_ ), .A2(_03849_ ), .ZN(_03850_ ) );
AOI21_X1 _11516_ ( .A(_03850_ ), .B1(\IF_ID_pc [18] ), .B2(_03737_ ), .ZN(_03851_ ) );
INV_X1 _11517_ ( .A(_03851_ ), .ZN(_03852_ ) );
AND2_X1 _11518_ ( .A1(_03852_ ), .A2(_03729_ ), .ZN(_03853_ ) );
AND2_X1 _11519_ ( .A1(_03717_ ), .A2(\IF_ID_pc [20] ), .ZN(_03854_ ) );
NOR2_X1 _11520_ ( .A1(_03727_ ), .A2(_02064_ ), .ZN(_03855_ ) );
AND2_X1 _11521_ ( .A1(_03721_ ), .A2(_03855_ ), .ZN(_03856_ ) );
NOR3_X1 _11522_ ( .A1(_03853_ ), .A2(_03854_ ), .A3(_03856_ ), .ZN(_03857_ ) );
NAND2_X1 _11523_ ( .A1(_03848_ ), .A2(_03857_ ), .ZN(_03858_ ) );
XNOR2_X1 _11524_ ( .A(_03718_ ), .B(_02032_ ), .ZN(_03859_ ) );
XNOR2_X1 _11525_ ( .A(_03718_ ), .B(_02166_ ), .ZN(_03860_ ) );
XNOR2_X1 _11526_ ( .A(_03717_ ), .B(_01951_ ), .ZN(_03861_ ) );
AND2_X1 _11527_ ( .A1(_03860_ ), .A2(_03861_ ), .ZN(_03862_ ) );
AND4_X1 _11528_ ( .A1(_03720_ ), .A2(_03858_ ), .A3(_03859_ ), .A4(_03862_ ), .ZN(_03863_ ) );
OAI21_X1 _11529_ ( .A(_03718_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_03864_ ) );
INV_X1 _11530_ ( .A(_03864_ ), .ZN(_03865_ ) );
NAND3_X1 _11531_ ( .A1(_03720_ ), .A2(_03859_ ), .A3(_03865_ ), .ZN(_03866_ ) );
NAND2_X1 _11532_ ( .A1(_03718_ ), .A2(\IF_ID_pc [24] ), .ZN(_03867_ ) );
NAND2_X1 _11533_ ( .A1(_03718_ ), .A2(\IF_ID_pc [23] ), .ZN(_03868_ ) );
AND3_X1 _11534_ ( .A1(_03866_ ), .A2(_03867_ ), .A3(_03868_ ), .ZN(_03869_ ) );
INV_X1 _11535_ ( .A(_03869_ ), .ZN(_03870_ ) );
OAI21_X2 _11536_ ( .A(_03719_ ), .B1(_03863_ ), .B2(_03870_ ), .ZN(_03871_ ) );
XNOR2_X1 _11537_ ( .A(_03718_ ), .B(_02111_ ), .ZN(_03872_ ) );
INV_X1 _11538_ ( .A(_03872_ ), .ZN(_03873_ ) );
NOR2_X1 _11539_ ( .A1(_03871_ ), .A2(_03873_ ), .ZN(_03874_ ) );
BUF_X4 _11540_ ( .A(_03718_ ), .Z(_03875_ ) );
XNOR2_X1 _11541_ ( .A(_03875_ ), .B(_02056_ ), .ZN(_03876_ ) );
XOR2_X1 _11542_ ( .A(_03718_ ), .B(\IF_ID_pc [27] ), .Z(_03877_ ) );
AND3_X1 _11543_ ( .A1(_03874_ ), .A2(_03876_ ), .A3(_03877_ ), .ZN(_03878_ ) );
OAI21_X1 _11544_ ( .A(_03875_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_03879_ ) );
INV_X1 _11545_ ( .A(_03879_ ), .ZN(_03880_ ) );
NAND3_X1 _11546_ ( .A1(_03877_ ), .A2(_03876_ ), .A3(_03880_ ), .ZN(_03881_ ) );
NAND2_X1 _11547_ ( .A1(_03875_ ), .A2(\IF_ID_pc [28] ), .ZN(_03882_ ) );
NAND2_X1 _11548_ ( .A1(_03875_ ), .A2(\IF_ID_pc [27] ), .ZN(_03883_ ) );
NAND3_X1 _11549_ ( .A1(_03881_ ), .A2(_03882_ ), .A3(_03883_ ), .ZN(_03884_ ) );
NOR2_X2 _11550_ ( .A1(_03878_ ), .A2(_03884_ ), .ZN(_03885_ ) );
XNOR2_X1 _11551_ ( .A(_03875_ ), .B(\IF_ID_pc [29] ), .ZN(_03886_ ) );
NOR2_X1 _11552_ ( .A1(_03885_ ), .A2(_03886_ ), .ZN(_03887_ ) );
NOR3_X1 _11553_ ( .A1(_03715_ ), .A2(_03724_ ), .A3(_02087_ ), .ZN(_03888_ ) );
NOR2_X1 _11554_ ( .A1(_03887_ ), .A2(_03888_ ), .ZN(_03889_ ) );
XNOR2_X1 _11555_ ( .A(_03875_ ), .B(\IF_ID_pc [30] ), .ZN(_03890_ ) );
OR2_X1 _11556_ ( .A1(_03889_ ), .A2(_03890_ ), .ZN(_03891_ ) );
AOI21_X1 _11557_ ( .A(_03538_ ), .B1(_03889_ ), .B2(_03890_ ), .ZN(_03892_ ) );
AOI221_X4 _11558_ ( .A(\myifu.to_reset ), .B1(\myexu.pc_jump [30] ), .B2(_03538_ ), .C1(_03891_ ), .C2(_03892_ ), .ZN(_03893_ ) );
BUF_X4 _11559_ ( .A(_03709_ ), .Z(_03894_ ) );
BUF_X4 _11560_ ( .A(_03894_ ), .Z(_03895_ ) );
NOR2_X1 _11561_ ( .A1(_03895_ ), .A2(\mtvec [30] ), .ZN(_03896_ ) );
NOR3_X1 _11562_ ( .A1(_03893_ ), .A2(fanout_net_4 ), .A3(_03896_ ), .ZN(_00282_ ) );
XOR2_X1 _11563_ ( .A(_03858_ ), .B(_03861_ ), .Z(_03897_ ) );
INV_X1 _11564_ ( .A(_03538_ ), .ZN(_03898_ ) );
BUF_X4 _11565_ ( .A(_03898_ ), .Z(_03899_ ) );
BUF_X4 _11566_ ( .A(_03899_ ), .Z(_03900_ ) );
MUX2_X1 _11567_ ( .A(\myexu.pc_jump [21] ), .B(_03897_ ), .S(_03900_ ), .Z(_03901_ ) );
MUX2_X1 _11568_ ( .A(\mtvec [21] ), .B(_03901_ ), .S(_03894_ ), .Z(_03902_ ) );
CLKBUF_X2 _11569_ ( .A(_01664_ ), .Z(_03903_ ) );
AND2_X1 _11570_ ( .A1(_03902_ ), .A2(_03903_ ), .ZN(_00283_ ) );
OAI21_X1 _11571_ ( .A(_03739_ ), .B1(_03832_ ), .B2(_03847_ ), .ZN(_03904_ ) );
NAND2_X1 _11572_ ( .A1(_03904_ ), .A2(_03851_ ), .ZN(_03905_ ) );
AOI21_X1 _11573_ ( .A(_03855_ ), .B1(_03905_ ), .B2(_03728_ ), .ZN(_03906_ ) );
XNOR2_X1 _11574_ ( .A(_03906_ ), .B(_03721_ ), .ZN(_03907_ ) );
MUX2_X1 _11575_ ( .A(\myexu.pc_jump [20] ), .B(_03907_ ), .S(_03900_ ), .Z(_03908_ ) );
MUX2_X1 _11576_ ( .A(\mtvec [20] ), .B(_03908_ ), .S(_03894_ ), .Z(_03909_ ) );
AND2_X1 _11577_ ( .A1(_03909_ ), .A2(_03903_ ), .ZN(_00284_ ) );
XNOR2_X1 _11578_ ( .A(_03905_ ), .B(_03728_ ), .ZN(_03910_ ) );
BUF_X4 _11579_ ( .A(_03900_ ), .Z(_03911_ ) );
NAND2_X1 _11580_ ( .A1(_03910_ ), .A2(_03911_ ), .ZN(_03912_ ) );
BUF_X4 _11581_ ( .A(_03900_ ), .Z(_03913_ ) );
OAI211_X1 _11582_ ( .A(_03912_ ), .B(_03895_ ), .C1(\myexu.pc_jump [19] ), .C2(_03913_ ), .ZN(_03914_ ) );
NAND2_X1 _11583_ ( .A1(\mtvec [19] ), .A2(\myifu.to_reset ), .ZN(_03915_ ) );
AOI21_X1 _11584_ ( .A(fanout_net_4 ), .B1(_03914_ ), .B2(_03915_ ), .ZN(_00285_ ) );
OAI21_X1 _11585_ ( .A(_03733_ ), .B1(_03832_ ), .B2(_03847_ ), .ZN(_03916_ ) );
INV_X1 _11586_ ( .A(_03849_ ), .ZN(_03917_ ) );
AND2_X1 _11587_ ( .A1(_03916_ ), .A2(_03917_ ), .ZN(_03918_ ) );
XNOR2_X1 _11588_ ( .A(_03918_ ), .B(_03738_ ), .ZN(_03919_ ) );
MUX2_X1 _11589_ ( .A(\myexu.pc_jump [18] ), .B(_03919_ ), .S(_03899_ ), .Z(_03920_ ) );
MUX2_X1 _11590_ ( .A(\mtvec [18] ), .B(_03920_ ), .S(_03894_ ), .Z(_03921_ ) );
AND2_X1 _11591_ ( .A1(_03921_ ), .A2(_03903_ ), .ZN(_00286_ ) );
NOR2_X1 _11592_ ( .A1(_03832_ ), .A2(_03847_ ), .ZN(_03922_ ) );
XOR2_X1 _11593_ ( .A(_03922_ ), .B(_03733_ ), .Z(_03923_ ) );
NAND2_X1 _11594_ ( .A1(_03923_ ), .A2(_03911_ ), .ZN(_03924_ ) );
OAI211_X1 _11595_ ( .A(_03924_ ), .B(_03895_ ), .C1(\myexu.pc_jump [17] ), .C2(_03913_ ), .ZN(_03925_ ) );
NAND2_X1 _11596_ ( .A1(\mtvec [17] ), .A2(\myifu.to_reset ), .ZN(_03926_ ) );
AOI21_X1 _11597_ ( .A(fanout_net_4 ), .B1(_03925_ ), .B2(_03926_ ), .ZN(_00287_ ) );
AOI21_X1 _11598_ ( .A(_03777_ ), .B1(_03829_ ), .B2(_03831_ ), .ZN(_03927_ ) );
INV_X1 _11599_ ( .A(_03927_ ), .ZN(_03928_ ) );
AND2_X1 _11600_ ( .A1(_03835_ ), .A2(_03838_ ), .ZN(_03929_ ) );
NAND2_X1 _11601_ ( .A1(_03928_ ), .A2(_03929_ ), .ZN(_03930_ ) );
AOI21_X1 _11602_ ( .A(_03842_ ), .B1(_03930_ ), .B2(_03748_ ), .ZN(_03931_ ) );
NOR2_X1 _11603_ ( .A1(_03931_ ), .A2(_03755_ ), .ZN(_03932_ ) );
NOR2_X1 _11604_ ( .A1(_03932_ ), .A2(_03844_ ), .ZN(_03933_ ) );
XNOR2_X1 _11605_ ( .A(_03933_ ), .B(_03751_ ), .ZN(_03934_ ) );
MUX2_X1 _11606_ ( .A(\myexu.pc_jump [16] ), .B(_03934_ ), .S(_03899_ ), .Z(_03935_ ) );
MUX2_X1 _11607_ ( .A(\mtvec [16] ), .B(_03935_ ), .S(_03894_ ), .Z(_03936_ ) );
AND2_X1 _11608_ ( .A1(_03936_ ), .A2(_03903_ ), .ZN(_00288_ ) );
XOR2_X1 _11609_ ( .A(_03931_ ), .B(_03755_ ), .Z(_03937_ ) );
MUX2_X1 _11610_ ( .A(\myexu.pc_jump [15] ), .B(_03937_ ), .S(_03899_ ), .Z(_03938_ ) );
MUX2_X1 _11611_ ( .A(\mtvec [15] ), .B(_03938_ ), .S(_03894_ ), .Z(_03939_ ) );
AND2_X1 _11612_ ( .A1(_03939_ ), .A2(_03903_ ), .ZN(_00289_ ) );
AND2_X1 _11613_ ( .A1(_03930_ ), .A2(_03744_ ), .ZN(_03940_ ) );
AOI21_X1 _11614_ ( .A(_03940_ ), .B1(\IF_ID_pc [13] ), .B2(_03742_ ), .ZN(_03941_ ) );
XNOR2_X1 _11615_ ( .A(_03941_ ), .B(_03747_ ), .ZN(_03942_ ) );
MUX2_X1 _11616_ ( .A(\myexu.pc_jump [14] ), .B(_03942_ ), .S(_03899_ ), .Z(_03943_ ) );
MUX2_X1 _11617_ ( .A(\mtvec [14] ), .B(_03943_ ), .S(_03894_ ), .Z(_03944_ ) );
AND2_X1 _11618_ ( .A1(_03944_ ), .A2(_03903_ ), .ZN(_00290_ ) );
NOR2_X1 _11619_ ( .A1(_03930_ ), .A2(_03744_ ), .ZN(_03945_ ) );
OAI21_X1 _11620_ ( .A(_03911_ ), .B1(_03940_ ), .B2(_03945_ ), .ZN(_03946_ ) );
OAI211_X1 _11621_ ( .A(_03946_ ), .B(_03895_ ), .C1(\myexu.pc_jump [13] ), .C2(_03913_ ), .ZN(_03947_ ) );
NAND2_X1 _11622_ ( .A1(\mtvec [13] ), .A2(\myifu.to_reset ), .ZN(_03948_ ) );
AOI21_X1 _11623_ ( .A(fanout_net_4 ), .B1(_03947_ ), .B2(_03948_ ), .ZN(_00291_ ) );
NOR2_X1 _11624_ ( .A1(_03710_ ), .A2(\mtvec [12] ), .ZN(_03949_ ) );
INV_X1 _11625_ ( .A(_03772_ ), .ZN(_03950_ ) );
AOI21_X1 _11626_ ( .A(_03950_ ), .B1(_03829_ ), .B2(_03831_ ), .ZN(_03951_ ) );
OR3_X1 _11627_ ( .A1(_03951_ ), .A2(_03833_ ), .A3(_03771_ ), .ZN(_03952_ ) );
AND2_X1 _11628_ ( .A1(_03775_ ), .A2(_02022_ ), .ZN(_03953_ ) );
INV_X1 _11629_ ( .A(_03953_ ), .ZN(_03954_ ) );
AND3_X1 _11630_ ( .A1(_03952_ ), .A2(_03761_ ), .A3(_03954_ ), .ZN(_03955_ ) );
OR3_X1 _11631_ ( .A1(_03955_ ), .A2(_03837_ ), .A3(_03764_ ), .ZN(_03956_ ) );
OAI21_X1 _11632_ ( .A(_03764_ ), .B1(_03955_ ), .B2(_03837_ ), .ZN(_03957_ ) );
NAND3_X1 _11633_ ( .A1(_03956_ ), .A2(_03913_ ), .A3(_03957_ ), .ZN(_03958_ ) );
BUF_X4 _11634_ ( .A(_03538_ ), .Z(_03959_ ) );
AOI21_X1 _11635_ ( .A(\myifu.to_reset ), .B1(_03959_ ), .B2(\myexu.pc_jump [12] ), .ZN(_03960_ ) );
AOI211_X1 _11636_ ( .A(fanout_net_4 ), .B(_03949_ ), .C1(_03958_ ), .C2(_03960_ ), .ZN(_00292_ ) );
AND2_X1 _11637_ ( .A1(_03885_ ), .A2(_03886_ ), .ZN(_03961_ ) );
OAI21_X1 _11638_ ( .A(_03911_ ), .B1(_03961_ ), .B2(_03887_ ), .ZN(_03962_ ) );
OAI211_X1 _11639_ ( .A(_03962_ ), .B(_03895_ ), .C1(\myexu.pc_jump [29] ), .C2(_03913_ ), .ZN(_03963_ ) );
NAND2_X1 _11640_ ( .A1(\mtvec [29] ), .A2(\myifu.to_reset ), .ZN(_03964_ ) );
AOI21_X1 _11641_ ( .A(fanout_net_4 ), .B1(_03963_ ), .B2(_03964_ ), .ZN(_00293_ ) );
AOI21_X1 _11642_ ( .A(_03761_ ), .B1(_03952_ ), .B2(_03954_ ), .ZN(_03965_ ) );
OAI21_X1 _11643_ ( .A(_03911_ ), .B1(_03955_ ), .B2(_03965_ ), .ZN(_03966_ ) );
OAI211_X1 _11644_ ( .A(_03966_ ), .B(_03710_ ), .C1(\myexu.pc_jump [11] ), .C2(_03913_ ), .ZN(_03967_ ) );
NAND2_X1 _11645_ ( .A1(\mtvec [11] ), .A2(\myifu.to_reset ), .ZN(_03968_ ) );
AOI21_X1 _11646_ ( .A(fanout_net_4 ), .B1(_03967_ ), .B2(_03968_ ), .ZN(_00294_ ) );
NOR2_X1 _11647_ ( .A1(_03951_ ), .A2(_03771_ ), .ZN(_03969_ ) );
INV_X1 _11648_ ( .A(_03969_ ), .ZN(_03970_ ) );
OAI21_X1 _11649_ ( .A(_03900_ ), .B1(_03970_ ), .B2(_03776_ ), .ZN(_03971_ ) );
AOI21_X1 _11650_ ( .A(_03971_ ), .B1(_03970_ ), .B2(_03776_ ), .ZN(_03972_ ) );
AOI211_X1 _11651_ ( .A(\myifu.to_reset ), .B(_03972_ ), .C1(\myexu.pc_jump [10] ), .C2(_03959_ ), .ZN(_03973_ ) );
NOR2_X1 _11652_ ( .A1(_03895_ ), .A2(\mtvec [10] ), .ZN(_03974_ ) );
NOR3_X1 _11653_ ( .A1(_03973_ ), .A2(fanout_net_4 ), .A3(_03974_ ), .ZN(_00295_ ) );
AND3_X1 _11654_ ( .A1(_03829_ ), .A2(_03831_ ), .A3(_03950_ ), .ZN(_03975_ ) );
OAI21_X1 _11655_ ( .A(_03911_ ), .B1(_03975_ ), .B2(_03951_ ), .ZN(_03976_ ) );
OAI211_X1 _11656_ ( .A(_03976_ ), .B(_03710_ ), .C1(\myexu.pc_jump [9] ), .C2(_03913_ ), .ZN(_03977_ ) );
NAND2_X1 _11657_ ( .A1(\mtvec [9] ), .A2(\myifu.to_reset ), .ZN(_03978_ ) );
AOI21_X1 _11658_ ( .A(fanout_net_4 ), .B1(_03977_ ), .B2(_03978_ ), .ZN(_00296_ ) );
NOR2_X1 _11659_ ( .A1(_03822_ ), .A2(_03824_ ), .ZN(_03979_ ) );
INV_X1 _11660_ ( .A(_03979_ ), .ZN(_03980_ ) );
XNOR2_X1 _11661_ ( .A(_03827_ ), .B(\IF_ID_pc [8] ), .ZN(_03981_ ) );
OAI21_X1 _11662_ ( .A(_03900_ ), .B1(_03980_ ), .B2(_03981_ ), .ZN(_03982_ ) );
AOI21_X1 _11663_ ( .A(_03982_ ), .B1(_03980_ ), .B2(_03981_ ), .ZN(_03983_ ) );
AOI211_X1 _11664_ ( .A(\myifu.to_reset ), .B(_03983_ ), .C1(\myexu.pc_jump [8] ), .C2(_03959_ ), .ZN(_03984_ ) );
NOR2_X1 _11665_ ( .A1(_03895_ ), .A2(\mtvec [8] ), .ZN(_03985_ ) );
NOR3_X1 _11666_ ( .A1(_03984_ ), .A2(fanout_net_4 ), .A3(_03985_ ), .ZN(_00297_ ) );
NAND2_X1 _11667_ ( .A1(_03816_ ), .A2(_03821_ ), .ZN(_03986_ ) );
XNOR2_X1 _11668_ ( .A(_03986_ ), .B(_03820_ ), .ZN(_03987_ ) );
MUX2_X1 _11669_ ( .A(\myexu.pc_jump [7] ), .B(_03987_ ), .S(_03899_ ), .Z(_03988_ ) );
MUX2_X1 _11670_ ( .A(\mtvec [7] ), .B(_03988_ ), .S(_03894_ ), .Z(_03989_ ) );
AND2_X1 _11671_ ( .A1(_03989_ ), .A2(_03903_ ), .ZN(_00298_ ) );
XNOR2_X1 _11672_ ( .A(_03813_ ), .B(_02133_ ), .ZN(_03990_ ) );
OR3_X1 _11673_ ( .A1(_03810_ ), .A2(_03815_ ), .A3(_03990_ ), .ZN(_03991_ ) );
OAI21_X1 _11674_ ( .A(_03990_ ), .B1(_03810_ ), .B2(_03815_ ), .ZN(_03992_ ) );
AOI21_X1 _11675_ ( .A(_03959_ ), .B1(_03991_ ), .B2(_03992_ ), .ZN(_03993_ ) );
AOI211_X1 _11676_ ( .A(\myifu.to_reset ), .B(_03993_ ), .C1(\myexu.pc_jump [6] ), .C2(_03959_ ), .ZN(_03994_ ) );
NOR2_X1 _11677_ ( .A1(_03895_ ), .A2(\mtvec [6] ), .ZN(_03995_ ) );
NOR3_X1 _11678_ ( .A1(_03994_ ), .A2(fanout_net_4 ), .A3(_03995_ ), .ZN(_00299_ ) );
AND3_X1 _11679_ ( .A1(_03808_ ), .A2(_03809_ ), .A3(_03783_ ), .ZN(_03996_ ) );
OAI21_X1 _11680_ ( .A(_03911_ ), .B1(_03996_ ), .B2(_03810_ ), .ZN(_03997_ ) );
OAI211_X1 _11681_ ( .A(_03997_ ), .B(_03710_ ), .C1(\myexu.pc_jump [5] ), .C2(_03913_ ), .ZN(_03998_ ) );
NAND2_X1 _11682_ ( .A1(\mtvec [5] ), .A2(\myifu.to_reset ), .ZN(_03999_ ) );
AOI21_X1 _11683_ ( .A(fanout_net_4 ), .B1(_03998_ ), .B2(_03999_ ), .ZN(_00300_ ) );
AND2_X1 _11684_ ( .A1(\mtvec [4] ), .A2(\myifu.to_reset ), .ZN(_04000_ ) );
XNOR2_X1 _11685_ ( .A(_03807_ ), .B(fanout_net_13 ), .ZN(_04001_ ) );
XNOR2_X1 _11686_ ( .A(_03803_ ), .B(_04001_ ), .ZN(_04002_ ) );
MUX2_X1 _11687_ ( .A(\myexu.pc_jump [4] ), .B(_04002_ ), .S(_03900_ ), .Z(_04003_ ) );
AOI21_X1 _11688_ ( .A(_04000_ ), .B1(_04003_ ), .B2(_03895_ ), .ZN(_04004_ ) );
NOR2_X1 _11689_ ( .A1(_04004_ ), .A2(fanout_net_4 ), .ZN(_00301_ ) );
XOR2_X1 _11690_ ( .A(_03795_ ), .B(_03800_ ), .Z(_04005_ ) );
MUX2_X1 _11691_ ( .A(\myexu.pc_jump [3] ), .B(_04005_ ), .S(_03898_ ), .Z(_04006_ ) );
AND2_X1 _11692_ ( .A1(_04006_ ), .A2(_03709_ ), .ZN(_04007_ ) );
AOI21_X1 _11693_ ( .A(_04007_ ), .B1(\mtvec [3] ), .B2(\myifu.to_reset ), .ZN(_04008_ ) );
NOR2_X1 _11694_ ( .A1(_04008_ ), .A2(fanout_net_4 ), .ZN(_00302_ ) );
AND2_X1 _11695_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
INV_X1 _11696_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_04009_ ) );
AOI211_X1 _11697_ ( .A(_04000_ ), .B(_04009_ ), .C1(_04003_ ), .C2(_03710_ ), .ZN(_04010_ ) );
INV_X1 _11698_ ( .A(fanout_net_13 ), .ZN(_04011_ ) );
BUF_X2 _11699_ ( .A(_04011_ ), .Z(_04012_ ) );
BUF_X2 _11700_ ( .A(_04012_ ), .Z(_04013_ ) );
BUF_X2 _11701_ ( .A(_04013_ ), .Z(_04014_ ) );
AOI211_X1 _11702_ ( .A(fanout_net_4 ), .B(_04010_ ), .C1(_04014_ ), .C2(_04009_ ), .ZN(_00303_ ) );
NOR2_X1 _11703_ ( .A1(_03787_ ), .A2(_03792_ ), .ZN(_04015_ ) );
OAI21_X1 _11704_ ( .A(_03911_ ), .B1(_03793_ ), .B2(_04015_ ), .ZN(_04016_ ) );
OAI211_X1 _11705_ ( .A(_04016_ ), .B(_03710_ ), .C1(\myexu.pc_jump [2] ), .C2(_03913_ ), .ZN(_04017_ ) );
NAND2_X1 _11706_ ( .A1(\mtvec [2] ), .A2(\myifu.to_reset ), .ZN(_04018_ ) );
AOI21_X1 _11707_ ( .A(fanout_net_4 ), .B1(_04017_ ), .B2(_04018_ ), .ZN(_00304_ ) );
AOI211_X1 _11708_ ( .A(_04009_ ), .B(_04007_ ), .C1(\mtvec [3] ), .C2(\myifu.to_reset ), .ZN(_04019_ ) );
BUF_X4 _11709_ ( .A(_03799_ ), .Z(_04020_ ) );
BUF_X2 _11710_ ( .A(_04020_ ), .Z(_04021_ ) );
AOI211_X1 _11711_ ( .A(fanout_net_4 ), .B(_04019_ ), .C1(_04021_ ), .C2(_04009_ ), .ZN(_00305_ ) );
OAI21_X1 _11712_ ( .A(_03877_ ), .B1(_03874_ ), .B2(_03880_ ), .ZN(_04022_ ) );
AND3_X1 _11713_ ( .A1(_04022_ ), .A2(_03876_ ), .A3(_03883_ ), .ZN(_04023_ ) );
AOI21_X1 _11714_ ( .A(_03876_ ), .B1(_04022_ ), .B2(_03883_ ), .ZN(_04024_ ) );
OR3_X1 _11715_ ( .A1(_04023_ ), .A2(_04024_ ), .A3(_03538_ ), .ZN(_04025_ ) );
OAI211_X1 _11716_ ( .A(_04025_ ), .B(_03710_ ), .C1(\myexu.pc_jump [28] ), .C2(_03911_ ), .ZN(_04026_ ) );
NAND2_X1 _11717_ ( .A1(\mtvec [28] ), .A2(\myifu.to_reset ), .ZN(_04027_ ) );
AOI21_X1 _11718_ ( .A(fanout_net_4 ), .B1(_04026_ ), .B2(_04027_ ), .ZN(_00306_ ) );
INV_X1 _11719_ ( .A(_03514_ ), .ZN(_04028_ ) );
INV_X1 _11720_ ( .A(_03535_ ), .ZN(_04029_ ) );
OAI211_X1 _11721_ ( .A(check_quest ), .B(\myexu.pc_jump [1] ), .C1(_04028_ ), .C2(_04029_ ), .ZN(_04030_ ) );
XNOR2_X1 _11722_ ( .A(_03790_ ), .B(_03791_ ), .ZN(_04031_ ) );
OAI211_X1 _11723_ ( .A(_03710_ ), .B(_04030_ ), .C1(_03959_ ), .C2(_04031_ ), .ZN(_04032_ ) );
OR2_X1 _11724_ ( .A1(_03894_ ), .A2(\mtvec [1] ), .ZN(_04033_ ) );
AND3_X1 _11725_ ( .A1(_04032_ ), .A2(_01758_ ), .A3(_04033_ ), .ZN(_00307_ ) );
OR3_X1 _11726_ ( .A1(_03874_ ), .A2(_03877_ ), .A3(_03880_ ), .ZN(_04034_ ) );
AND3_X1 _11727_ ( .A1(_04034_ ), .A2(_03900_ ), .A3(_04022_ ), .ZN(_04035_ ) );
AOI211_X1 _11728_ ( .A(\myifu.to_reset ), .B(_04035_ ), .C1(\myexu.pc_jump [27] ), .C2(_03959_ ), .ZN(_04036_ ) );
NOR2_X1 _11729_ ( .A1(_03895_ ), .A2(\mtvec [27] ), .ZN(_04037_ ) );
NOR3_X1 _11730_ ( .A1(_04036_ ), .A2(fanout_net_4 ), .A3(_04037_ ), .ZN(_00308_ ) );
NAND2_X1 _11731_ ( .A1(_03875_ ), .A2(\IF_ID_pc [25] ), .ZN(_04038_ ) );
NAND2_X1 _11732_ ( .A1(_03871_ ), .A2(_04038_ ), .ZN(_04039_ ) );
XNOR2_X1 _11733_ ( .A(_04039_ ), .B(_03873_ ), .ZN(_04040_ ) );
MUX2_X1 _11734_ ( .A(\myexu.pc_jump [26] ), .B(_04040_ ), .S(_03899_ ), .Z(_04041_ ) );
MUX2_X1 _11735_ ( .A(\mtvec [26] ), .B(_04041_ ), .S(_03894_ ), .Z(_04042_ ) );
AND2_X1 _11736_ ( .A1(_04042_ ), .A2(_03903_ ), .ZN(_00309_ ) );
INV_X1 _11737_ ( .A(_03871_ ), .ZN(_04043_ ) );
NOR3_X1 _11738_ ( .A1(_03863_ ), .A2(_03870_ ), .A3(_03719_ ), .ZN(_04044_ ) );
OAI21_X1 _11739_ ( .A(_03900_ ), .B1(_04043_ ), .B2(_04044_ ), .ZN(_04045_ ) );
OAI211_X1 _11740_ ( .A(_04045_ ), .B(_03710_ ), .C1(\myexu.pc_jump [25] ), .C2(_03911_ ), .ZN(_04046_ ) );
NAND2_X1 _11741_ ( .A1(\mtvec [25] ), .A2(\myifu.to_reset ), .ZN(_04047_ ) );
AOI21_X1 _11742_ ( .A(fanout_net_4 ), .B1(_04046_ ), .B2(_04047_ ), .ZN(_00310_ ) );
NAND2_X1 _11743_ ( .A1(_03858_ ), .A2(_03862_ ), .ZN(_04048_ ) );
NAND2_X1 _11744_ ( .A1(_04048_ ), .A2(_03864_ ), .ZN(_04049_ ) );
NAND2_X1 _11745_ ( .A1(_04049_ ), .A2(_03859_ ), .ZN(_04050_ ) );
AND2_X1 _11746_ ( .A1(_04050_ ), .A2(_03868_ ), .ZN(_04051_ ) );
XNOR2_X1 _11747_ ( .A(_04051_ ), .B(_03720_ ), .ZN(_04052_ ) );
MUX2_X1 _11748_ ( .A(\myexu.pc_jump [24] ), .B(_04052_ ), .S(_03899_ ), .Z(_04053_ ) );
MUX2_X1 _11749_ ( .A(\mtvec [24] ), .B(_04053_ ), .S(_03709_ ), .Z(_04054_ ) );
AND2_X1 _11750_ ( .A1(_04054_ ), .A2(_01813_ ), .ZN(_00311_ ) );
XOR2_X1 _11751_ ( .A(_04049_ ), .B(_03859_ ), .Z(_04055_ ) );
MUX2_X1 _11752_ ( .A(\myexu.pc_jump [23] ), .B(_04055_ ), .S(_03899_ ), .Z(_04056_ ) );
MUX2_X1 _11753_ ( .A(\mtvec [23] ), .B(_04056_ ), .S(_03709_ ), .Z(_04057_ ) );
AND2_X1 _11754_ ( .A1(_04057_ ), .A2(_01813_ ), .ZN(_00312_ ) );
AND2_X1 _11755_ ( .A1(_03858_ ), .A2(_03861_ ), .ZN(_04058_ ) );
AND2_X1 _11756_ ( .A1(_03875_ ), .A2(\IF_ID_pc [21] ), .ZN(_04059_ ) );
NOR2_X1 _11757_ ( .A1(_04058_ ), .A2(_04059_ ), .ZN(_04060_ ) );
XNOR2_X1 _11758_ ( .A(_04060_ ), .B(_03860_ ), .ZN(_04061_ ) );
MUX2_X1 _11759_ ( .A(\myexu.pc_jump [22] ), .B(_04061_ ), .S(_03899_ ), .Z(_04062_ ) );
MUX2_X1 _11760_ ( .A(\mtvec [22] ), .B(_04062_ ), .S(_03709_ ), .Z(_04063_ ) );
AND2_X1 _11761_ ( .A1(_04063_ ), .A2(_01813_ ), .ZN(_00313_ ) );
OAI21_X1 _11762_ ( .A(_03709_ ), .B1(_03900_ ), .B2(\myexu.pc_jump [31] ), .ZN(_04064_ ) );
OR3_X1 _11763_ ( .A1(_03885_ ), .A2(_03886_ ), .A3(_03890_ ), .ZN(_04065_ ) );
OAI21_X1 _11764_ ( .A(_03875_ ), .B1(\IF_ID_pc [30] ), .B2(\IF_ID_pc [29] ), .ZN(_04066_ ) );
AND2_X1 _11765_ ( .A1(_04065_ ), .A2(_04066_ ), .ZN(_04067_ ) );
XNOR2_X1 _11766_ ( .A(_03875_ ), .B(_02042_ ), .ZN(_04068_ ) );
OR2_X1 _11767_ ( .A1(_04067_ ), .A2(_04068_ ), .ZN(_04069_ ) );
AOI21_X2 _11768_ ( .A(_03959_ ), .B1(_04067_ ), .B2(_04068_ ), .ZN(_04070_ ) );
AOI21_X1 _11769_ ( .A(_04064_ ), .B1(_04069_ ), .B2(_04070_ ), .ZN(_04071_ ) );
AND2_X1 _11770_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_04072_ ) );
OR3_X1 _11771_ ( .A1(_04071_ ), .A2(fanout_net_5 ), .A3(_04072_ ), .ZN(_00314_ ) );
OR2_X1 _11772_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [19] ), .ZN(_04073_ ) );
NOR3_X1 _11773_ ( .A1(_04073_ ), .A2(\io_master_araddr [22] ), .A3(\io_master_araddr [16] ), .ZN(_04074_ ) );
AND4_X1 _11774_ ( .A1(_02193_ ), .A2(_02211_ ), .A3(_02158_ ), .A4(_02174_ ), .ZN(_04075_ ) );
NAND2_X1 _11775_ ( .A1(_04074_ ), .A2(_04075_ ), .ZN(_04076_ ) );
AND4_X1 _11776_ ( .A1(_02162_ ), .A2(_02178_ ), .A3(_02197_ ), .A4(_02215_ ), .ZN(_04077_ ) );
AND4_X1 _11777_ ( .A1(_02201_ ), .A2(_02219_ ), .A3(_02206_ ), .A4(\io_master_araddr [25] ), .ZN(_04078_ ) );
NAND2_X4 _11778_ ( .A1(_04077_ ), .A2(_04078_ ), .ZN(_04079_ ) );
NOR2_X4 _11779_ ( .A1(_04076_ ), .A2(_04079_ ), .ZN(_04080_ ) );
INV_X1 _11780_ ( .A(_04080_ ), .ZN(_04081_ ) );
NOR2_X1 _11781_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_04082_ ) );
NOR2_X1 _11782_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_04083_ ) );
INV_X1 _11783_ ( .A(\io_master_rid [1] ), .ZN(_04084_ ) );
NAND4_X1 _11784_ ( .A1(_04082_ ), .A2(_04083_ ), .A3(_04084_ ), .A4(\io_master_rid [0] ), .ZN(_04085_ ) );
AOI21_X1 _11785_ ( .A(_02167_ ), .B1(_04081_ ), .B2(_04085_ ), .ZN(_04086_ ) );
OR3_X1 _11786_ ( .A1(_04076_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .A3(_04079_ ), .ZN(_04087_ ) );
OAI21_X1 _11787_ ( .A(io_master_rvalid ), .B1(_04076_ ), .B2(_04079_ ), .ZN(_04088_ ) );
NAND2_X2 _11788_ ( .A1(_04087_ ), .A2(_04088_ ), .ZN(_04089_ ) );
AND2_X1 _11789_ ( .A1(_04086_ ), .A2(_04089_ ), .ZN(_04090_ ) );
BUF_X4 _11790_ ( .A(_04090_ ), .Z(_04091_ ) );
OR2_X1 _11791_ ( .A1(_04080_ ), .A2(io_master_rlast ), .ZN(_04092_ ) );
AND2_X1 _11792_ ( .A1(_04091_ ), .A2(_04092_ ), .ZN(_04093_ ) );
INV_X1 _11793_ ( .A(_04093_ ), .ZN(_04094_ ) );
INV_X1 _11794_ ( .A(\myifu.tmp_offset [2] ), .ZN(_04095_ ) );
NAND3_X1 _11795_ ( .A1(_04094_ ), .A2(_03903_ ), .A3(_04095_ ), .ZN(_04096_ ) );
INV_X1 _11796_ ( .A(_04096_ ), .ZN(_00315_ ) );
NOR3_X1 _11797_ ( .A1(fanout_net_5 ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00316_ ) );
AND3_X1 _11798_ ( .A1(_02312_ ), .A2(_03539_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_04097_ ) );
INV_X1 _11799_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_04098_ ) );
MUX2_X1 _11800_ ( .A(_02312_ ), .B(_04098_ ), .S(\myifu.to_reset ), .Z(_04099_ ) );
AOI211_X1 _11801_ ( .A(fanout_net_5 ), .B(_04097_ ), .C1(_04099_ ), .C2(\myifu.state [1] ), .ZN(_00317_ ) );
INV_X1 _11802_ ( .A(_02256_ ), .ZN(_04100_ ) );
NOR2_X1 _11803_ ( .A1(_02265_ ), .A2(_04100_ ), .ZN(_04101_ ) );
INV_X2 _11804_ ( .A(_04101_ ), .ZN(_04102_ ) );
BUF_X2 _11805_ ( .A(_04102_ ), .Z(_04103_ ) );
AND2_X2 _11806_ ( .A1(_02255_ ), .A2(\EX_LS_flag [2] ), .ZN(_04104_ ) );
BUF_X4 _11807_ ( .A(_04104_ ), .Z(_04105_ ) );
MUX2_X1 _11808_ ( .A(\LS_WB_waddr_csreg [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_04105_ ), .Z(_04106_ ) );
NOR2_X1 _11809_ ( .A1(_02145_ ), .A2(\EX_LS_flag [1] ), .ZN(_04107_ ) );
OR2_X1 _11810_ ( .A1(_04107_ ), .A2(_02243_ ), .ZN(_04108_ ) );
AND2_X2 _11811_ ( .A1(_02377_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_04109_ ) );
NOR2_X1 _11812_ ( .A1(_04108_ ), .A2(_04109_ ), .ZN(_04110_ ) );
BUF_X2 _11813_ ( .A(_04110_ ), .Z(_04111_ ) );
AND3_X1 _11814_ ( .A1(_04103_ ), .A2(_04106_ ), .A3(_04111_ ), .ZN(_00320_ ) );
BUF_X4 _11815_ ( .A(_02244_ ), .Z(_04112_ ) );
NOR2_X1 _11816_ ( .A1(_04101_ ), .A2(_04109_ ), .ZN(_04113_ ) );
INV_X1 _11817_ ( .A(_04113_ ), .ZN(_04114_ ) );
BUF_X4 _11818_ ( .A(_02255_ ), .Z(_04115_ ) );
NAND3_X1 _11819_ ( .A1(_04115_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_04116_ ) );
BUF_X4 _11820_ ( .A(_02145_ ), .Z(_04117_ ) );
BUF_X4 _11821_ ( .A(_04117_ ), .Z(_04118_ ) );
NAND2_X1 _11822_ ( .A1(_04118_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_04119_ ) );
AOI211_X1 _11823_ ( .A(_04112_ ), .B(_04114_ ), .C1(_04116_ ), .C2(_04119_ ), .ZN(_00321_ ) );
NAND3_X1 _11824_ ( .A1(_04115_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_04120_ ) );
NAND2_X1 _11825_ ( .A1(_04118_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_04121_ ) );
AOI211_X1 _11826_ ( .A(_04112_ ), .B(_04114_ ), .C1(_04120_ ), .C2(_04121_ ), .ZN(_00322_ ) );
NAND3_X1 _11827_ ( .A1(_04115_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_04122_ ) );
NAND2_X1 _11828_ ( .A1(_04118_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_04123_ ) );
AOI211_X1 _11829_ ( .A(_04112_ ), .B(_04114_ ), .C1(_04122_ ), .C2(_04123_ ), .ZN(_00323_ ) );
NAND3_X1 _11830_ ( .A1(_04115_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_04124_ ) );
NAND2_X1 _11831_ ( .A1(_04118_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_04125_ ) );
AOI211_X1 _11832_ ( .A(_04112_ ), .B(_04114_ ), .C1(_04124_ ), .C2(_04125_ ), .ZN(_00324_ ) );
NAND3_X1 _11833_ ( .A1(_04115_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_04126_ ) );
NAND2_X1 _11834_ ( .A1(_04118_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_04127_ ) );
AOI211_X1 _11835_ ( .A(_04112_ ), .B(_04114_ ), .C1(_04126_ ), .C2(_04127_ ), .ZN(_00325_ ) );
NAND3_X1 _11836_ ( .A1(_04115_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_04128_ ) );
NAND2_X1 _11837_ ( .A1(_04118_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_04129_ ) );
AOI211_X1 _11838_ ( .A(_04112_ ), .B(_04114_ ), .C1(_04128_ ), .C2(_04129_ ), .ZN(_00326_ ) );
NAND3_X1 _11839_ ( .A1(_04115_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_flag [2] ), .ZN(_04130_ ) );
NAND2_X1 _11840_ ( .A1(_04118_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_04131_ ) );
AOI211_X1 _11841_ ( .A(_04112_ ), .B(_04114_ ), .C1(_04130_ ), .C2(_04131_ ), .ZN(_00327_ ) );
INV_X1 _11842_ ( .A(_04112_ ), .ZN(_04132_ ) );
NOR4_X1 _11843_ ( .A1(_04118_ ), .A2(_02254_ ), .A3(\EX_LS_dest_csreg_mem [9] ), .A4(\EX_LS_flag [0] ), .ZN(_04133_ ) );
NOR2_X1 _11844_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_04134_ ) );
OAI211_X1 _11845_ ( .A(_04113_ ), .B(_04132_ ), .C1(_04133_ ), .C2(_04134_ ), .ZN(_00328_ ) );
NOR4_X1 _11846_ ( .A1(_04118_ ), .A2(_02254_ ), .A3(\EX_LS_dest_csreg_mem [8] ), .A4(\EX_LS_flag [0] ), .ZN(_04135_ ) );
NOR2_X1 _11847_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_04136_ ) );
OAI211_X1 _11848_ ( .A(_04113_ ), .B(_04132_ ), .C1(_04135_ ), .C2(_04136_ ), .ZN(_00329_ ) );
NOR4_X1 _11849_ ( .A1(_04118_ ), .A2(_02254_ ), .A3(\EX_LS_dest_csreg_mem [6] ), .A4(\EX_LS_flag [0] ), .ZN(_04137_ ) );
NOR2_X1 _11850_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_04138_ ) );
OAI211_X1 _11851_ ( .A(_04113_ ), .B(_04132_ ), .C1(_04137_ ), .C2(_04138_ ), .ZN(_00330_ ) );
NOR4_X1 _11852_ ( .A1(_04117_ ), .A2(_02254_ ), .A3(fanout_net_6 ), .A4(\EX_LS_flag [0] ), .ZN(_04139_ ) );
NOR2_X1 _11853_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_04140_ ) );
OAI211_X1 _11854_ ( .A(_04113_ ), .B(_04132_ ), .C1(_04139_ ), .C2(_04140_ ), .ZN(_00331_ ) );
INV_X1 _11855_ ( .A(\mysc.state [2] ), .ZN(_04141_ ) );
NOR2_X1 _11856_ ( .A1(_04141_ ), .A2(fanout_net_5 ), .ZN(_00339_ ) );
INV_X2 _11857_ ( .A(_03338_ ), .ZN(_04142_ ) );
NOR2_X1 _11858_ ( .A1(_03592_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _11859_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_04143_ ) );
NOR2_X1 _11860_ ( .A1(_03605_ ), .A2(\ID_EX_typ [6] ), .ZN(_04144_ ) );
AND2_X1 _11861_ ( .A1(_04144_ ), .A2(\ID_EX_typ [5] ), .ZN(_04145_ ) );
INV_X2 _11862_ ( .A(fanout_net_7 ), .ZN(_04146_ ) );
AND2_X2 _11863_ ( .A1(_04145_ ), .A2(_04146_ ), .ZN(_04147_ ) );
INV_X1 _11864_ ( .A(_04147_ ), .ZN(_04148_ ) );
INV_X1 _11865_ ( .A(\ID_EX_typ [5] ), .ZN(_04149_ ) );
BUF_X2 _11866_ ( .A(_04149_ ), .Z(_04150_ ) );
INV_X1 _11867_ ( .A(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04151_ ) );
NAND3_X1 _11868_ ( .A1(_04144_ ), .A2(_04150_ ), .A3(_04151_ ), .ZN(_04152_ ) );
AOI21_X1 _11869_ ( .A(_04143_ ), .B1(_04148_ ), .B2(_04152_ ), .ZN(_04153_ ) );
OR2_X1 _11870_ ( .A1(_03537_ ), .A2(check_assert ), .ZN(_04154_ ) );
INV_X1 _11871_ ( .A(\ID_EX_typ [6] ), .ZN(_04155_ ) );
CLKBUF_X2 _11872_ ( .A(_02187_ ), .Z(_04156_ ) );
AND4_X1 _11873_ ( .A1(\ID_EX_typ [7] ), .A2(_04155_ ), .A3(_04156_ ), .A4(IDU_valid_EXU ), .ZN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _11874_ ( .A(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_04157_ ) );
AOI211_X1 _11875_ ( .A(_04142_ ), .B(_04153_ ), .C1(_04154_ ), .C2(_04157_ ), .ZN(_00132_ ) );
CLKBUF_X2 _11876_ ( .A(_03338_ ), .Z(_04158_ ) );
AND2_X1 _11877_ ( .A1(_04158_ ), .A2(\ID_EX_rd [4] ), .ZN(_00153_ ) );
AND2_X1 _11878_ ( .A1(_04158_ ), .A2(\ID_EX_rd [3] ), .ZN(_00154_ ) );
AND2_X1 _11879_ ( .A1(_04158_ ), .A2(\ID_EX_rd [2] ), .ZN(_00155_ ) );
AND2_X1 _11880_ ( .A1(_04158_ ), .A2(\ID_EX_rd [1] ), .ZN(_00156_ ) );
AND2_X1 _11881_ ( .A1(_04158_ ), .A2(\ID_EX_rd [0] ), .ZN(_00157_ ) );
BUF_X4 _11882_ ( .A(_04142_ ), .Z(_04159_ ) );
AND2_X1 _11883_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_04160_ ) );
AND2_X1 _11884_ ( .A1(_04160_ ), .A2(\ID_EX_pc [4] ), .ZN(_04161_ ) );
AND2_X1 _11885_ ( .A1(_04161_ ), .A2(\ID_EX_pc [5] ), .ZN(_04162_ ) );
AND2_X1 _11886_ ( .A1(_04162_ ), .A2(\ID_EX_pc [6] ), .ZN(_04163_ ) );
AND2_X1 _11887_ ( .A1(_04163_ ), .A2(\ID_EX_pc [7] ), .ZN(_04164_ ) );
AND2_X1 _11888_ ( .A1(_04164_ ), .A2(\ID_EX_pc [8] ), .ZN(_04165_ ) );
AND2_X1 _11889_ ( .A1(_04165_ ), .A2(\ID_EX_pc [9] ), .ZN(_04166_ ) );
AND2_X1 _11890_ ( .A1(_04166_ ), .A2(\ID_EX_pc [10] ), .ZN(_04167_ ) );
AND2_X1 _11891_ ( .A1(_04167_ ), .A2(\ID_EX_pc [11] ), .ZN(_04168_ ) );
AND2_X1 _11892_ ( .A1(_04168_ ), .A2(\ID_EX_pc [12] ), .ZN(_04169_ ) );
AND2_X1 _11893_ ( .A1(_04169_ ), .A2(\ID_EX_pc [13] ), .ZN(_04170_ ) );
AND3_X1 _11894_ ( .A1(_04170_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_04171_ ) );
AND3_X1 _11895_ ( .A1(_04171_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_04172_ ) );
AND3_X1 _11896_ ( .A1(_04172_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_04173_ ) );
AND3_X1 _11897_ ( .A1(_04173_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_04174_ ) );
AND3_X1 _11898_ ( .A1(_04174_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_04175_ ) );
AND3_X1 _11899_ ( .A1(_04175_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_04176_ ) );
AND3_X1 _11900_ ( .A1(_04176_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_04177_ ) );
NAND3_X1 _11901_ ( .A1(_04177_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_04178_ ) );
XNOR2_X1 _11902_ ( .A(_04178_ ), .B(\ID_EX_pc [30] ), .ZN(_04179_ ) );
XOR2_X1 _11903_ ( .A(\ID_EX_pc [25] ), .B(\ID_EX_imm [25] ), .Z(_04180_ ) );
XOR2_X1 _11904_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_04181_ ) );
NOR2_X1 _11905_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04182_ ) );
XOR2_X1 _11906_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_04183_ ) );
XOR2_X1 _11907_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_04184_ ) );
XOR2_X1 _11908_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_04185_ ) );
AND2_X1 _11909_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_04186_ ) );
AND2_X1 _11910_ ( .A1(_04185_ ), .A2(_04186_ ), .ZN(_04187_ ) );
AND2_X1 _11911_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_04188_ ) );
OAI21_X1 _11912_ ( .A(_04184_ ), .B1(_04187_ ), .B2(_04188_ ), .ZN(_04189_ ) );
NAND2_X1 _11913_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_04190_ ) );
INV_X1 _11914_ ( .A(\ID_EX_pc [3] ), .ZN(_04191_ ) );
AOI22_X1 _11915_ ( .A1(_04189_ ), .A2(_04190_ ), .B1(_04191_ ), .B2(_02911_ ), .ZN(_04192_ ) );
AND2_X1 _11916_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_04193_ ) );
OAI21_X1 _11917_ ( .A(_04183_ ), .B1(_04192_ ), .B2(_04193_ ), .ZN(_04194_ ) );
NAND2_X1 _11918_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_04195_ ) );
NAND2_X1 _11919_ ( .A1(_04194_ ), .A2(_04195_ ), .ZN(_04196_ ) );
OAI21_X1 _11920_ ( .A(_04196_ ), .B1(\ID_EX_pc [5] ), .B2(\ID_EX_imm [5] ), .ZN(_04197_ ) );
AND2_X1 _11921_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_04198_ ) );
INV_X1 _11922_ ( .A(_04198_ ), .ZN(_04199_ ) );
NAND2_X1 _11923_ ( .A1(_04197_ ), .A2(_04199_ ), .ZN(_04200_ ) );
XOR2_X1 _11924_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_04201_ ) );
NAND2_X1 _11925_ ( .A1(_04200_ ), .A2(_04201_ ), .ZN(_04202_ ) );
NAND2_X1 _11926_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_04203_ ) );
AOI21_X1 _11927_ ( .A(_04182_ ), .B1(_04202_ ), .B2(_04203_ ), .ZN(_04204_ ) );
AND2_X1 _11928_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04205_ ) );
OR2_X1 _11929_ ( .A1(_04204_ ), .A2(_04205_ ), .ZN(_04206_ ) );
XOR2_X1 _11930_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_04207_ ) );
XOR2_X1 _11931_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_04208_ ) );
AND2_X1 _11932_ ( .A1(_04207_ ), .A2(_04208_ ), .ZN(_04209_ ) );
XOR2_X1 _11933_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_04210_ ) );
XOR2_X1 _11934_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_04211_ ) );
AND2_X1 _11935_ ( .A1(_04210_ ), .A2(_04211_ ), .ZN(_04212_ ) );
AND3_X1 _11936_ ( .A1(_04206_ ), .A2(_04209_ ), .A3(_04212_ ), .ZN(_04213_ ) );
AND2_X1 _11937_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_04214_ ) );
AND2_X1 _11938_ ( .A1(_04207_ ), .A2(_04214_ ), .ZN(_04215_ ) );
AOI21_X1 _11939_ ( .A(_04215_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_04216_ ) );
AND2_X1 _11940_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_04217_ ) );
AND2_X1 _11941_ ( .A1(_04211_ ), .A2(_04217_ ), .ZN(_04218_ ) );
AOI21_X1 _11942_ ( .A(_04218_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_04219_ ) );
INV_X1 _11943_ ( .A(_04209_ ), .ZN(_04220_ ) );
OAI21_X1 _11944_ ( .A(_04216_ ), .B1(_04219_ ), .B2(_04220_ ), .ZN(_04221_ ) );
OR2_X1 _11945_ ( .A1(_04213_ ), .A2(_04221_ ), .ZN(_04222_ ) );
XOR2_X1 _11946_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_04223_ ) );
XOR2_X1 _11947_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_04224_ ) );
AND2_X1 _11948_ ( .A1(_04223_ ), .A2(_04224_ ), .ZN(_04225_ ) );
XOR2_X1 _11949_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_04226_ ) );
INV_X1 _11950_ ( .A(_04226_ ), .ZN(_04227_ ) );
XNOR2_X1 _11951_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .ZN(_04228_ ) );
NOR2_X1 _11952_ ( .A1(_04227_ ), .A2(_04228_ ), .ZN(_04229_ ) );
AND3_X1 _11953_ ( .A1(_04222_ ), .A2(_04225_ ), .A3(_04229_ ), .ZN(_04230_ ) );
AND2_X1 _11954_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04231_ ) );
AND2_X1 _11955_ ( .A1(_04223_ ), .A2(_04231_ ), .ZN(_04232_ ) );
AOI21_X1 _11956_ ( .A(_04232_ ), .B1(\ID_EX_pc [15] ), .B2(\ID_EX_imm [15] ), .ZN(_04233_ ) );
INV_X1 _11957_ ( .A(_04225_ ), .ZN(_04234_ ) );
NAND2_X1 _11958_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_04235_ ) );
NOR2_X1 _11959_ ( .A1(_04228_ ), .A2(_04235_ ), .ZN(_04236_ ) );
AOI21_X1 _11960_ ( .A(_04236_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_04237_ ) );
OAI21_X1 _11961_ ( .A(_04233_ ), .B1(_04234_ ), .B2(_04237_ ), .ZN(_04238_ ) );
OR2_X1 _11962_ ( .A1(_04230_ ), .A2(_04238_ ), .ZN(_04239_ ) );
XOR2_X1 _11963_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_04240_ ) );
XOR2_X1 _11964_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_04241_ ) );
AND2_X1 _11965_ ( .A1(_04240_ ), .A2(_04241_ ), .ZN(_04242_ ) );
XOR2_X1 _11966_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_04243_ ) );
XOR2_X1 _11967_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_04244_ ) );
AND2_X1 _11968_ ( .A1(_04243_ ), .A2(_04244_ ), .ZN(_04245_ ) );
AND3_X1 _11969_ ( .A1(_04239_ ), .A2(_04242_ ), .A3(_04245_ ), .ZN(_04246_ ) );
AND2_X1 _11970_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_04247_ ) );
AND2_X1 _11971_ ( .A1(_04240_ ), .A2(_04247_ ), .ZN(_04248_ ) );
AOI21_X1 _11972_ ( .A(_04248_ ), .B1(\ID_EX_pc [19] ), .B2(\ID_EX_imm [19] ), .ZN(_04249_ ) );
AND2_X1 _11973_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_04250_ ) );
AND2_X1 _11974_ ( .A1(_04244_ ), .A2(_04250_ ), .ZN(_04251_ ) );
AOI21_X1 _11975_ ( .A(_04251_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_04252_ ) );
INV_X1 _11976_ ( .A(_04242_ ), .ZN(_04253_ ) );
OAI21_X1 _11977_ ( .A(_04249_ ), .B1(_04252_ ), .B2(_04253_ ), .ZN(_04254_ ) );
OR2_X1 _11978_ ( .A1(_04246_ ), .A2(_04254_ ), .ZN(_04255_ ) );
XOR2_X1 _11979_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_04256_ ) );
XOR2_X1 _11980_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_04257_ ) );
AND2_X1 _11981_ ( .A1(_04256_ ), .A2(_04257_ ), .ZN(_04258_ ) );
XOR2_X1 _11982_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_04259_ ) );
XOR2_X1 _11983_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_04260_ ) );
AND2_X1 _11984_ ( .A1(_04259_ ), .A2(_04260_ ), .ZN(_04261_ ) );
AND3_X1 _11985_ ( .A1(_04255_ ), .A2(_04258_ ), .A3(_04261_ ), .ZN(_04262_ ) );
AND2_X1 _11986_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_04263_ ) );
AND2_X1 _11987_ ( .A1(_04256_ ), .A2(_04263_ ), .ZN(_04264_ ) );
AOI21_X1 _11988_ ( .A(_04264_ ), .B1(\ID_EX_pc [23] ), .B2(\ID_EX_imm [23] ), .ZN(_04265_ ) );
AND2_X1 _11989_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_04266_ ) );
AND2_X1 _11990_ ( .A1(_04259_ ), .A2(_04266_ ), .ZN(_04267_ ) );
AOI21_X1 _11991_ ( .A(_04267_ ), .B1(\ID_EX_pc [21] ), .B2(\ID_EX_imm [21] ), .ZN(_04268_ ) );
INV_X1 _11992_ ( .A(_04258_ ), .ZN(_04269_ ) );
OAI21_X1 _11993_ ( .A(_04265_ ), .B1(_04268_ ), .B2(_04269_ ), .ZN(_04270_ ) );
OAI211_X1 _11994_ ( .A(_04180_ ), .B(_04181_ ), .C1(_04262_ ), .C2(_04270_ ), .ZN(_04271_ ) );
AND2_X1 _11995_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_04272_ ) );
AND2_X1 _11996_ ( .A1(_04180_ ), .A2(_04272_ ), .ZN(_04273_ ) );
AOI21_X1 _11997_ ( .A(_04273_ ), .B1(\ID_EX_pc [25] ), .B2(\ID_EX_imm [25] ), .ZN(_04274_ ) );
NAND2_X1 _11998_ ( .A1(_04271_ ), .A2(_04274_ ), .ZN(_04275_ ) );
XOR2_X1 _11999_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_04276_ ) );
XOR2_X1 _12000_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_04277_ ) );
NAND3_X1 _12001_ ( .A1(_04275_ ), .A2(_04276_ ), .A3(_04277_ ), .ZN(_04278_ ) );
AND3_X1 _12002_ ( .A1(_04276_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_04279_ ) );
AOI21_X1 _12003_ ( .A(_04279_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_04280_ ) );
NAND2_X1 _12004_ ( .A1(_04278_ ), .A2(_04280_ ), .ZN(_04281_ ) );
XOR2_X1 _12005_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_04282_ ) );
NAND2_X1 _12006_ ( .A1(_04281_ ), .A2(_04282_ ), .ZN(_04283_ ) );
NAND2_X1 _12007_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_04284_ ) );
INV_X1 _12008_ ( .A(\ID_EX_pc [29] ), .ZN(_04285_ ) );
AOI22_X1 _12009_ ( .A1(_04283_ ), .A2(_04284_ ), .B1(_04285_ ), .B2(_02426_ ), .ZN(_04286_ ) );
AND2_X1 _12010_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_04287_ ) );
OR2_X1 _12011_ ( .A1(_04286_ ), .A2(_04287_ ), .ZN(_04288_ ) );
XOR2_X1 _12012_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_04289_ ) );
XOR2_X1 _12013_ ( .A(_04288_ ), .B(_04289_ ), .Z(_04290_ ) );
NOR2_X1 _12014_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_7 ), .ZN(_04291_ ) );
AND2_X1 _12015_ ( .A1(_04291_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04292_ ) );
OAI21_X2 _12016_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02385_ ), .B2(\ID_EX_rs2 [1] ), .ZN(_04293_ ) );
AOI211_X2 _12017_ ( .A(_04293_ ), .B(_02454_ ), .C1(_02385_ ), .C2(\ID_EX_rs2 [1] ), .ZN(_04294_ ) );
XNOR2_X1 _12018_ ( .A(\EX_LS_dest_reg [3] ), .B(\ID_EX_rs2 [3] ), .ZN(_04295_ ) );
XNOR2_X1 _12019_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_04296_ ) );
XNOR2_X1 _12020_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_04297_ ) );
XNOR2_X1 _12021_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_04298_ ) );
AND4_X4 _12022_ ( .A1(_04295_ ), .A2(_04296_ ), .A3(_04297_ ), .A4(_04298_ ), .ZN(_04299_ ) );
NAND2_X2 _12023_ ( .A1(_04294_ ), .A2(_04299_ ), .ZN(_04300_ ) );
BUF_X8 _12024_ ( .A(_04300_ ), .Z(_04301_ ) );
BUF_X16 _12025_ ( .A(_04301_ ), .Z(_04302_ ) );
BUF_X4 _12026_ ( .A(_04302_ ), .Z(_04303_ ) );
BUF_X8 _12027_ ( .A(_02379_ ), .Z(_04304_ ) );
BUF_X16 _12028_ ( .A(_04304_ ), .Z(_04305_ ) );
BUF_X4 _12029_ ( .A(_04305_ ), .Z(_04306_ ) );
OR3_X1 _12030_ ( .A1(_04303_ ), .A2(\EX_LS_result_reg [16] ), .A3(_04306_ ), .ZN(_04307_ ) );
INV_X1 _12031_ ( .A(fanout_net_41 ), .ZN(_04308_ ) );
BUF_X4 _12032_ ( .A(_04308_ ), .Z(_04309_ ) );
BUF_X4 _12033_ ( .A(_04309_ ), .Z(_04310_ ) );
BUF_X4 _12034_ ( .A(_04310_ ), .Z(_04311_ ) );
OR2_X1 _12035_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[4][16] ), .ZN(_04312_ ) );
INV_X2 _12036_ ( .A(fanout_net_38 ), .ZN(_04313_ ) );
BUF_X4 _12037_ ( .A(_04313_ ), .Z(_04314_ ) );
BUF_X4 _12038_ ( .A(_04314_ ), .Z(_04315_ ) );
BUF_X4 _12039_ ( .A(_04315_ ), .Z(_04316_ ) );
BUF_X4 _12040_ ( .A(_04316_ ), .Z(_04317_ ) );
BUF_X4 _12041_ ( .A(_04317_ ), .Z(_04318_ ) );
INV_X32 _12042_ ( .A(fanout_net_30 ), .ZN(_04319_ ) );
BUF_X32 _12043_ ( .A(_04319_ ), .Z(_04320_ ) );
BUF_X4 _12044_ ( .A(_04320_ ), .Z(_04321_ ) );
BUF_X8 _12045_ ( .A(_04321_ ), .Z(_04322_ ) );
BUF_X2 _12046_ ( .A(_04322_ ), .Z(_04323_ ) );
BUF_X2 _12047_ ( .A(_04323_ ), .Z(_04324_ ) );
OAI211_X1 _12048_ ( .A(_04312_ ), .B(_04318_ ), .C1(_04324_ ), .C2(\myreg.Reg[5][16] ), .ZN(_04325_ ) );
OR2_X1 _12049_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[6][16] ), .ZN(_04326_ ) );
OAI211_X1 _12050_ ( .A(_04326_ ), .B(fanout_net_38 ), .C1(_04324_ ), .C2(\myreg.Reg[7][16] ), .ZN(_04327_ ) );
NAND3_X1 _12051_ ( .A1(_04325_ ), .A2(_04327_ ), .A3(fanout_net_40 ), .ZN(_04328_ ) );
MUX2_X1 _12052_ ( .A(\myreg.Reg[2][16] ), .B(\myreg.Reg[3][16] ), .S(fanout_net_30 ), .Z(_04329_ ) );
MUX2_X1 _12053_ ( .A(\myreg.Reg[0][16] ), .B(\myreg.Reg[1][16] ), .S(fanout_net_30 ), .Z(_04330_ ) );
BUF_X4 _12054_ ( .A(_04315_ ), .Z(_04331_ ) );
BUF_X4 _12055_ ( .A(_04331_ ), .Z(_04332_ ) );
MUX2_X1 _12056_ ( .A(_04329_ ), .B(_04330_ ), .S(_04332_ ), .Z(_04333_ ) );
OAI211_X1 _12057_ ( .A(_04311_ ), .B(_04328_ ), .C1(_04333_ ), .C2(fanout_net_40 ), .ZN(_04334_ ) );
INV_X2 _12058_ ( .A(fanout_net_40 ), .ZN(_04335_ ) );
BUF_X4 _12059_ ( .A(_04335_ ), .Z(_04336_ ) );
BUF_X4 _12060_ ( .A(_04336_ ), .Z(_04337_ ) );
BUF_X4 _12061_ ( .A(_04337_ ), .Z(_04338_ ) );
BUF_X2 _12062_ ( .A(_04322_ ), .Z(_04339_ ) );
BUF_X2 _12063_ ( .A(_04339_ ), .Z(_04340_ ) );
NOR2_X1 _12064_ ( .A1(_04340_ ), .A2(\myreg.Reg[11][16] ), .ZN(_04341_ ) );
OAI21_X1 _12065_ ( .A(fanout_net_38 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][16] ), .ZN(_04342_ ) );
NOR2_X1 _12066_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][16] ), .ZN(_04343_ ) );
OAI21_X1 _12067_ ( .A(_04332_ ), .B1(_04340_ ), .B2(\myreg.Reg[9][16] ), .ZN(_04344_ ) );
OAI221_X1 _12068_ ( .A(_04338_ ), .B1(_04341_ ), .B2(_04342_ ), .C1(_04343_ ), .C2(_04344_ ), .ZN(_04345_ ) );
MUX2_X1 _12069_ ( .A(\myreg.Reg[12][16] ), .B(\myreg.Reg[13][16] ), .S(fanout_net_30 ), .Z(_04346_ ) );
MUX2_X1 _12070_ ( .A(\myreg.Reg[14][16] ), .B(\myreg.Reg[15][16] ), .S(fanout_net_30 ), .Z(_04347_ ) );
MUX2_X1 _12071_ ( .A(_04346_ ), .B(_04347_ ), .S(fanout_net_38 ), .Z(_04348_ ) );
BUF_X4 _12072_ ( .A(_04338_ ), .Z(_04349_ ) );
OAI211_X1 _12073_ ( .A(fanout_net_41 ), .B(_04345_ ), .C1(_04348_ ), .C2(_04349_ ), .ZN(_04350_ ) );
OAI211_X1 _12074_ ( .A(_04334_ ), .B(_04350_ ), .C1(_04303_ ), .C2(_04306_ ), .ZN(_04351_ ) );
NAND2_X1 _12075_ ( .A1(_04307_ ), .A2(_04351_ ), .ZN(_04352_ ) );
XOR2_X1 _12076_ ( .A(_02709_ ), .B(_04352_ ), .Z(_04353_ ) );
BUF_X16 _12077_ ( .A(_04305_ ), .Z(_04354_ ) );
OR3_X1 _12078_ ( .A1(_04303_ ), .A2(\EX_LS_result_reg [17] ), .A3(_04354_ ), .ZN(_04355_ ) );
OR2_X1 _12079_ ( .A1(_04339_ ), .A2(\myreg.Reg[1][17] ), .ZN(_04356_ ) );
OAI211_X1 _12080_ ( .A(_04356_ ), .B(_04317_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[0][17] ), .ZN(_04357_ ) );
OR2_X1 _12081_ ( .A1(_04339_ ), .A2(\myreg.Reg[3][17] ), .ZN(_04358_ ) );
OAI211_X1 _12082_ ( .A(_04358_ ), .B(fanout_net_38 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[2][17] ), .ZN(_04359_ ) );
NAND3_X1 _12083_ ( .A1(_04357_ ), .A2(_04359_ ), .A3(_04338_ ), .ZN(_04360_ ) );
MUX2_X1 _12084_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_30 ), .Z(_04361_ ) );
MUX2_X1 _12085_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_30 ), .Z(_04362_ ) );
MUX2_X1 _12086_ ( .A(_04361_ ), .B(_04362_ ), .S(_04317_ ), .Z(_04363_ ) );
OAI211_X1 _12087_ ( .A(_04311_ ), .B(_04360_ ), .C1(_04363_ ), .C2(_04349_ ), .ZN(_04364_ ) );
OR2_X1 _12088_ ( .A1(_04339_ ), .A2(\myreg.Reg[15][17] ), .ZN(_04365_ ) );
OAI211_X1 _12089_ ( .A(_04365_ ), .B(fanout_net_38 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[14][17] ), .ZN(_04366_ ) );
OR2_X1 _12090_ ( .A1(_04339_ ), .A2(\myreg.Reg[13][17] ), .ZN(_04367_ ) );
OAI211_X1 _12091_ ( .A(_04367_ ), .B(_04317_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[12][17] ), .ZN(_04368_ ) );
NAND3_X1 _12092_ ( .A1(_04366_ ), .A2(_04368_ ), .A3(fanout_net_40 ), .ZN(_04369_ ) );
MUX2_X1 _12093_ ( .A(\myreg.Reg[8][17] ), .B(\myreg.Reg[9][17] ), .S(fanout_net_30 ), .Z(_04370_ ) );
MUX2_X1 _12094_ ( .A(\myreg.Reg[10][17] ), .B(\myreg.Reg[11][17] ), .S(fanout_net_30 ), .Z(_04371_ ) );
MUX2_X1 _12095_ ( .A(_04370_ ), .B(_04371_ ), .S(fanout_net_38 ), .Z(_04372_ ) );
OAI211_X1 _12096_ ( .A(fanout_net_41 ), .B(_04369_ ), .C1(_04372_ ), .C2(fanout_net_40 ), .ZN(_04373_ ) );
OAI211_X1 _12097_ ( .A(_04364_ ), .B(_04373_ ), .C1(_04303_ ), .C2(_04306_ ), .ZN(_04374_ ) );
NAND2_X1 _12098_ ( .A1(_04355_ ), .A2(_04374_ ), .ZN(_04375_ ) );
AND2_X1 _12099_ ( .A1(_02684_ ), .A2(_04375_ ), .ZN(_04376_ ) );
NOR2_X1 _12100_ ( .A1(_02684_ ), .A2(_04375_ ), .ZN(_04377_ ) );
NOR2_X1 _12101_ ( .A1(_04376_ ), .A2(_04377_ ), .ZN(_04378_ ) );
AND2_X1 _12102_ ( .A1(_04353_ ), .A2(_04378_ ), .ZN(_04379_ ) );
AND2_X4 _12103_ ( .A1(_02638_ ), .A2(_02658_ ), .ZN(_04380_ ) );
OR3_X2 _12104_ ( .A1(_04302_ ), .A2(\EX_LS_result_reg [19] ), .A3(_04305_ ), .ZN(_04381_ ) );
OR2_X1 _12105_ ( .A1(_04322_ ), .A2(\myreg.Reg[5][19] ), .ZN(_04382_ ) );
OAI211_X1 _12106_ ( .A(_04382_ ), .B(_04331_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[4][19] ), .ZN(_04383_ ) );
OR2_X1 _12107_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[6][19] ), .ZN(_04384_ ) );
OAI211_X1 _12108_ ( .A(_04384_ ), .B(fanout_net_38 ), .C1(_04339_ ), .C2(\myreg.Reg[7][19] ), .ZN(_04385_ ) );
NAND3_X1 _12109_ ( .A1(_04383_ ), .A2(fanout_net_40 ), .A3(_04385_ ), .ZN(_04386_ ) );
MUX2_X1 _12110_ ( .A(\myreg.Reg[2][19] ), .B(\myreg.Reg[3][19] ), .S(fanout_net_30 ), .Z(_04387_ ) );
MUX2_X1 _12111_ ( .A(\myreg.Reg[0][19] ), .B(\myreg.Reg[1][19] ), .S(fanout_net_30 ), .Z(_04388_ ) );
MUX2_X1 _12112_ ( .A(_04387_ ), .B(_04388_ ), .S(_04316_ ), .Z(_04389_ ) );
OAI211_X1 _12113_ ( .A(_04310_ ), .B(_04386_ ), .C1(_04389_ ), .C2(fanout_net_40 ), .ZN(_04390_ ) );
BUF_X2 _12114_ ( .A(_04319_ ), .Z(_04391_ ) );
BUF_X2 _12115_ ( .A(_04391_ ), .Z(_04392_ ) );
BUF_X2 _12116_ ( .A(_04392_ ), .Z(_04393_ ) );
NOR2_X1 _12117_ ( .A1(_04393_ ), .A2(\myreg.Reg[11][19] ), .ZN(_04394_ ) );
OAI21_X1 _12118_ ( .A(fanout_net_38 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][19] ), .ZN(_04395_ ) );
NOR2_X1 _12119_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][19] ), .ZN(_04396_ ) );
OAI21_X1 _12120_ ( .A(_04316_ ), .B1(_04393_ ), .B2(\myreg.Reg[9][19] ), .ZN(_04397_ ) );
OAI221_X1 _12121_ ( .A(_04337_ ), .B1(_04394_ ), .B2(_04395_ ), .C1(_04396_ ), .C2(_04397_ ), .ZN(_04398_ ) );
MUX2_X1 _12122_ ( .A(\myreg.Reg[12][19] ), .B(\myreg.Reg[13][19] ), .S(fanout_net_30 ), .Z(_04399_ ) );
MUX2_X1 _12123_ ( .A(\myreg.Reg[14][19] ), .B(\myreg.Reg[15][19] ), .S(fanout_net_30 ), .Z(_04400_ ) );
MUX2_X1 _12124_ ( .A(_04399_ ), .B(_04400_ ), .S(fanout_net_38 ), .Z(_04401_ ) );
BUF_X4 _12125_ ( .A(_04337_ ), .Z(_04402_ ) );
OAI211_X1 _12126_ ( .A(fanout_net_41 ), .B(_04398_ ), .C1(_04401_ ), .C2(_04402_ ), .ZN(_04403_ ) );
BUF_X16 _12127_ ( .A(_04302_ ), .Z(_04404_ ) );
OAI211_X2 _12128_ ( .A(_04390_ ), .B(_04403_ ), .C1(_04404_ ), .C2(_04354_ ), .ZN(_04405_ ) );
NAND2_X1 _12129_ ( .A1(_04381_ ), .A2(_04405_ ), .ZN(_04406_ ) );
INV_X1 _12130_ ( .A(_04406_ ), .ZN(_04407_ ) );
XNOR2_X1 _12131_ ( .A(_04380_ ), .B(_04407_ ), .ZN(_04408_ ) );
OR3_X4 _12132_ ( .A1(_04404_ ), .A2(\EX_LS_result_reg [18] ), .A3(_04354_ ), .ZN(_04409_ ) );
OR2_X1 _12133_ ( .A1(_04322_ ), .A2(\myreg.Reg[1][18] ), .ZN(_04410_ ) );
OAI211_X1 _12134_ ( .A(_04410_ ), .B(_04331_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[0][18] ), .ZN(_04411_ ) );
OR2_X1 _12135_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[2][18] ), .ZN(_04412_ ) );
OAI211_X1 _12136_ ( .A(_04412_ ), .B(fanout_net_38 ), .C1(_04339_ ), .C2(\myreg.Reg[3][18] ), .ZN(_04413_ ) );
NAND3_X1 _12137_ ( .A1(_04411_ ), .A2(_04402_ ), .A3(_04413_ ), .ZN(_04414_ ) );
MUX2_X1 _12138_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_30 ), .Z(_04415_ ) );
MUX2_X1 _12139_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_30 ), .Z(_04416_ ) );
MUX2_X1 _12140_ ( .A(_04415_ ), .B(_04416_ ), .S(_04331_ ), .Z(_04417_ ) );
OAI211_X1 _12141_ ( .A(_04310_ ), .B(_04414_ ), .C1(_04417_ ), .C2(_04338_ ), .ZN(_04418_ ) );
OR2_X1 _12142_ ( .A1(_04322_ ), .A2(\myreg.Reg[13][18] ), .ZN(_04419_ ) );
OAI211_X1 _12143_ ( .A(_04419_ ), .B(_04331_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[12][18] ), .ZN(_04420_ ) );
OR2_X1 _12144_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][18] ), .ZN(_04421_ ) );
OAI211_X1 _12145_ ( .A(_04421_ ), .B(fanout_net_38 ), .C1(_04339_ ), .C2(\myreg.Reg[15][18] ), .ZN(_04422_ ) );
NAND3_X1 _12146_ ( .A1(_04420_ ), .A2(fanout_net_40 ), .A3(_04422_ ), .ZN(_04423_ ) );
MUX2_X1 _12147_ ( .A(\myreg.Reg[8][18] ), .B(\myreg.Reg[9][18] ), .S(fanout_net_31 ), .Z(_04424_ ) );
MUX2_X1 _12148_ ( .A(\myreg.Reg[10][18] ), .B(\myreg.Reg[11][18] ), .S(fanout_net_31 ), .Z(_04425_ ) );
MUX2_X1 _12149_ ( .A(_04424_ ), .B(_04425_ ), .S(fanout_net_38 ), .Z(_04426_ ) );
OAI211_X1 _12150_ ( .A(fanout_net_41 ), .B(_04423_ ), .C1(_04426_ ), .C2(fanout_net_40 ), .ZN(_04427_ ) );
OAI211_X2 _12151_ ( .A(_04418_ ), .B(_04427_ ), .C1(_04404_ ), .C2(_04354_ ), .ZN(_04428_ ) );
NAND2_X1 _12152_ ( .A1(_04409_ ), .A2(_04428_ ), .ZN(_04429_ ) );
INV_X1 _12153_ ( .A(_04429_ ), .ZN(_04430_ ) );
XNOR2_X1 _12154_ ( .A(_02635_ ), .B(_04430_ ), .ZN(_04431_ ) );
AND3_X1 _12155_ ( .A1(_04379_ ), .A2(_04408_ ), .A3(_04431_ ), .ZN(_04432_ ) );
INV_X1 _12156_ ( .A(_04432_ ), .ZN(_04433_ ) );
OR3_X2 _12157_ ( .A1(_04302_ ), .A2(\EX_LS_result_reg [22] ), .A3(_04305_ ), .ZN(_04434_ ) );
OR2_X2 _12158_ ( .A1(_04322_ ), .A2(\myreg.Reg[5][22] ), .ZN(_04435_ ) );
OAI211_X1 _12159_ ( .A(_04435_ ), .B(_04316_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[4][22] ), .ZN(_04436_ ) );
OR2_X1 _12160_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[6][22] ), .ZN(_04437_ ) );
OAI211_X1 _12161_ ( .A(_04437_ ), .B(fanout_net_38 ), .C1(_04393_ ), .C2(\myreg.Reg[7][22] ), .ZN(_04438_ ) );
NAND3_X1 _12162_ ( .A1(_04436_ ), .A2(fanout_net_40 ), .A3(_04438_ ), .ZN(_04439_ ) );
MUX2_X1 _12163_ ( .A(\myreg.Reg[2][22] ), .B(\myreg.Reg[3][22] ), .S(fanout_net_31 ), .Z(_04440_ ) );
MUX2_X1 _12164_ ( .A(\myreg.Reg[0][22] ), .B(\myreg.Reg[1][22] ), .S(fanout_net_31 ), .Z(_04441_ ) );
MUX2_X1 _12165_ ( .A(_04440_ ), .B(_04441_ ), .S(_04316_ ), .Z(_04442_ ) );
OAI211_X1 _12166_ ( .A(_04310_ ), .B(_04439_ ), .C1(_04442_ ), .C2(fanout_net_40 ), .ZN(_04443_ ) );
NOR2_X1 _12167_ ( .A1(_04322_ ), .A2(\myreg.Reg[11][22] ), .ZN(_04444_ ) );
OAI21_X1 _12168_ ( .A(fanout_net_38 ), .B1(fanout_net_31 ), .B2(\myreg.Reg[10][22] ), .ZN(_04445_ ) );
NOR2_X1 _12169_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][22] ), .ZN(_04446_ ) );
OAI21_X1 _12170_ ( .A(_04315_ ), .B1(_04322_ ), .B2(\myreg.Reg[9][22] ), .ZN(_04447_ ) );
OAI221_X1 _12171_ ( .A(_04337_ ), .B1(_04444_ ), .B2(_04445_ ), .C1(_04446_ ), .C2(_04447_ ), .ZN(_04448_ ) );
MUX2_X1 _12172_ ( .A(\myreg.Reg[12][22] ), .B(\myreg.Reg[13][22] ), .S(fanout_net_31 ), .Z(_04449_ ) );
MUX2_X1 _12173_ ( .A(\myreg.Reg[14][22] ), .B(\myreg.Reg[15][22] ), .S(fanout_net_31 ), .Z(_04450_ ) );
MUX2_X1 _12174_ ( .A(_04449_ ), .B(_04450_ ), .S(fanout_net_38 ), .Z(_04451_ ) );
OAI211_X1 _12175_ ( .A(fanout_net_41 ), .B(_04448_ ), .C1(_04451_ ), .C2(_04402_ ), .ZN(_04452_ ) );
OAI211_X2 _12176_ ( .A(_04443_ ), .B(_04452_ ), .C1(_04404_ ), .C2(_04354_ ), .ZN(_04453_ ) );
NAND2_X2 _12177_ ( .A1(_04434_ ), .A2(_04453_ ), .ZN(_04454_ ) );
INV_X1 _12178_ ( .A(_04454_ ), .ZN(_04455_ ) );
XNOR2_X1 _12179_ ( .A(_02535_ ), .B(_04455_ ), .ZN(_04456_ ) );
INV_X1 _12180_ ( .A(\EX_LS_result_reg [23] ), .ZN(_04457_ ) );
OR3_X4 _12181_ ( .A1(_04302_ ), .A2(_04457_ ), .A3(_04305_ ), .ZN(_04458_ ) );
OR2_X1 _12182_ ( .A1(_04392_ ), .A2(\myreg.Reg[1][23] ), .ZN(_04459_ ) );
OAI211_X1 _12183_ ( .A(_04459_ ), .B(_04316_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[0][23] ), .ZN(_04460_ ) );
OR2_X1 _12184_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][23] ), .ZN(_04461_ ) );
OAI211_X1 _12185_ ( .A(_04461_ ), .B(fanout_net_38 ), .C1(_04393_ ), .C2(\myreg.Reg[3][23] ), .ZN(_04462_ ) );
NAND3_X1 _12186_ ( .A1(_04460_ ), .A2(_04337_ ), .A3(_04462_ ), .ZN(_04463_ ) );
MUX2_X1 _12187_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_31 ), .Z(_04464_ ) );
MUX2_X1 _12188_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_31 ), .Z(_04465_ ) );
MUX2_X1 _12189_ ( .A(_04464_ ), .B(_04465_ ), .S(_04315_ ), .Z(_04466_ ) );
OAI211_X1 _12190_ ( .A(_04310_ ), .B(_04463_ ), .C1(_04466_ ), .C2(_04402_ ), .ZN(_04467_ ) );
OR2_X1 _12191_ ( .A1(_04392_ ), .A2(\myreg.Reg[13][23] ), .ZN(_04468_ ) );
OAI211_X1 _12192_ ( .A(_04468_ ), .B(_04315_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[12][23] ), .ZN(_04469_ ) );
OR2_X1 _12193_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][23] ), .ZN(_04470_ ) );
OAI211_X1 _12194_ ( .A(_04470_ ), .B(fanout_net_38 ), .C1(_04322_ ), .C2(\myreg.Reg[15][23] ), .ZN(_04471_ ) );
NAND3_X1 _12195_ ( .A1(_04469_ ), .A2(fanout_net_40 ), .A3(_04471_ ), .ZN(_04472_ ) );
MUX2_X1 _12196_ ( .A(\myreg.Reg[8][23] ), .B(\myreg.Reg[9][23] ), .S(fanout_net_31 ), .Z(_04473_ ) );
MUX2_X1 _12197_ ( .A(\myreg.Reg[10][23] ), .B(\myreg.Reg[11][23] ), .S(fanout_net_31 ), .Z(_04474_ ) );
MUX2_X1 _12198_ ( .A(_04473_ ), .B(_04474_ ), .S(fanout_net_38 ), .Z(_04475_ ) );
OAI211_X1 _12199_ ( .A(fanout_net_41 ), .B(_04472_ ), .C1(_04475_ ), .C2(fanout_net_40 ), .ZN(_04476_ ) );
NAND2_X1 _12200_ ( .A1(_04467_ ), .A2(_04476_ ), .ZN(_04477_ ) );
OAI21_X2 _12201_ ( .A(_04477_ ), .B1(_04354_ ), .B2(_04404_ ), .ZN(_04478_ ) );
AND2_X2 _12202_ ( .A1(_04458_ ), .A2(_04478_ ), .ZN(_04479_ ) );
INV_X1 _12203_ ( .A(_04479_ ), .ZN(_04480_ ) );
XNOR2_X1 _12204_ ( .A(_04480_ ), .B(_02561_ ), .ZN(_04481_ ) );
AND2_X1 _12205_ ( .A1(_04456_ ), .A2(_04481_ ), .ZN(_04482_ ) );
OR3_X4 _12206_ ( .A1(_04404_ ), .A2(\EX_LS_result_reg [20] ), .A3(_04354_ ), .ZN(_04483_ ) );
OR2_X1 _12207_ ( .A1(_04393_ ), .A2(\myreg.Reg[11][20] ), .ZN(_04484_ ) );
OAI211_X1 _12208_ ( .A(_04484_ ), .B(fanout_net_38 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[10][20] ), .ZN(_04485_ ) );
OR2_X1 _12209_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][20] ), .ZN(_04486_ ) );
OAI211_X1 _12210_ ( .A(_04486_ ), .B(_04317_ ), .C1(_04323_ ), .C2(\myreg.Reg[9][20] ), .ZN(_04487_ ) );
NAND3_X1 _12211_ ( .A1(_04485_ ), .A2(_04402_ ), .A3(_04487_ ), .ZN(_04488_ ) );
MUX2_X1 _12212_ ( .A(\myreg.Reg[14][20] ), .B(\myreg.Reg[15][20] ), .S(fanout_net_31 ), .Z(_04489_ ) );
MUX2_X1 _12213_ ( .A(\myreg.Reg[12][20] ), .B(\myreg.Reg[13][20] ), .S(fanout_net_31 ), .Z(_04490_ ) );
MUX2_X1 _12214_ ( .A(_04489_ ), .B(_04490_ ), .S(_04317_ ), .Z(_04491_ ) );
OAI211_X1 _12215_ ( .A(fanout_net_41 ), .B(_04488_ ), .C1(_04491_ ), .C2(_04338_ ), .ZN(_04492_ ) );
NOR2_X1 _12216_ ( .A1(_04323_ ), .A2(\myreg.Reg[3][20] ), .ZN(_04493_ ) );
OAI21_X1 _12217_ ( .A(fanout_net_38 ), .B1(fanout_net_31 ), .B2(\myreg.Reg[2][20] ), .ZN(_04494_ ) );
NOR2_X1 _12218_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][20] ), .ZN(_04495_ ) );
OAI21_X1 _12219_ ( .A(_04331_ ), .B1(_04323_ ), .B2(\myreg.Reg[1][20] ), .ZN(_04496_ ) );
OAI221_X1 _12220_ ( .A(_04402_ ), .B1(_04493_ ), .B2(_04494_ ), .C1(_04495_ ), .C2(_04496_ ), .ZN(_04497_ ) );
MUX2_X1 _12221_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_31 ), .Z(_04498_ ) );
MUX2_X1 _12222_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_31 ), .Z(_04499_ ) );
MUX2_X1 _12223_ ( .A(_04498_ ), .B(_04499_ ), .S(_04317_ ), .Z(_04500_ ) );
OAI211_X1 _12224_ ( .A(_04310_ ), .B(_04497_ ), .C1(_04500_ ), .C2(_04338_ ), .ZN(_04501_ ) );
OAI211_X2 _12225_ ( .A(_04492_ ), .B(_04501_ ), .C1(_04303_ ), .C2(_04306_ ), .ZN(_04502_ ) );
NAND2_X1 _12226_ ( .A1(_04483_ ), .A2(_04502_ ), .ZN(_04503_ ) );
XOR2_X1 _12227_ ( .A(_02610_ ), .B(_04503_ ), .Z(_04504_ ) );
AND2_X4 _12228_ ( .A1(_02565_ ), .A2(_02585_ ), .ZN(_04505_ ) );
OR3_X2 _12229_ ( .A1(_04302_ ), .A2(\EX_LS_result_reg [21] ), .A3(_04305_ ), .ZN(_04506_ ) );
OR2_X1 _12230_ ( .A1(\myreg.Reg[0][21] ), .A2(fanout_net_31 ), .ZN(_04507_ ) );
OAI211_X1 _12231_ ( .A(_04507_ ), .B(_04316_ ), .C1(\myreg.Reg[1][21] ), .C2(_04393_ ), .ZN(_04508_ ) );
OR2_X1 _12232_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][21] ), .ZN(_04509_ ) );
OAI211_X1 _12233_ ( .A(_04509_ ), .B(fanout_net_38 ), .C1(_04393_ ), .C2(\myreg.Reg[3][21] ), .ZN(_04510_ ) );
NAND3_X1 _12234_ ( .A1(_04508_ ), .A2(_04510_ ), .A3(_04337_ ), .ZN(_04511_ ) );
MUX2_X1 _12235_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_31 ), .Z(_04512_ ) );
MUX2_X1 _12236_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_32 ), .Z(_04513_ ) );
MUX2_X1 _12237_ ( .A(_04512_ ), .B(_04513_ ), .S(_04316_ ), .Z(_04514_ ) );
OAI211_X1 _12238_ ( .A(_04310_ ), .B(_04511_ ), .C1(_04514_ ), .C2(_04402_ ), .ZN(_04515_ ) );
OR2_X1 _12239_ ( .A1(_04392_ ), .A2(\myreg.Reg[15][21] ), .ZN(_04516_ ) );
OAI211_X1 _12240_ ( .A(_04516_ ), .B(fanout_net_38 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[14][21] ), .ZN(_04517_ ) );
OR2_X1 _12241_ ( .A1(_04392_ ), .A2(\myreg.Reg[13][21] ), .ZN(_04518_ ) );
OAI211_X1 _12242_ ( .A(_04518_ ), .B(_04316_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[12][21] ), .ZN(_04519_ ) );
NAND3_X1 _12243_ ( .A1(_04517_ ), .A2(_04519_ ), .A3(fanout_net_40 ), .ZN(_04520_ ) );
MUX2_X1 _12244_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_32 ), .Z(_04521_ ) );
MUX2_X1 _12245_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_32 ), .Z(_04522_ ) );
MUX2_X1 _12246_ ( .A(_04521_ ), .B(_04522_ ), .S(fanout_net_38 ), .Z(_04523_ ) );
OAI211_X1 _12247_ ( .A(fanout_net_41 ), .B(_04520_ ), .C1(_04523_ ), .C2(fanout_net_40 ), .ZN(_04524_ ) );
OAI211_X2 _12248_ ( .A(_04515_ ), .B(_04524_ ), .C1(_04404_ ), .C2(_04354_ ), .ZN(_04525_ ) );
NAND2_X1 _12249_ ( .A1(_04506_ ), .A2(_04525_ ), .ZN(_04526_ ) );
AND2_X1 _12250_ ( .A1(_04505_ ), .A2(_04526_ ), .ZN(_04527_ ) );
NOR2_X1 _12251_ ( .A1(_04505_ ), .A2(_04526_ ), .ZN(_04528_ ) );
NOR2_X1 _12252_ ( .A1(_04527_ ), .A2(_04528_ ), .ZN(_04529_ ) );
NAND3_X1 _12253_ ( .A1(_04482_ ), .A2(_04504_ ), .A3(_04529_ ), .ZN(_04530_ ) );
NOR2_X1 _12254_ ( .A1(_04433_ ), .A2(_04530_ ), .ZN(_04531_ ) );
NOR2_X1 _12255_ ( .A1(_04300_ ), .A2(_02379_ ), .ZN(_04532_ ) );
NAND2_X1 _12256_ ( .A1(_04532_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_04533_ ) );
NOR2_X1 _12257_ ( .A1(_04324_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04534_ ) );
OAI21_X1 _12258_ ( .A(fanout_net_38 ), .B1(fanout_net_32 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04535_ ) );
NOR2_X1 _12259_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04536_ ) );
BUF_X4 _12260_ ( .A(_04340_ ), .Z(_04537_ ) );
OAI21_X1 _12261_ ( .A(_04318_ ), .B1(_04537_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04538_ ) );
OAI221_X1 _12262_ ( .A(_04349_ ), .B1(_04534_ ), .B2(_04535_ ), .C1(_04536_ ), .C2(_04538_ ), .ZN(_04539_ ) );
MUX2_X1 _12263_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04540_ ) );
MUX2_X1 _12264_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04541_ ) );
MUX2_X1 _12265_ ( .A(_04540_ ), .B(_04541_ ), .S(fanout_net_38 ), .Z(_04542_ ) );
BUF_X4 _12266_ ( .A(_04338_ ), .Z(_04543_ ) );
OAI211_X1 _12267_ ( .A(fanout_net_41 ), .B(_04539_ ), .C1(_04542_ ), .C2(_04543_ ), .ZN(_04544_ ) );
OR2_X1 _12268_ ( .A1(_04340_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04545_ ) );
BUF_X4 _12269_ ( .A(_04332_ ), .Z(_04546_ ) );
OAI211_X1 _12270_ ( .A(_04545_ ), .B(_04546_ ), .C1(fanout_net_32 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04547_ ) );
OR2_X1 _12271_ ( .A1(_04340_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04548_ ) );
OAI211_X1 _12272_ ( .A(_04548_ ), .B(fanout_net_38 ), .C1(fanout_net_32 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04549_ ) );
NAND3_X1 _12273_ ( .A1(_04547_ ), .A2(_04549_ ), .A3(fanout_net_40 ), .ZN(_04550_ ) );
MUX2_X1 _12274_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04551_ ) );
MUX2_X1 _12275_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04552_ ) );
MUX2_X1 _12276_ ( .A(_04551_ ), .B(_04552_ ), .S(_04318_ ), .Z(_04553_ ) );
OAI211_X1 _12277_ ( .A(_04311_ ), .B(_04550_ ), .C1(_04553_ ), .C2(fanout_net_40 ), .ZN(_04554_ ) );
NAND2_X1 _12278_ ( .A1(_04544_ ), .A2(_04554_ ), .ZN(_04555_ ) );
BUF_X2 _12279_ ( .A(_04306_ ), .Z(_04556_ ) );
BUF_X2 _12280_ ( .A(_04303_ ), .Z(_04557_ ) );
OAI21_X1 _12281_ ( .A(_04555_ ), .B1(_04556_ ), .B2(_04557_ ), .ZN(_04558_ ) );
AND2_X1 _12282_ ( .A1(_04533_ ), .A2(_04558_ ), .ZN(_04559_ ) );
XNOR2_X1 _12283_ ( .A(_02448_ ), .B(_04559_ ), .ZN(_04560_ ) );
OR3_X1 _12284_ ( .A1(_04303_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04306_ ), .ZN(_04561_ ) );
OR2_X1 _12285_ ( .A1(_04340_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04562_ ) );
OAI211_X1 _12286_ ( .A(_04562_ ), .B(fanout_net_38 ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04563_ ) );
OR2_X1 _12287_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04564_ ) );
OAI211_X1 _12288_ ( .A(_04564_ ), .B(_04318_ ), .C1(_04537_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04565_ ) );
NAND3_X1 _12289_ ( .A1(_04563_ ), .A2(_04543_ ), .A3(_04565_ ), .ZN(_04566_ ) );
MUX2_X1 _12290_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04567_ ) );
MUX2_X1 _12291_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04568_ ) );
MUX2_X1 _12292_ ( .A(_04567_ ), .B(_04568_ ), .S(_04318_ ), .Z(_04569_ ) );
OAI211_X1 _12293_ ( .A(_04311_ ), .B(_04566_ ), .C1(_04569_ ), .C2(_04543_ ), .ZN(_04570_ ) );
OR2_X1 _12294_ ( .A1(_04340_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04571_ ) );
OAI211_X1 _12295_ ( .A(_04571_ ), .B(_04546_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04572_ ) );
OR2_X1 _12296_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04573_ ) );
OAI211_X1 _12297_ ( .A(_04573_ ), .B(fanout_net_38 ), .C1(_04537_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04574_ ) );
NAND3_X1 _12298_ ( .A1(_04572_ ), .A2(fanout_net_40 ), .A3(_04574_ ), .ZN(_04575_ ) );
MUX2_X1 _12299_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04576_ ) );
MUX2_X1 _12300_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04577_ ) );
MUX2_X1 _12301_ ( .A(_04576_ ), .B(_04577_ ), .S(fanout_net_38 ), .Z(_04578_ ) );
OAI211_X1 _12302_ ( .A(fanout_net_41 ), .B(_04575_ ), .C1(_04578_ ), .C2(fanout_net_40 ), .ZN(_04579_ ) );
OAI211_X1 _12303_ ( .A(_04570_ ), .B(_04579_ ), .C1(_04557_ ), .C2(_04556_ ), .ZN(_04580_ ) );
NAND2_X1 _12304_ ( .A1(_04561_ ), .A2(_04580_ ), .ZN(_04581_ ) );
AND3_X1 _12305_ ( .A1(_02423_ ), .A2(_02424_ ), .A3(_04581_ ), .ZN(_04582_ ) );
AOI21_X1 _12306_ ( .A(_04581_ ), .B1(_02423_ ), .B2(_02424_ ), .ZN(_04583_ ) );
NOR2_X1 _12307_ ( .A1(_04582_ ), .A2(_04583_ ), .ZN(_04584_ ) );
AND2_X1 _12308_ ( .A1(_04560_ ), .A2(_04584_ ), .ZN(_04585_ ) );
OR3_X1 _12309_ ( .A1(_04557_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_04556_ ), .ZN(_04586_ ) );
OR2_X1 _12310_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04587_ ) );
OAI211_X1 _12311_ ( .A(_04587_ ), .B(_04546_ ), .C1(_04537_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04588_ ) );
OR2_X1 _12312_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04589_ ) );
OAI211_X1 _12313_ ( .A(_04589_ ), .B(fanout_net_39 ), .C1(_04537_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04590_ ) );
NAND3_X1 _12314_ ( .A1(_04588_ ), .A2(_04590_ ), .A3(fanout_net_40 ), .ZN(_04591_ ) );
MUX2_X1 _12315_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04592_ ) );
MUX2_X1 _12316_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04593_ ) );
MUX2_X1 _12317_ ( .A(_04592_ ), .B(_04593_ ), .S(_04546_ ), .Z(_04594_ ) );
OAI211_X1 _12318_ ( .A(_04311_ ), .B(_04591_ ), .C1(_04594_ ), .C2(fanout_net_40 ), .ZN(_04595_ ) );
NOR2_X1 _12319_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04596_ ) );
OAI21_X1 _12320_ ( .A(_04546_ ), .B1(_04537_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04597_ ) );
MUX2_X1 _12321_ ( .A(_02358_ ), .B(_02359_ ), .S(fanout_net_32 ), .Z(_04598_ ) );
OAI221_X1 _12322_ ( .A(_04543_ ), .B1(_04596_ ), .B2(_04597_ ), .C1(_04598_ ), .C2(_04546_ ), .ZN(_04599_ ) );
MUX2_X1 _12323_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04600_ ) );
MUX2_X1 _12324_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04601_ ) );
MUX2_X1 _12325_ ( .A(_04600_ ), .B(_04601_ ), .S(fanout_net_39 ), .Z(_04602_ ) );
OAI211_X1 _12326_ ( .A(fanout_net_41 ), .B(_04599_ ), .C1(_04602_ ), .C2(_04543_ ), .ZN(_04603_ ) );
OAI211_X1 _12327_ ( .A(_04595_ ), .B(_04603_ ), .C1(_04557_ ), .C2(_04556_ ), .ZN(_04604_ ) );
NAND2_X1 _12328_ ( .A1(_04586_ ), .A2(_04604_ ), .ZN(_04605_ ) );
INV_X1 _12329_ ( .A(_04605_ ), .ZN(_04606_ ) );
XNOR2_X1 _12330_ ( .A(_02401_ ), .B(_04606_ ), .ZN(_04607_ ) );
NAND2_X1 _12331_ ( .A1(_04532_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04608_ ) );
OR2_X1 _12332_ ( .A1(_04323_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04609_ ) );
OAI211_X1 _12333_ ( .A(_04609_ ), .B(_04332_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04610_ ) );
OR2_X1 _12334_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04611_ ) );
OAI211_X1 _12335_ ( .A(_04611_ ), .B(fanout_net_39 ), .C1(_04324_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04612_ ) );
NAND3_X1 _12336_ ( .A1(_04610_ ), .A2(_04349_ ), .A3(_04612_ ), .ZN(_04613_ ) );
MUX2_X1 _12337_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04614_ ) );
MUX2_X1 _12338_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04615_ ) );
MUX2_X1 _12339_ ( .A(_04614_ ), .B(_04615_ ), .S(_04332_ ), .Z(_04616_ ) );
OAI211_X1 _12340_ ( .A(_04311_ ), .B(_04613_ ), .C1(_04616_ ), .C2(_04349_ ), .ZN(_04617_ ) );
OR2_X1 _12341_ ( .A1(_04323_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04618_ ) );
OAI211_X1 _12342_ ( .A(_04618_ ), .B(fanout_net_39 ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04619_ ) );
OR2_X1 _12343_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04620_ ) );
OAI211_X1 _12344_ ( .A(_04620_ ), .B(_04332_ ), .C1(_04324_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04621_ ) );
NAND3_X1 _12345_ ( .A1(_04619_ ), .A2(fanout_net_40 ), .A3(_04621_ ), .ZN(_04622_ ) );
MUX2_X1 _12346_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04623_ ) );
MUX2_X1 _12347_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04624_ ) );
MUX2_X1 _12348_ ( .A(_04623_ ), .B(_04624_ ), .S(fanout_net_39 ), .Z(_04625_ ) );
OAI211_X1 _12349_ ( .A(fanout_net_41 ), .B(_04622_ ), .C1(_04625_ ), .C2(fanout_net_40 ), .ZN(_04626_ ) );
NAND2_X1 _12350_ ( .A1(_04617_ ), .A2(_04626_ ), .ZN(_04627_ ) );
OAI21_X1 _12351_ ( .A(_04627_ ), .B1(_04556_ ), .B2(_04557_ ), .ZN(_04628_ ) );
AND2_X1 _12352_ ( .A1(_04608_ ), .A2(_04628_ ), .ZN(_04629_ ) );
XNOR2_X1 _12353_ ( .A(_03243_ ), .B(_04629_ ), .ZN(_04630_ ) );
AND3_X1 _12354_ ( .A1(_04585_ ), .A2(_04607_ ), .A3(_04630_ ), .ZN(_04631_ ) );
OR3_X1 _12355_ ( .A1(_04303_ ), .A2(\EX_LS_result_reg [24] ), .A3(_04306_ ), .ZN(_04632_ ) );
NOR2_X1 _12356_ ( .A1(_04340_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04633_ ) );
OAI21_X1 _12357_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04634_ ) );
NOR2_X1 _12358_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04635_ ) );
OAI21_X1 _12359_ ( .A(_04332_ ), .B1(_04324_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04636_ ) );
OAI221_X1 _12360_ ( .A(_04349_ ), .B1(_04633_ ), .B2(_04634_ ), .C1(_04635_ ), .C2(_04636_ ), .ZN(_04637_ ) );
MUX2_X1 _12361_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04638_ ) );
MUX2_X1 _12362_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04639_ ) );
MUX2_X1 _12363_ ( .A(_04638_ ), .B(_04639_ ), .S(fanout_net_39 ), .Z(_04640_ ) );
OAI211_X1 _12364_ ( .A(fanout_net_41 ), .B(_04637_ ), .C1(_04640_ ), .C2(_04349_ ), .ZN(_04641_ ) );
OR2_X1 _12365_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04642_ ) );
OAI211_X1 _12366_ ( .A(_04642_ ), .B(_04318_ ), .C1(_04324_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04643_ ) );
OR2_X1 _12367_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04644_ ) );
OAI211_X1 _12368_ ( .A(_04644_ ), .B(fanout_net_39 ), .C1(_04324_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04645_ ) );
NAND3_X1 _12369_ ( .A1(_04643_ ), .A2(_04645_ ), .A3(fanout_net_40 ), .ZN(_04646_ ) );
MUX2_X1 _12370_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04647_ ) );
MUX2_X1 _12371_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04648_ ) );
MUX2_X1 _12372_ ( .A(_04647_ ), .B(_04648_ ), .S(_04332_ ), .Z(_04649_ ) );
OAI211_X1 _12373_ ( .A(_04311_ ), .B(_04646_ ), .C1(_04649_ ), .C2(fanout_net_40 ), .ZN(_04650_ ) );
NAND2_X1 _12374_ ( .A1(_04641_ ), .A2(_04650_ ), .ZN(_04651_ ) );
OAI21_X1 _12375_ ( .A(_04651_ ), .B1(_04556_ ), .B2(_04557_ ), .ZN(_04652_ ) );
AND2_X1 _12376_ ( .A1(_04632_ ), .A2(_04652_ ), .ZN(_04653_ ) );
XNOR2_X1 _12377_ ( .A(_02510_ ), .B(_04653_ ), .ZN(_04654_ ) );
INV_X1 _12378_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04655_ ) );
OR3_X1 _12379_ ( .A1(_04557_ ), .A2(_04655_ ), .A3(_04306_ ), .ZN(_04656_ ) );
OR2_X1 _12380_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04657_ ) );
OAI211_X1 _12381_ ( .A(_04657_ ), .B(fanout_net_39 ), .C1(_04537_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04658_ ) );
NAND2_X1 _12382_ ( .A1(_03166_ ), .A2(fanout_net_33 ), .ZN(_04659_ ) );
OAI211_X1 _12383_ ( .A(_04659_ ), .B(_04318_ ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04660_ ) );
NAND3_X1 _12384_ ( .A1(_04658_ ), .A2(_04660_ ), .A3(_04543_ ), .ZN(_04661_ ) );
MUX2_X1 _12385_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04662_ ) );
MUX2_X1 _12386_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04663_ ) );
MUX2_X1 _12387_ ( .A(_04662_ ), .B(_04663_ ), .S(_04318_ ), .Z(_04664_ ) );
OAI211_X1 _12388_ ( .A(fanout_net_41 ), .B(_04661_ ), .C1(_04664_ ), .C2(_04543_ ), .ZN(_04665_ ) );
OR2_X1 _12389_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04666_ ) );
OAI211_X1 _12390_ ( .A(_04666_ ), .B(_04318_ ), .C1(_04537_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04667_ ) );
NOR2_X1 _12391_ ( .A1(_04537_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04668_ ) );
OAI21_X1 _12392_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04669_ ) );
OAI211_X1 _12393_ ( .A(_04667_ ), .B(_04349_ ), .C1(_04668_ ), .C2(_04669_ ), .ZN(_04670_ ) );
MUX2_X1 _12394_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04671_ ) );
MUX2_X1 _12395_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04672_ ) );
MUX2_X1 _12396_ ( .A(_04671_ ), .B(_04672_ ), .S(_04318_ ), .Z(_04673_ ) );
OAI211_X1 _12397_ ( .A(_04311_ ), .B(_04670_ ), .C1(_04673_ ), .C2(_04543_ ), .ZN(_04674_ ) );
OAI211_X1 _12398_ ( .A(_04665_ ), .B(_04674_ ), .C1(_04557_ ), .C2(_04556_ ), .ZN(_04675_ ) );
NAND2_X1 _12399_ ( .A1(_04656_ ), .A2(_04675_ ), .ZN(_04676_ ) );
XNOR2_X1 _12400_ ( .A(_03184_ ), .B(_04676_ ), .ZN(_04677_ ) );
AND2_X1 _12401_ ( .A1(_04654_ ), .A2(_04677_ ), .ZN(_04678_ ) );
OR3_X1 _12402_ ( .A1(_04303_ ), .A2(\EX_LS_result_reg [26] ), .A3(_04306_ ), .ZN(_04679_ ) );
NOR2_X1 _12403_ ( .A1(_04323_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04680_ ) );
OAI21_X1 _12404_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04681_ ) );
NOR2_X1 _12405_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04682_ ) );
OAI21_X1 _12406_ ( .A(_04317_ ), .B1(_04340_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04683_ ) );
OAI221_X1 _12407_ ( .A(_04338_ ), .B1(_04680_ ), .B2(_04681_ ), .C1(_04682_ ), .C2(_04683_ ), .ZN(_04684_ ) );
MUX2_X1 _12408_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04685_ ) );
MUX2_X1 _12409_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04686_ ) );
MUX2_X1 _12410_ ( .A(_04685_ ), .B(_04686_ ), .S(_04332_ ), .Z(_04687_ ) );
OAI211_X1 _12411_ ( .A(_04311_ ), .B(_04684_ ), .C1(_04687_ ), .C2(_04349_ ), .ZN(_04688_ ) );
OR2_X1 _12412_ ( .A1(_04323_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04689_ ) );
OAI211_X1 _12413_ ( .A(_04689_ ), .B(fanout_net_39 ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04690_ ) );
OR2_X1 _12414_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04691_ ) );
OAI211_X1 _12415_ ( .A(_04691_ ), .B(_04332_ ), .C1(_04340_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04692_ ) );
NAND3_X1 _12416_ ( .A1(_04690_ ), .A2(_04338_ ), .A3(_04692_ ), .ZN(_04693_ ) );
MUX2_X1 _12417_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04694_ ) );
MUX2_X1 _12418_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04695_ ) );
MUX2_X1 _12419_ ( .A(_04694_ ), .B(_04695_ ), .S(_04317_ ), .Z(_04696_ ) );
OAI211_X1 _12420_ ( .A(fanout_net_41 ), .B(_04693_ ), .C1(_04696_ ), .C2(_04349_ ), .ZN(_04697_ ) );
NAND2_X1 _12421_ ( .A1(_04688_ ), .A2(_04697_ ), .ZN(_04698_ ) );
OAI21_X1 _12422_ ( .A(_04698_ ), .B1(_04556_ ), .B2(_04303_ ), .ZN(_04699_ ) );
AND2_X1 _12423_ ( .A1(_04679_ ), .A2(_04699_ ), .ZN(_04700_ ) );
XNOR2_X1 _12424_ ( .A(_03207_ ), .B(_04700_ ), .ZN(_04701_ ) );
INV_X1 _12425_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04702_ ) );
OR3_X1 _12426_ ( .A1(_04557_ ), .A2(_04702_ ), .A3(_04556_ ), .ZN(_04703_ ) );
OR2_X1 _12427_ ( .A1(_04324_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04704_ ) );
OAI211_X1 _12428_ ( .A(_04704_ ), .B(_04546_ ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04705_ ) );
OR2_X1 _12429_ ( .A1(_04324_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04706_ ) );
OAI211_X1 _12430_ ( .A(_04706_ ), .B(fanout_net_39 ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04707_ ) );
NAND3_X1 _12431_ ( .A1(_04705_ ), .A2(_04707_ ), .A3(fanout_net_40 ), .ZN(_04708_ ) );
MUX2_X1 _12432_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04709_ ) );
MUX2_X1 _12433_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04710_ ) );
MUX2_X1 _12434_ ( .A(_04709_ ), .B(_04710_ ), .S(_04546_ ), .Z(_04711_ ) );
OAI211_X1 _12435_ ( .A(_04311_ ), .B(_04708_ ), .C1(_04711_ ), .C2(fanout_net_40 ), .ZN(_04712_ ) );
NOR2_X1 _12436_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04713_ ) );
OAI21_X1 _12437_ ( .A(_04546_ ), .B1(_04537_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04714_ ) );
MUX2_X1 _12438_ ( .A(_02464_ ), .B(_02465_ ), .S(fanout_net_34 ), .Z(_04715_ ) );
OAI221_X1 _12439_ ( .A(_04543_ ), .B1(_04713_ ), .B2(_04714_ ), .C1(_04715_ ), .C2(_04546_ ), .ZN(_04716_ ) );
MUX2_X1 _12440_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04717_ ) );
MUX2_X1 _12441_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04718_ ) );
MUX2_X1 _12442_ ( .A(_04717_ ), .B(_04718_ ), .S(fanout_net_39 ), .Z(_04719_ ) );
OAI211_X1 _12443_ ( .A(fanout_net_41 ), .B(_04716_ ), .C1(_04719_ ), .C2(_04543_ ), .ZN(_04720_ ) );
OAI211_X1 _12444_ ( .A(_04712_ ), .B(_04720_ ), .C1(_04557_ ), .C2(_04556_ ), .ZN(_04721_ ) );
NAND2_X1 _12445_ ( .A1(_04703_ ), .A2(_04721_ ), .ZN(_04722_ ) );
XNOR2_X1 _12446_ ( .A(_02487_ ), .B(_04722_ ), .ZN(_04723_ ) );
AND2_X1 _12447_ ( .A1(_04701_ ), .A2(_04723_ ), .ZN(_04724_ ) );
AND2_X1 _12448_ ( .A1(_04678_ ), .A2(_04724_ ), .ZN(_04725_ ) );
AND2_X1 _12449_ ( .A1(_04631_ ), .A2(_04725_ ), .ZN(_04726_ ) );
AND2_X1 _12450_ ( .A1(_04531_ ), .A2(_04726_ ), .ZN(_04727_ ) );
OR3_X1 _12451_ ( .A1(_04300_ ), .A2(\EX_LS_result_reg [14] ), .A3(_02379_ ), .ZN(_04728_ ) );
OR2_X1 _12452_ ( .A1(_04391_ ), .A2(\myreg.Reg[9][14] ), .ZN(_04729_ ) );
BUF_X4 _12453_ ( .A(_04313_ ), .Z(_04730_ ) );
OAI211_X1 _12454_ ( .A(_04729_ ), .B(_04730_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[8][14] ), .ZN(_04731_ ) );
OR2_X1 _12455_ ( .A1(_04320_ ), .A2(\myreg.Reg[11][14] ), .ZN(_04732_ ) );
OAI211_X1 _12456_ ( .A(_04732_ ), .B(fanout_net_39 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[10][14] ), .ZN(_04733_ ) );
NAND3_X1 _12457_ ( .A1(_04731_ ), .A2(_04733_ ), .A3(_04336_ ), .ZN(_04734_ ) );
MUX2_X1 _12458_ ( .A(\myreg.Reg[14][14] ), .B(\myreg.Reg[15][14] ), .S(fanout_net_34 ), .Z(_04735_ ) );
MUX2_X1 _12459_ ( .A(\myreg.Reg[12][14] ), .B(\myreg.Reg[13][14] ), .S(fanout_net_34 ), .Z(_04736_ ) );
MUX2_X1 _12460_ ( .A(_04735_ ), .B(_04736_ ), .S(_04314_ ), .Z(_04737_ ) );
BUF_X4 _12461_ ( .A(_04335_ ), .Z(_04738_ ) );
OAI211_X1 _12462_ ( .A(fanout_net_41 ), .B(_04734_ ), .C1(_04737_ ), .C2(_04738_ ), .ZN(_04739_ ) );
OR2_X1 _12463_ ( .A1(_04391_ ), .A2(\myreg.Reg[1][14] ), .ZN(_04740_ ) );
OAI211_X1 _12464_ ( .A(_04740_ ), .B(_04730_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[0][14] ), .ZN(_04741_ ) );
OR2_X1 _12465_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[2][14] ), .ZN(_04742_ ) );
OAI211_X1 _12466_ ( .A(_04742_ ), .B(fanout_net_39 ), .C1(_04321_ ), .C2(\myreg.Reg[3][14] ), .ZN(_04743_ ) );
NAND3_X1 _12467_ ( .A1(_04741_ ), .A2(_04336_ ), .A3(_04743_ ), .ZN(_04744_ ) );
MUX2_X1 _12468_ ( .A(\myreg.Reg[6][14] ), .B(\myreg.Reg[7][14] ), .S(fanout_net_34 ), .Z(_04745_ ) );
MUX2_X1 _12469_ ( .A(\myreg.Reg[4][14] ), .B(\myreg.Reg[5][14] ), .S(fanout_net_34 ), .Z(_04746_ ) );
MUX2_X1 _12470_ ( .A(_04745_ ), .B(_04746_ ), .S(_04314_ ), .Z(_04747_ ) );
BUF_X4 _12471_ ( .A(_04335_ ), .Z(_04748_ ) );
OAI211_X1 _12472_ ( .A(_04309_ ), .B(_04744_ ), .C1(_04747_ ), .C2(_04748_ ), .ZN(_04749_ ) );
BUF_X4 _12473_ ( .A(_02379_ ), .Z(_04750_ ) );
OAI211_X2 _12474_ ( .A(_04739_ ), .B(_04749_ ), .C1(_04301_ ), .C2(_04750_ ), .ZN(_04751_ ) );
NAND2_X2 _12475_ ( .A1(_04728_ ), .A2(_04751_ ), .ZN(_04752_ ) );
XOR2_X1 _12476_ ( .A(_03020_ ), .B(_04752_ ), .Z(_04753_ ) );
OR3_X4 _12477_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [15] ), .A3(_04304_ ), .ZN(_04754_ ) );
OR2_X1 _12478_ ( .A1(_04391_ ), .A2(\myreg.Reg[11][15] ), .ZN(_04755_ ) );
OAI211_X1 _12479_ ( .A(_04755_ ), .B(fanout_net_39 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[10][15] ), .ZN(_04756_ ) );
OR2_X1 _12480_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[8][15] ), .ZN(_04757_ ) );
BUF_X4 _12481_ ( .A(_04313_ ), .Z(_04758_ ) );
BUF_X4 _12482_ ( .A(_04391_ ), .Z(_04759_ ) );
OAI211_X1 _12483_ ( .A(_04757_ ), .B(_04758_ ), .C1(_04759_ ), .C2(\myreg.Reg[9][15] ), .ZN(_04760_ ) );
NAND3_X1 _12484_ ( .A1(_04756_ ), .A2(_04748_ ), .A3(_04760_ ), .ZN(_04761_ ) );
MUX2_X1 _12485_ ( .A(\myreg.Reg[14][15] ), .B(\myreg.Reg[15][15] ), .S(fanout_net_34 ), .Z(_04762_ ) );
MUX2_X1 _12486_ ( .A(\myreg.Reg[12][15] ), .B(\myreg.Reg[13][15] ), .S(fanout_net_34 ), .Z(_04763_ ) );
MUX2_X1 _12487_ ( .A(_04762_ ), .B(_04763_ ), .S(_04730_ ), .Z(_04764_ ) );
OAI211_X1 _12488_ ( .A(fanout_net_41 ), .B(_04761_ ), .C1(_04764_ ), .C2(_04738_ ), .ZN(_04765_ ) );
OR2_X1 _12489_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[0][15] ), .ZN(_04766_ ) );
OAI211_X1 _12490_ ( .A(_04766_ ), .B(_04730_ ), .C1(_04759_ ), .C2(\myreg.Reg[1][15] ), .ZN(_04767_ ) );
NOR2_X1 _12491_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[2][15] ), .ZN(_04768_ ) );
OAI21_X1 _12492_ ( .A(fanout_net_39 ), .B1(_04759_ ), .B2(\myreg.Reg[3][15] ), .ZN(_04769_ ) );
OAI211_X1 _12493_ ( .A(_04767_ ), .B(_04336_ ), .C1(_04768_ ), .C2(_04769_ ), .ZN(_04770_ ) );
MUX2_X1 _12494_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_34 ), .Z(_04771_ ) );
MUX2_X1 _12495_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_34 ), .Z(_04772_ ) );
MUX2_X1 _12496_ ( .A(_04771_ ), .B(_04772_ ), .S(_04730_ ), .Z(_04773_ ) );
OAI211_X1 _12497_ ( .A(_04309_ ), .B(_04770_ ), .C1(_04773_ ), .C2(_04738_ ), .ZN(_04774_ ) );
BUF_X4 _12498_ ( .A(_04300_ ), .Z(_04775_ ) );
OAI211_X1 _12499_ ( .A(_04765_ ), .B(_04774_ ), .C1(_04775_ ), .C2(_04750_ ), .ZN(_04776_ ) );
NAND2_X1 _12500_ ( .A1(_04754_ ), .A2(_04776_ ), .ZN(_04777_ ) );
INV_X1 _12501_ ( .A(_04777_ ), .ZN(_04778_ ) );
XNOR2_X1 _12502_ ( .A(_02996_ ), .B(_04778_ ), .ZN(_04779_ ) );
AND2_X1 _12503_ ( .A1(_04753_ ), .A2(_04779_ ), .ZN(_04780_ ) );
AND2_X4 _12504_ ( .A1(_02950_ ), .A2(_02970_ ), .ZN(_04781_ ) );
OR3_X1 _12505_ ( .A1(_04300_ ), .A2(\EX_LS_result_reg [13] ), .A3(_02379_ ), .ZN(_04782_ ) );
OR2_X1 _12506_ ( .A1(_04320_ ), .A2(\myreg.Reg[11][13] ), .ZN(_04783_ ) );
OAI211_X1 _12507_ ( .A(_04783_ ), .B(fanout_net_39 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[10][13] ), .ZN(_04784_ ) );
OR2_X1 _12508_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[8][13] ), .ZN(_04785_ ) );
BUF_X4 _12509_ ( .A(_04320_ ), .Z(_04786_ ) );
OAI211_X1 _12510_ ( .A(_04785_ ), .B(_04314_ ), .C1(_04786_ ), .C2(\myreg.Reg[9][13] ), .ZN(_04787_ ) );
NAND3_X1 _12511_ ( .A1(_04784_ ), .A2(_04336_ ), .A3(_04787_ ), .ZN(_04788_ ) );
MUX2_X1 _12512_ ( .A(\myreg.Reg[14][13] ), .B(\myreg.Reg[15][13] ), .S(fanout_net_34 ), .Z(_04789_ ) );
MUX2_X1 _12513_ ( .A(\myreg.Reg[12][13] ), .B(\myreg.Reg[13][13] ), .S(fanout_net_34 ), .Z(_04790_ ) );
BUF_X4 _12514_ ( .A(_04313_ ), .Z(_04791_ ) );
MUX2_X1 _12515_ ( .A(_04789_ ), .B(_04790_ ), .S(_04791_ ), .Z(_04792_ ) );
OAI211_X1 _12516_ ( .A(fanout_net_41 ), .B(_04788_ ), .C1(_04792_ ), .C2(_04748_ ), .ZN(_04793_ ) );
OR2_X1 _12517_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][13] ), .ZN(_04794_ ) );
OAI211_X1 _12518_ ( .A(_04794_ ), .B(_04791_ ), .C1(_04391_ ), .C2(\myreg.Reg[1][13] ), .ZN(_04795_ ) );
NOR2_X1 _12519_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][13] ), .ZN(_04796_ ) );
OAI21_X1 _12520_ ( .A(fanout_net_39 ), .B1(_04786_ ), .B2(\myreg.Reg[3][13] ), .ZN(_04797_ ) );
OAI211_X1 _12521_ ( .A(_04795_ ), .B(_04335_ ), .C1(_04796_ ), .C2(_04797_ ), .ZN(_04798_ ) );
MUX2_X1 _12522_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_35 ), .Z(_04799_ ) );
MUX2_X1 _12523_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_35 ), .Z(_04800_ ) );
MUX2_X1 _12524_ ( .A(_04799_ ), .B(_04800_ ), .S(_04791_ ), .Z(_04801_ ) );
OAI211_X1 _12525_ ( .A(_04308_ ), .B(_04798_ ), .C1(_04801_ ), .C2(_04748_ ), .ZN(_04802_ ) );
OAI211_X2 _12526_ ( .A(_04793_ ), .B(_04802_ ), .C1(_04301_ ), .C2(_04304_ ), .ZN(_04803_ ) );
NAND2_X1 _12527_ ( .A1(_04782_ ), .A2(_04803_ ), .ZN(_04804_ ) );
INV_X1 _12528_ ( .A(_04804_ ), .ZN(_04805_ ) );
XNOR2_X1 _12529_ ( .A(_04781_ ), .B(_04805_ ), .ZN(_04806_ ) );
OR3_X2 _12530_ ( .A1(_04775_ ), .A2(\EX_LS_result_reg [12] ), .A3(_04750_ ), .ZN(_04807_ ) );
OR2_X1 _12531_ ( .A1(_04786_ ), .A2(\myreg.Reg[9][12] ), .ZN(_04808_ ) );
OAI211_X1 _12532_ ( .A(_04808_ ), .B(_04758_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[8][12] ), .ZN(_04809_ ) );
OR2_X1 _12533_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[10][12] ), .ZN(_04810_ ) );
OAI211_X1 _12534_ ( .A(_04810_ ), .B(fanout_net_39 ), .C1(_04392_ ), .C2(\myreg.Reg[11][12] ), .ZN(_04811_ ) );
NAND3_X1 _12535_ ( .A1(_04809_ ), .A2(_04738_ ), .A3(_04811_ ), .ZN(_04812_ ) );
MUX2_X1 _12536_ ( .A(\myreg.Reg[14][12] ), .B(\myreg.Reg[15][12] ), .S(fanout_net_35 ), .Z(_04813_ ) );
MUX2_X1 _12537_ ( .A(\myreg.Reg[12][12] ), .B(\myreg.Reg[13][12] ), .S(fanout_net_35 ), .Z(_04814_ ) );
MUX2_X1 _12538_ ( .A(_04813_ ), .B(_04814_ ), .S(_04758_ ), .Z(_04815_ ) );
OAI211_X1 _12539_ ( .A(fanout_net_41 ), .B(_04812_ ), .C1(_04815_ ), .C2(_04337_ ), .ZN(_04816_ ) );
NOR2_X1 _12540_ ( .A1(_04759_ ), .A2(\myreg.Reg[3][12] ), .ZN(_04817_ ) );
OAI21_X1 _12541_ ( .A(fanout_net_39 ), .B1(fanout_net_35 ), .B2(\myreg.Reg[2][12] ), .ZN(_04818_ ) );
NOR2_X1 _12542_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][12] ), .ZN(_04819_ ) );
OAI21_X1 _12543_ ( .A(_04758_ ), .B1(_04759_ ), .B2(\myreg.Reg[1][12] ), .ZN(_04820_ ) );
OAI221_X1 _12544_ ( .A(_04748_ ), .B1(_04817_ ), .B2(_04818_ ), .C1(_04819_ ), .C2(_04820_ ), .ZN(_04821_ ) );
MUX2_X1 _12545_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_35 ), .Z(_04822_ ) );
MUX2_X1 _12546_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_35 ), .Z(_04823_ ) );
MUX2_X1 _12547_ ( .A(_04822_ ), .B(_04823_ ), .S(_04758_ ), .Z(_04824_ ) );
OAI211_X1 _12548_ ( .A(_04309_ ), .B(_04821_ ), .C1(_04824_ ), .C2(_04337_ ), .ZN(_04825_ ) );
OAI211_X4 _12549_ ( .A(_04816_ ), .B(_04825_ ), .C1(_04302_ ), .C2(_04305_ ), .ZN(_04826_ ) );
NAND2_X1 _12550_ ( .A1(_04807_ ), .A2(_04826_ ), .ZN(_04827_ ) );
XOR2_X1 _12551_ ( .A(_02948_ ), .B(_04827_ ), .Z(_04828_ ) );
AND3_X1 _12552_ ( .A1(_04780_ ), .A2(_04806_ ), .A3(_04828_ ), .ZN(_04829_ ) );
INV_X1 _12553_ ( .A(\EX_LS_result_reg [11] ), .ZN(_04830_ ) );
OR3_X2 _12554_ ( .A1(_04300_ ), .A2(_04830_ ), .A3(_02379_ ), .ZN(_04831_ ) );
OR2_X1 _12555_ ( .A1(_04319_ ), .A2(\myreg.Reg[1][11] ), .ZN(_04832_ ) );
OAI211_X1 _12556_ ( .A(_04832_ ), .B(_04313_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[0][11] ), .ZN(_04833_ ) );
OR2_X1 _12557_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][11] ), .ZN(_04834_ ) );
OAI211_X1 _12558_ ( .A(_04834_ ), .B(fanout_net_39 ), .C1(_04319_ ), .C2(\myreg.Reg[3][11] ), .ZN(_04835_ ) );
NAND3_X1 _12559_ ( .A1(_04833_ ), .A2(_04335_ ), .A3(_04835_ ), .ZN(_04836_ ) );
MUX2_X1 _12560_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_35 ), .Z(_04837_ ) );
MUX2_X1 _12561_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_35 ), .Z(_04838_ ) );
MUX2_X1 _12562_ ( .A(_04837_ ), .B(_04838_ ), .S(_04313_ ), .Z(_04839_ ) );
OAI211_X1 _12563_ ( .A(_04308_ ), .B(_04836_ ), .C1(_04839_ ), .C2(_04335_ ), .ZN(_04840_ ) );
OR2_X1 _12564_ ( .A1(_04319_ ), .A2(\myreg.Reg[15][11] ), .ZN(_04841_ ) );
OAI211_X1 _12565_ ( .A(_04841_ ), .B(fanout_net_39 ), .C1(fanout_net_35 ), .C2(\myreg.Reg[14][11] ), .ZN(_04842_ ) );
OR2_X1 _12566_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[12][11] ), .ZN(_04843_ ) );
OAI211_X1 _12567_ ( .A(_04843_ ), .B(_04313_ ), .C1(_04319_ ), .C2(\myreg.Reg[13][11] ), .ZN(_04844_ ) );
NAND3_X1 _12568_ ( .A1(_04842_ ), .A2(fanout_net_40 ), .A3(_04844_ ), .ZN(_04845_ ) );
MUX2_X1 _12569_ ( .A(\myreg.Reg[8][11] ), .B(\myreg.Reg[9][11] ), .S(fanout_net_35 ), .Z(_04846_ ) );
MUX2_X1 _12570_ ( .A(\myreg.Reg[10][11] ), .B(\myreg.Reg[11][11] ), .S(fanout_net_35 ), .Z(_04847_ ) );
MUX2_X1 _12571_ ( .A(_04846_ ), .B(_04847_ ), .S(fanout_net_39 ), .Z(_04848_ ) );
OAI211_X1 _12572_ ( .A(fanout_net_41 ), .B(_04845_ ), .C1(_04848_ ), .C2(fanout_net_40 ), .ZN(_04849_ ) );
NAND2_X1 _12573_ ( .A1(_04840_ ), .A2(_04849_ ), .ZN(_04850_ ) );
OAI21_X1 _12574_ ( .A(_04850_ ), .B1(_02379_ ), .B2(_04300_ ), .ZN(_04851_ ) );
AND2_X2 _12575_ ( .A1(_04831_ ), .A2(_04851_ ), .ZN(_04852_ ) );
INV_X1 _12576_ ( .A(_04852_ ), .ZN(_04853_ ) );
AND2_X2 _12577_ ( .A1(_03098_ ), .A2(_03118_ ), .ZN(_04854_ ) );
XNOR2_X1 _12578_ ( .A(_04853_ ), .B(_04854_ ), .ZN(_04855_ ) );
OR3_X1 _12579_ ( .A1(_04775_ ), .A2(\EX_LS_result_reg [10] ), .A3(_04304_ ), .ZN(_04856_ ) );
OR2_X1 _12580_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][10] ), .ZN(_04857_ ) );
OAI211_X1 _12581_ ( .A(_04857_ ), .B(_04758_ ), .C1(_04759_ ), .C2(\myreg.Reg[1][10] ), .ZN(_04858_ ) );
OR2_X1 _12582_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][10] ), .ZN(_04859_ ) );
OAI211_X1 _12583_ ( .A(_04859_ ), .B(fanout_net_39 ), .C1(_04759_ ), .C2(\myreg.Reg[3][10] ), .ZN(_04860_ ) );
NAND3_X1 _12584_ ( .A1(_04858_ ), .A2(_04860_ ), .A3(_04748_ ), .ZN(_04861_ ) );
MUX2_X1 _12585_ ( .A(\myreg.Reg[6][10] ), .B(\myreg.Reg[7][10] ), .S(fanout_net_35 ), .Z(_04862_ ) );
MUX2_X1 _12586_ ( .A(\myreg.Reg[4][10] ), .B(\myreg.Reg[5][10] ), .S(fanout_net_35 ), .Z(_04863_ ) );
MUX2_X1 _12587_ ( .A(_04862_ ), .B(_04863_ ), .S(_04758_ ), .Z(_04864_ ) );
OAI211_X1 _12588_ ( .A(_04309_ ), .B(_04861_ ), .C1(_04864_ ), .C2(_04738_ ), .ZN(_04865_ ) );
OR2_X1 _12589_ ( .A1(_04391_ ), .A2(\myreg.Reg[15][10] ), .ZN(_04866_ ) );
OAI211_X1 _12590_ ( .A(_04866_ ), .B(fanout_net_39 ), .C1(fanout_net_35 ), .C2(\myreg.Reg[14][10] ), .ZN(_04867_ ) );
OR2_X1 _12591_ ( .A1(_04391_ ), .A2(\myreg.Reg[13][10] ), .ZN(_04868_ ) );
OAI211_X1 _12592_ ( .A(_04868_ ), .B(_04758_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[12][10] ), .ZN(_04869_ ) );
NAND3_X1 _12593_ ( .A1(_04867_ ), .A2(_04869_ ), .A3(fanout_net_40 ), .ZN(_04870_ ) );
MUX2_X1 _12594_ ( .A(\myreg.Reg[8][10] ), .B(\myreg.Reg[9][10] ), .S(fanout_net_35 ), .Z(_04871_ ) );
MUX2_X1 _12595_ ( .A(\myreg.Reg[10][10] ), .B(\myreg.Reg[11][10] ), .S(fanout_net_35 ), .Z(_04872_ ) );
MUX2_X1 _12596_ ( .A(_04871_ ), .B(_04872_ ), .S(fanout_net_39 ), .Z(_04873_ ) );
OAI211_X1 _12597_ ( .A(fanout_net_41 ), .B(_04870_ ), .C1(_04873_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04874_ ) );
OAI211_X1 _12598_ ( .A(_04865_ ), .B(_04874_ ), .C1(_04775_ ), .C2(_04750_ ), .ZN(_04875_ ) );
NAND2_X1 _12599_ ( .A1(_04856_ ), .A2(_04875_ ), .ZN(_04876_ ) );
INV_X1 _12600_ ( .A(_04876_ ), .ZN(_04877_ ) );
XNOR2_X1 _12601_ ( .A(_03095_ ), .B(_04877_ ), .ZN(_04878_ ) );
AND2_X1 _12602_ ( .A1(_04855_ ), .A2(_04878_ ), .ZN(_04879_ ) );
OR3_X1 _12603_ ( .A1(_04775_ ), .A2(\EX_LS_result_reg [8] ), .A3(_04750_ ), .ZN(_04880_ ) );
OR2_X1 _12604_ ( .A1(_04321_ ), .A2(\myreg.Reg[1][8] ), .ZN(_04881_ ) );
OAI211_X1 _12605_ ( .A(_04881_ ), .B(_04315_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[0][8] ), .ZN(_04882_ ) );
OR2_X1 _12606_ ( .A1(_04786_ ), .A2(\myreg.Reg[3][8] ), .ZN(_04883_ ) );
OAI211_X1 _12607_ ( .A(_04883_ ), .B(fanout_net_39 ), .C1(fanout_net_35 ), .C2(\myreg.Reg[2][8] ), .ZN(_04884_ ) );
NAND3_X1 _12608_ ( .A1(_04882_ ), .A2(_04884_ ), .A3(_04738_ ), .ZN(_04885_ ) );
MUX2_X1 _12609_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_36 ), .Z(_04886_ ) );
MUX2_X1 _12610_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_36 ), .Z(_04887_ ) );
MUX2_X1 _12611_ ( .A(_04886_ ), .B(_04887_ ), .S(_04315_ ), .Z(_04888_ ) );
OAI211_X1 _12612_ ( .A(_04310_ ), .B(_04885_ ), .C1(_04888_ ), .C2(_04337_ ), .ZN(_04889_ ) );
OR2_X1 _12613_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][8] ), .ZN(_04890_ ) );
OAI211_X1 _12614_ ( .A(_04890_ ), .B(fanout_net_39 ), .C1(_04392_ ), .C2(\myreg.Reg[15][8] ), .ZN(_04891_ ) );
OR2_X1 _12615_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[12][8] ), .ZN(_04892_ ) );
OAI211_X1 _12616_ ( .A(_04892_ ), .B(_04315_ ), .C1(_04392_ ), .C2(\myreg.Reg[13][8] ), .ZN(_04893_ ) );
NAND3_X1 _12617_ ( .A1(_04891_ ), .A2(_04893_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04894_ ) );
MUX2_X1 _12618_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_36 ), .Z(_04895_ ) );
MUX2_X1 _12619_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_36 ), .Z(_04896_ ) );
MUX2_X1 _12620_ ( .A(_04895_ ), .B(_04896_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04897_ ) );
OAI211_X1 _12621_ ( .A(fanout_net_41 ), .B(_04894_ ), .C1(_04897_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04898_ ) );
OAI211_X1 _12622_ ( .A(_04889_ ), .B(_04898_ ), .C1(_04302_ ), .C2(_04305_ ), .ZN(_04899_ ) );
NAND2_X1 _12623_ ( .A1(_04880_ ), .A2(_04899_ ), .ZN(_04900_ ) );
INV_X1 _12624_ ( .A(_04900_ ), .ZN(_04901_ ) );
XNOR2_X1 _12625_ ( .A(_03045_ ), .B(_04901_ ), .ZN(_04902_ ) );
OR2_X1 _12626_ ( .A1(_04320_ ), .A2(\myreg.Reg[1][9] ), .ZN(_04903_ ) );
OAI211_X1 _12627_ ( .A(_04903_ ), .B(_04791_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[0][9] ), .ZN(_04904_ ) );
OR2_X1 _12628_ ( .A1(_04320_ ), .A2(\myreg.Reg[3][9] ), .ZN(_04905_ ) );
OAI211_X1 _12629_ ( .A(_04905_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_36 ), .C2(\myreg.Reg[2][9] ), .ZN(_04906_ ) );
NAND3_X1 _12630_ ( .A1(_04904_ ), .A2(_04906_ ), .A3(_04335_ ), .ZN(_04907_ ) );
MUX2_X1 _12631_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_36 ), .Z(_04908_ ) );
MUX2_X1 _12632_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_36 ), .Z(_04909_ ) );
MUX2_X1 _12633_ ( .A(_04908_ ), .B(_04909_ ), .S(_04791_ ), .Z(_04910_ ) );
OAI211_X1 _12634_ ( .A(_04308_ ), .B(_04907_ ), .C1(_04910_ ), .C2(_04336_ ), .ZN(_04911_ ) );
OR2_X1 _12635_ ( .A1(_04320_ ), .A2(\myreg.Reg[13][9] ), .ZN(_04912_ ) );
OAI211_X1 _12636_ ( .A(_04912_ ), .B(_04791_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[12][9] ), .ZN(_04913_ ) );
OR2_X1 _12637_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][9] ), .ZN(_04914_ ) );
OAI211_X1 _12638_ ( .A(_04914_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04391_ ), .C2(\myreg.Reg[15][9] ), .ZN(_04915_ ) );
NAND3_X1 _12639_ ( .A1(_04913_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04915_ ), .ZN(_04916_ ) );
MUX2_X1 _12640_ ( .A(\myreg.Reg[8][9] ), .B(\myreg.Reg[9][9] ), .S(fanout_net_36 ), .Z(_04917_ ) );
MUX2_X1 _12641_ ( .A(\myreg.Reg[10][9] ), .B(\myreg.Reg[11][9] ), .S(fanout_net_36 ), .Z(_04918_ ) );
MUX2_X1 _12642_ ( .A(_04917_ ), .B(_04918_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04919_ ) );
OAI211_X1 _12643_ ( .A(fanout_net_41 ), .B(_04916_ ), .C1(_04919_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04920_ ) );
AOI21_X1 _12644_ ( .A(_04532_ ), .B1(_04911_ ), .B2(_04920_ ), .ZN(_04921_ ) );
INV_X1 _12645_ ( .A(\EX_LS_result_reg [9] ), .ZN(_04922_ ) );
NOR3_X1 _12646_ ( .A1(_04301_ ), .A2(_04922_ ), .A3(_04304_ ), .ZN(_04923_ ) );
NOR2_X1 _12647_ ( .A1(_04921_ ), .A2(_04923_ ), .ZN(_04924_ ) );
AND2_X1 _12648_ ( .A1(_04924_ ), .A2(_03068_ ), .ZN(_04925_ ) );
NOR2_X1 _12649_ ( .A1(_04924_ ), .A2(_03068_ ), .ZN(_04926_ ) );
NOR2_X1 _12650_ ( .A1(_04925_ ), .A2(_04926_ ), .ZN(_04927_ ) );
AND3_X1 _12651_ ( .A1(_04879_ ), .A2(_04902_ ), .A3(_04927_ ), .ZN(_04928_ ) );
AND2_X1 _12652_ ( .A1(_04829_ ), .A2(_04928_ ), .ZN(_04929_ ) );
INV_X1 _12653_ ( .A(_04929_ ), .ZN(_04930_ ) );
OR3_X1 _12654_ ( .A1(_04300_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02379_ ), .ZN(_04931_ ) );
OR2_X1 _12655_ ( .A1(_04320_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04932_ ) );
OAI211_X1 _12656_ ( .A(_04932_ ), .B(_04314_ ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04933_ ) );
OR2_X1 _12657_ ( .A1(_04320_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04934_ ) );
OAI211_X1 _12658_ ( .A(_04934_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04935_ ) );
NAND3_X1 _12659_ ( .A1(_04933_ ), .A2(_04935_ ), .A3(_04335_ ), .ZN(_04936_ ) );
MUX2_X1 _12660_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04937_ ) );
MUX2_X1 _12661_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04938_ ) );
MUX2_X1 _12662_ ( .A(_04937_ ), .B(_04938_ ), .S(_04791_ ), .Z(_04939_ ) );
OAI211_X1 _12663_ ( .A(_04308_ ), .B(_04936_ ), .C1(_04939_ ), .C2(_04336_ ), .ZN(_04940_ ) );
OR2_X1 _12664_ ( .A1(_04320_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04941_ ) );
OAI211_X1 _12665_ ( .A(_04941_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04942_ ) );
OR2_X1 _12666_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04943_ ) );
OAI211_X1 _12667_ ( .A(_04943_ ), .B(_04791_ ), .C1(_04786_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04944_ ) );
NAND3_X1 _12668_ ( .A1(_04942_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04944_ ), .ZN(_04945_ ) );
MUX2_X1 _12669_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04946_ ) );
MUX2_X1 _12670_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04947_ ) );
MUX2_X1 _12671_ ( .A(_04946_ ), .B(_04947_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04948_ ) );
OAI211_X1 _12672_ ( .A(fanout_net_41 ), .B(_04945_ ), .C1(_04948_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04949_ ) );
OAI211_X4 _12673_ ( .A(_04940_ ), .B(_04949_ ), .C1(_04301_ ), .C2(_04304_ ), .ZN(_04950_ ) );
NAND2_X1 _12674_ ( .A1(_04931_ ), .A2(_04950_ ), .ZN(_04951_ ) );
XNOR2_X1 _12675_ ( .A(_02910_ ), .B(_04951_ ), .ZN(_04952_ ) );
INV_X1 _12676_ ( .A(_04952_ ), .ZN(_04953_ ) );
INV_X1 _12677_ ( .A(\EX_LS_result_reg [0] ), .ZN(_04954_ ) );
OR3_X1 _12678_ ( .A1(_04301_ ), .A2(_04954_ ), .A3(_04304_ ), .ZN(_04955_ ) );
OR2_X1 _12679_ ( .A1(_04391_ ), .A2(\myreg.Reg[1][0] ), .ZN(_04956_ ) );
OAI211_X1 _12680_ ( .A(_04956_ ), .B(_04314_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[0][0] ), .ZN(_04957_ ) );
OR2_X1 _12681_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[2][0] ), .ZN(_04958_ ) );
OAI211_X1 _12682_ ( .A(_04958_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04321_ ), .C2(\myreg.Reg[3][0] ), .ZN(_04959_ ) );
NAND3_X1 _12683_ ( .A1(_04957_ ), .A2(_04336_ ), .A3(_04959_ ), .ZN(_04960_ ) );
MUX2_X1 _12684_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_36 ), .Z(_04961_ ) );
MUX2_X1 _12685_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_36 ), .Z(_04962_ ) );
MUX2_X1 _12686_ ( .A(_04961_ ), .B(_04962_ ), .S(_04791_ ), .Z(_04963_ ) );
OAI211_X1 _12687_ ( .A(_04309_ ), .B(_04960_ ), .C1(_04963_ ), .C2(_04748_ ), .ZN(_04964_ ) );
OR2_X1 _12688_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][0] ), .ZN(_04965_ ) );
OAI211_X1 _12689_ ( .A(_04965_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04321_ ), .C2(\myreg.Reg[15][0] ), .ZN(_04966_ ) );
OR2_X1 _12690_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[12][0] ), .ZN(_04967_ ) );
OAI211_X1 _12691_ ( .A(_04967_ ), .B(_04314_ ), .C1(_04786_ ), .C2(\myreg.Reg[13][0] ), .ZN(_04968_ ) );
NAND3_X1 _12692_ ( .A1(_04966_ ), .A2(_04968_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04969_ ) );
MUX2_X1 _12693_ ( .A(\myreg.Reg[8][0] ), .B(\myreg.Reg[9][0] ), .S(fanout_net_36 ), .Z(_04970_ ) );
MUX2_X1 _12694_ ( .A(\myreg.Reg[10][0] ), .B(\myreg.Reg[11][0] ), .S(fanout_net_36 ), .Z(_04971_ ) );
MUX2_X1 _12695_ ( .A(_04970_ ), .B(_04971_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04972_ ) );
OAI211_X1 _12696_ ( .A(fanout_net_41 ), .B(_04969_ ), .C1(_04972_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04973_ ) );
NAND2_X1 _12697_ ( .A1(_04964_ ), .A2(_04973_ ), .ZN(_04974_ ) );
OAI21_X2 _12698_ ( .A(_04974_ ), .B1(_04750_ ), .B2(_04775_ ), .ZN(_04975_ ) );
AND2_X1 _12699_ ( .A1(_04955_ ), .A2(_04975_ ), .ZN(_04976_ ) );
AND3_X1 _12700_ ( .A1(_04976_ ), .A2(_02859_ ), .A3(_02838_ ), .ZN(_04977_ ) );
OR3_X1 _12701_ ( .A1(_04775_ ), .A2(\EX_LS_result_reg [4] ), .A3(_04750_ ), .ZN(_04978_ ) );
OR2_X1 _12702_ ( .A1(_04321_ ), .A2(\myreg.Reg[1][4] ), .ZN(_04979_ ) );
OAI211_X1 _12703_ ( .A(_04979_ ), .B(_04315_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[0][4] ), .ZN(_04980_ ) );
OR2_X1 _12704_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][4] ), .ZN(_04981_ ) );
OAI211_X1 _12705_ ( .A(_04981_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04392_ ), .C2(\myreg.Reg[3][4] ), .ZN(_04982_ ) );
NAND3_X1 _12706_ ( .A1(_04980_ ), .A2(_04738_ ), .A3(_04982_ ), .ZN(_04983_ ) );
MUX2_X1 _12707_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_37 ), .Z(_04984_ ) );
MUX2_X1 _12708_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_37 ), .Z(_04985_ ) );
MUX2_X1 _12709_ ( .A(_04984_ ), .B(_04985_ ), .S(_04758_ ), .Z(_04986_ ) );
OAI211_X1 _12710_ ( .A(_04309_ ), .B(_04983_ ), .C1(_04986_ ), .C2(_04337_ ), .ZN(_04987_ ) );
OR2_X1 _12711_ ( .A1(_04786_ ), .A2(\myreg.Reg[15][4] ), .ZN(_04988_ ) );
OAI211_X1 _12712_ ( .A(_04988_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][4] ), .ZN(_04989_ ) );
OR2_X1 _12713_ ( .A1(_04786_ ), .A2(\myreg.Reg[13][4] ), .ZN(_04990_ ) );
OAI211_X1 _12714_ ( .A(_04990_ ), .B(_04315_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[12][4] ), .ZN(_04991_ ) );
NAND3_X1 _12715_ ( .A1(_04989_ ), .A2(_04991_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04992_ ) );
MUX2_X1 _12716_ ( .A(\myreg.Reg[8][4] ), .B(\myreg.Reg[9][4] ), .S(fanout_net_37 ), .Z(_04993_ ) );
MUX2_X1 _12717_ ( .A(\myreg.Reg[10][4] ), .B(\myreg.Reg[11][4] ), .S(fanout_net_37 ), .Z(_04994_ ) );
MUX2_X1 _12718_ ( .A(_04993_ ), .B(_04994_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04995_ ) );
OAI211_X1 _12719_ ( .A(fanout_net_41 ), .B(_04992_ ), .C1(_04995_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04996_ ) );
OAI211_X2 _12720_ ( .A(_04987_ ), .B(_04996_ ), .C1(_04302_ ), .C2(_04305_ ), .ZN(_04997_ ) );
NAND2_X2 _12721_ ( .A1(_04978_ ), .A2(_04997_ ), .ZN(_04998_ ) );
XOR2_X1 _12722_ ( .A(_02735_ ), .B(_04998_ ), .Z(_04999_ ) );
OR3_X4 _12723_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [2] ), .A3(_04304_ ), .ZN(_05000_ ) );
OR2_X1 _12724_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][2] ), .ZN(_05001_ ) );
OAI211_X1 _12725_ ( .A(_05001_ ), .B(_04758_ ), .C1(_04759_ ), .C2(\myreg.Reg[9][2] ), .ZN(_05002_ ) );
OR2_X1 _12726_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[10][2] ), .ZN(_05003_ ) );
OAI211_X1 _12727_ ( .A(_05003_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04759_ ), .C2(\myreg.Reg[11][2] ), .ZN(_05004_ ) );
NAND3_X1 _12728_ ( .A1(_05002_ ), .A2(_05004_ ), .A3(_04748_ ), .ZN(_05005_ ) );
MUX2_X1 _12729_ ( .A(\myreg.Reg[14][2] ), .B(\myreg.Reg[15][2] ), .S(fanout_net_37 ), .Z(_05006_ ) );
MUX2_X1 _12730_ ( .A(\myreg.Reg[12][2] ), .B(\myreg.Reg[13][2] ), .S(fanout_net_37 ), .Z(_05007_ ) );
MUX2_X1 _12731_ ( .A(_05006_ ), .B(_05007_ ), .S(_04730_ ), .Z(_05008_ ) );
OAI211_X1 _12732_ ( .A(fanout_net_41 ), .B(_05005_ ), .C1(_05008_ ), .C2(_04738_ ), .ZN(_05009_ ) );
OR2_X1 _12733_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][2] ), .ZN(_05010_ ) );
OAI211_X1 _12734_ ( .A(_05010_ ), .B(_04730_ ), .C1(_04759_ ), .C2(\myreg.Reg[1][2] ), .ZN(_05011_ ) );
NOR2_X1 _12735_ ( .A1(_04392_ ), .A2(\myreg.Reg[3][2] ), .ZN(_05012_ ) );
OAI21_X1 _12736_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_37 ), .B2(\myreg.Reg[2][2] ), .ZN(_05013_ ) );
OAI211_X1 _12737_ ( .A(_05011_ ), .B(_04336_ ), .C1(_05012_ ), .C2(_05013_ ), .ZN(_05014_ ) );
MUX2_X1 _12738_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_37 ), .Z(_05015_ ) );
MUX2_X1 _12739_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_37 ), .Z(_05016_ ) );
MUX2_X1 _12740_ ( .A(_05015_ ), .B(_05016_ ), .S(_04730_ ), .Z(_05017_ ) );
OAI211_X1 _12741_ ( .A(_04309_ ), .B(_05014_ ), .C1(_05017_ ), .C2(_04738_ ), .ZN(_05018_ ) );
OAI211_X1 _12742_ ( .A(_05009_ ), .B(_05018_ ), .C1(_04775_ ), .C2(_04750_ ), .ZN(_05019_ ) );
NAND2_X1 _12743_ ( .A1(_05000_ ), .A2(_05019_ ), .ZN(_05020_ ) );
INV_X1 _12744_ ( .A(_05020_ ), .ZN(_05021_ ) );
XNOR2_X1 _12745_ ( .A(_02886_ ), .B(_05021_ ), .ZN(_05022_ ) );
NAND2_X1 _12746_ ( .A1(_04999_ ), .A2(_05022_ ), .ZN(_05023_ ) );
NOR3_X1 _12747_ ( .A1(_04953_ ), .A2(_04977_ ), .A3(_05023_ ), .ZN(_05024_ ) );
OR3_X1 _12748_ ( .A1(_04404_ ), .A2(\EX_LS_result_reg [7] ), .A3(_04354_ ), .ZN(_05025_ ) );
OR2_X1 _12749_ ( .A1(_04393_ ), .A2(\myreg.Reg[5][7] ), .ZN(_05026_ ) );
OAI211_X1 _12750_ ( .A(_05026_ ), .B(_04317_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[4][7] ), .ZN(_05027_ ) );
OR2_X1 _12751_ ( .A1(_04393_ ), .A2(\myreg.Reg[7][7] ), .ZN(_05028_ ) );
OAI211_X1 _12752_ ( .A(_05028_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[6][7] ), .ZN(_05029_ ) );
NAND3_X1 _12753_ ( .A1(_05027_ ), .A2(_05029_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05030_ ) );
MUX2_X1 _12754_ ( .A(\myreg.Reg[2][7] ), .B(\myreg.Reg[3][7] ), .S(fanout_net_37 ), .Z(_05031_ ) );
MUX2_X1 _12755_ ( .A(\myreg.Reg[0][7] ), .B(\myreg.Reg[1][7] ), .S(fanout_net_37 ), .Z(_05032_ ) );
MUX2_X1 _12756_ ( .A(_05031_ ), .B(_05032_ ), .S(_04331_ ), .Z(_05033_ ) );
OAI211_X1 _12757_ ( .A(_04310_ ), .B(_05030_ ), .C1(_05033_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05034_ ) );
NOR2_X1 _12758_ ( .A1(_04323_ ), .A2(\myreg.Reg[11][7] ), .ZN(_05035_ ) );
OAI21_X1 _12759_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_37 ), .B2(\myreg.Reg[10][7] ), .ZN(_05036_ ) );
NOR2_X1 _12760_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][7] ), .ZN(_05037_ ) );
OAI21_X1 _12761_ ( .A(_04331_ ), .B1(_04323_ ), .B2(\myreg.Reg[9][7] ), .ZN(_05038_ ) );
OAI221_X1 _12762_ ( .A(_04402_ ), .B1(_05035_ ), .B2(_05036_ ), .C1(_05037_ ), .C2(_05038_ ), .ZN(_05039_ ) );
MUX2_X1 _12763_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_37 ), .Z(_05040_ ) );
MUX2_X1 _12764_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_37 ), .Z(_05041_ ) );
MUX2_X1 _12765_ ( .A(_05040_ ), .B(_05041_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_05042_ ) );
OAI211_X1 _12766_ ( .A(fanout_net_41 ), .B(_05039_ ), .C1(_05042_ ), .C2(_04338_ ), .ZN(_05043_ ) );
OAI211_X1 _12767_ ( .A(_05034_ ), .B(_05043_ ), .C1(_04404_ ), .C2(_04306_ ), .ZN(_05044_ ) );
NAND2_X1 _12768_ ( .A1(_05025_ ), .A2(_05044_ ), .ZN(_05045_ ) );
INV_X1 _12769_ ( .A(_05045_ ), .ZN(_05046_ ) );
XNOR2_X1 _12770_ ( .A(_02812_ ), .B(_05046_ ), .ZN(_05047_ ) );
INV_X1 _12771_ ( .A(_05047_ ), .ZN(_05048_ ) );
OR3_X1 _12772_ ( .A1(_04302_ ), .A2(\EX_LS_result_reg [6] ), .A3(_04305_ ), .ZN(_05049_ ) );
OR2_X1 _12773_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][6] ), .ZN(_05050_ ) );
OAI211_X1 _12774_ ( .A(_05050_ ), .B(_04331_ ), .C1(_04339_ ), .C2(\myreg.Reg[1][6] ), .ZN(_05051_ ) );
OR2_X1 _12775_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][6] ), .ZN(_05052_ ) );
OAI211_X1 _12776_ ( .A(_05052_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04339_ ), .C2(\myreg.Reg[3][6] ), .ZN(_05053_ ) );
NAND3_X1 _12777_ ( .A1(_05051_ ), .A2(_05053_ ), .A3(_04402_ ), .ZN(_05054_ ) );
MUX2_X1 _12778_ ( .A(\myreg.Reg[6][6] ), .B(\myreg.Reg[7][6] ), .S(fanout_net_37 ), .Z(_05055_ ) );
MUX2_X1 _12779_ ( .A(\myreg.Reg[4][6] ), .B(\myreg.Reg[5][6] ), .S(fanout_net_37 ), .Z(_05056_ ) );
MUX2_X1 _12780_ ( .A(_05055_ ), .B(_05056_ ), .S(_04316_ ), .Z(_05057_ ) );
OAI211_X1 _12781_ ( .A(_04310_ ), .B(_05054_ ), .C1(_05057_ ), .C2(_04402_ ), .ZN(_05058_ ) );
OR2_X1 _12782_ ( .A1(_04322_ ), .A2(\myreg.Reg[15][6] ), .ZN(_05059_ ) );
OAI211_X1 _12783_ ( .A(_05059_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][6] ), .ZN(_05060_ ) );
OR2_X1 _12784_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][6] ), .ZN(_05061_ ) );
OAI211_X1 _12785_ ( .A(_05061_ ), .B(_04331_ ), .C1(_04393_ ), .C2(\myreg.Reg[13][6] ), .ZN(_05062_ ) );
NAND3_X1 _12786_ ( .A1(_05060_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_05062_ ), .ZN(_05063_ ) );
MUX2_X1 _12787_ ( .A(\myreg.Reg[8][6] ), .B(\myreg.Reg[9][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05064_ ) );
MUX2_X1 _12788_ ( .A(\myreg.Reg[10][6] ), .B(\myreg.Reg[11][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05065_ ) );
MUX2_X1 _12789_ ( .A(_05064_ ), .B(_05065_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_05066_ ) );
OAI211_X1 _12790_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05063_ ), .C1(_05066_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05067_ ) );
OAI211_X1 _12791_ ( .A(_05058_ ), .B(_05067_ ), .C1(_04404_ ), .C2(_04354_ ), .ZN(_05068_ ) );
NAND2_X2 _12792_ ( .A1(_05049_ ), .A2(_05068_ ), .ZN(_05069_ ) );
XNOR2_X1 _12793_ ( .A(_02788_ ), .B(_05069_ ), .ZN(_05070_ ) );
NOR2_X1 _12794_ ( .A1(_05048_ ), .A2(_05070_ ), .ZN(_05071_ ) );
OR2_X1 _12795_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05072_ ) );
OAI211_X1 _12796_ ( .A(_05072_ ), .B(_04730_ ), .C1(_04321_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05073_ ) );
OR2_X1 _12797_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_05074_ ) );
OAI211_X1 _12798_ ( .A(_05074_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04321_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05075_ ) );
NAND3_X1 _12799_ ( .A1(_05073_ ), .A2(_05075_ ), .A3(_04336_ ), .ZN(_05076_ ) );
MUX2_X1 _12800_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05077_ ) );
MUX2_X1 _12801_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05078_ ) );
MUX2_X1 _12802_ ( .A(_05077_ ), .B(_05078_ ), .S(_04314_ ), .Z(_05079_ ) );
OAI211_X1 _12803_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05076_ ), .C1(_05079_ ), .C2(_04738_ ), .ZN(_05080_ ) );
NOR2_X1 _12804_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05081_ ) );
AOI211_X1 _12805_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B(_05081_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(_02742_ ), .ZN(_05082_ ) );
MUX2_X1 _12806_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05083_ ) );
AOI211_X1 _12807_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_05082_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C2(_05083_ ), .ZN(_05084_ ) );
MUX2_X1 _12808_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05085_ ) );
MUX2_X1 _12809_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05086_ ) );
MUX2_X1 _12810_ ( .A(_05085_ ), .B(_05086_ ), .S(_04791_ ), .Z(_05087_ ) );
OAI21_X1 _12811_ ( .A(_04309_ ), .B1(_05087_ ), .B2(_04748_ ), .ZN(_05088_ ) );
OAI221_X2 _12812_ ( .A(_05080_ ), .B1(_05084_ ), .B2(_05088_ ), .C1(_04775_ ), .C2(_04750_ ), .ZN(_05089_ ) );
OR3_X4 _12813_ ( .A1(_04301_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04304_ ), .ZN(_05090_ ) );
NAND2_X4 _12814_ ( .A1(_05089_ ), .A2(_05090_ ), .ZN(_05091_ ) );
XNOR2_X1 _12815_ ( .A(_02764_ ), .B(_05091_ ), .ZN(_05092_ ) );
OR3_X4 _12816_ ( .A1(_04301_ ), .A2(\EX_LS_result_reg [1] ), .A3(_04304_ ), .ZN(_05093_ ) );
OR2_X1 _12817_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[4][1] ), .ZN(_05094_ ) );
OAI211_X1 _12818_ ( .A(_05094_ ), .B(_04730_ ), .C1(_04321_ ), .C2(\myreg.Reg[5][1] ), .ZN(_05095_ ) );
OR2_X1 _12819_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[6][1] ), .ZN(_05096_ ) );
OAI211_X1 _12820_ ( .A(_05096_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04321_ ), .C2(\myreg.Reg[7][1] ), .ZN(_05097_ ) );
NAND3_X1 _12821_ ( .A1(_05095_ ), .A2(_05097_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05098_ ) );
MUX2_X1 _12822_ ( .A(\myreg.Reg[2][1] ), .B(\myreg.Reg[3][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05099_ ) );
MUX2_X1 _12823_ ( .A(\myreg.Reg[0][1] ), .B(\myreg.Reg[1][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05100_ ) );
MUX2_X1 _12824_ ( .A(_05099_ ), .B(_05100_ ), .S(_04314_ ), .Z(_05101_ ) );
OAI211_X1 _12825_ ( .A(_04309_ ), .B(_05098_ ), .C1(_05101_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05102_ ) );
NOR2_X1 _12826_ ( .A1(_04786_ ), .A2(\myreg.Reg[11][1] ), .ZN(_05103_ ) );
OAI21_X1 _12827_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myreg.Reg[10][1] ), .ZN(_05104_ ) );
NOR2_X1 _12828_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[8][1] ), .ZN(_05105_ ) );
OAI21_X1 _12829_ ( .A(_04314_ ), .B1(_04786_ ), .B2(\myreg.Reg[9][1] ), .ZN(_05106_ ) );
OAI221_X1 _12830_ ( .A(_04335_ ), .B1(_05103_ ), .B2(_05104_ ), .C1(_05105_ ), .C2(_05106_ ), .ZN(_05107_ ) );
MUX2_X1 _12831_ ( .A(\myreg.Reg[12][1] ), .B(\myreg.Reg[13][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05108_ ) );
MUX2_X1 _12832_ ( .A(\myreg.Reg[14][1] ), .B(\myreg.Reg[15][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05109_ ) );
MUX2_X1 _12833_ ( .A(_05108_ ), .B(_05109_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_05110_ ) );
OAI211_X1 _12834_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05107_ ), .C1(_05110_ ), .C2(_04748_ ), .ZN(_05111_ ) );
OAI211_X2 _12835_ ( .A(_05102_ ), .B(_05111_ ), .C1(_04775_ ), .C2(_04750_ ), .ZN(_05112_ ) );
NAND2_X4 _12836_ ( .A1(_05093_ ), .A2(_05112_ ), .ZN(_05113_ ) );
INV_X1 _12837_ ( .A(_05113_ ), .ZN(_05114_ ) );
XNOR2_X1 _12838_ ( .A(_02835_ ), .B(_05114_ ), .ZN(_05115_ ) );
AND2_X4 _12839_ ( .A1(_02838_ ), .A2(_02859_ ), .ZN(_05116_ ) );
NOR2_X1 _12840_ ( .A1(_05116_ ), .A2(_04976_ ), .ZN(_05117_ ) );
INV_X1 _12841_ ( .A(_05117_ ), .ZN(_05118_ ) );
AND2_X1 _12842_ ( .A1(_05115_ ), .A2(_05118_ ), .ZN(_05119_ ) );
NAND4_X1 _12843_ ( .A1(_05024_ ), .A2(_05071_ ), .A3(_05092_ ), .A4(_05119_ ), .ZN(_05120_ ) );
NOR2_X1 _12844_ ( .A1(_04930_ ), .A2(_05120_ ), .ZN(_05121_ ) );
NAND2_X1 _12845_ ( .A1(_04727_ ), .A2(_05121_ ), .ZN(_05122_ ) );
NOR2_X1 _12846_ ( .A1(_04146_ ), .A2(\ID_EX_typ [1] ), .ZN(_05123_ ) );
AND2_X1 _12847_ ( .A1(_05123_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05124_ ) );
INV_X1 _12848_ ( .A(\ID_EX_typ [1] ), .ZN(_05125_ ) );
NOR2_X1 _12849_ ( .A1(_05125_ ), .A2(fanout_net_7 ), .ZN(_05126_ ) );
INV_X1 _12850_ ( .A(\ID_EX_typ [2] ), .ZN(_05127_ ) );
AND2_X1 _12851_ ( .A1(_05126_ ), .A2(_05127_ ), .ZN(_05128_ ) );
BUF_X4 _12852_ ( .A(_05128_ ), .Z(_05129_ ) );
INV_X1 _12853_ ( .A(_05129_ ), .ZN(_05130_ ) );
NAND2_X1 _12854_ ( .A1(_04291_ ), .A2(\ID_EX_typ [2] ), .ZN(_05131_ ) );
OR2_X1 _12855_ ( .A1(_04629_ ), .A2(fanout_net_8 ), .ZN(_05132_ ) );
INV_X1 _12856_ ( .A(\ID_EX_imm [31] ), .ZN(_05133_ ) );
NAND2_X1 _12857_ ( .A1(_05133_ ), .A2(fanout_net_8 ), .ZN(_05134_ ) );
NAND2_X1 _12858_ ( .A1(_05132_ ), .A2(_05134_ ), .ZN(_05135_ ) );
INV_X1 _12859_ ( .A(_03243_ ), .ZN(_05136_ ) );
NAND2_X1 _12860_ ( .A1(_05135_ ), .A2(_05136_ ), .ZN(_05137_ ) );
NAND3_X1 _12861_ ( .A1(_05132_ ), .A2(_03243_ ), .A3(_05134_ ), .ZN(_05138_ ) );
NAND2_X1 _12862_ ( .A1(_05137_ ), .A2(_05138_ ), .ZN(_05139_ ) );
INV_X1 _12863_ ( .A(_05139_ ), .ZN(_05140_ ) );
INV_X1 _12864_ ( .A(fanout_net_8 ), .ZN(_05141_ ) );
BUF_X4 _12865_ ( .A(_05141_ ), .Z(_05142_ ) );
BUF_X4 _12866_ ( .A(_05142_ ), .Z(_05143_ ) );
BUF_X2 _12867_ ( .A(_05143_ ), .Z(_05144_ ) );
NAND3_X1 _12868_ ( .A1(_04586_ ), .A2(_05144_ ), .A3(_04604_ ), .ZN(_05145_ ) );
NAND2_X1 _12869_ ( .A1(fanout_net_8 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05146_ ) );
AND2_X1 _12870_ ( .A1(_05145_ ), .A2(_05146_ ), .ZN(_05147_ ) );
XNOR2_X1 _12871_ ( .A(_02401_ ), .B(_05147_ ), .ZN(_05148_ ) );
NOR2_X1 _12872_ ( .A1(_05140_ ), .A2(_05148_ ), .ZN(_05149_ ) );
INV_X1 _12873_ ( .A(_05149_ ), .ZN(_05150_ ) );
NAND2_X1 _12874_ ( .A1(_04581_ ), .A2(_05144_ ), .ZN(_05151_ ) );
NAND2_X1 _12875_ ( .A1(_03219_ ), .A2(fanout_net_8 ), .ZN(_05152_ ) );
NAND2_X1 _12876_ ( .A1(_05151_ ), .A2(_05152_ ), .ZN(_05153_ ) );
AND2_X1 _12877_ ( .A1(_05153_ ), .A2(_02425_ ), .ZN(_05154_ ) );
NOR2_X1 _12878_ ( .A1(_05153_ ), .A2(_02425_ ), .ZN(_05155_ ) );
NOR2_X1 _12879_ ( .A1(_05154_ ), .A2(_05155_ ), .ZN(_05156_ ) );
OR2_X1 _12880_ ( .A1(_04559_ ), .A2(fanout_net_8 ), .ZN(_05157_ ) );
NAND2_X1 _12881_ ( .A1(fanout_net_8 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05158_ ) );
AND2_X2 _12882_ ( .A1(_05157_ ), .A2(_05158_ ), .ZN(_05159_ ) );
INV_X1 _12883_ ( .A(_02448_ ), .ZN(_05160_ ) );
XNOR2_X1 _12884_ ( .A(_05159_ ), .B(_05160_ ), .ZN(_05161_ ) );
OR3_X1 _12885_ ( .A1(_05150_ ), .A2(_05156_ ), .A3(_05161_ ), .ZN(_05162_ ) );
NAND2_X1 _12886_ ( .A1(_04752_ ), .A2(_05142_ ), .ZN(_05163_ ) );
OR2_X1 _12887_ ( .A1(_05141_ ), .A2(\ID_EX_imm [14] ), .ZN(_05164_ ) );
NAND2_X4 _12888_ ( .A1(_05163_ ), .A2(_05164_ ), .ZN(_05165_ ) );
XNOR2_X2 _12889_ ( .A(_05165_ ), .B(_03020_ ), .ZN(_05166_ ) );
INV_X2 _12890_ ( .A(_05166_ ), .ZN(_05167_ ) );
NAND3_X1 _12891_ ( .A1(_04754_ ), .A2(_05142_ ), .A3(_04776_ ), .ZN(_05168_ ) );
NAND2_X1 _12892_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [15] ), .ZN(_05169_ ) );
AND2_X4 _12893_ ( .A1(_05168_ ), .A2(_05169_ ), .ZN(_05170_ ) );
XNOR2_X2 _12894_ ( .A(_05170_ ), .B(_02996_ ), .ZN(_05171_ ) );
INV_X2 _12895_ ( .A(_05171_ ), .ZN(_05172_ ) );
NAND3_X1 _12896_ ( .A1(_04807_ ), .A2(_04826_ ), .A3(_05142_ ), .ZN(_05173_ ) );
NAND2_X1 _12897_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [12] ), .ZN(_05174_ ) );
AND2_X4 _12898_ ( .A1(_05173_ ), .A2(_05174_ ), .ZN(_05175_ ) );
XNOR2_X2 _12899_ ( .A(_05175_ ), .B(_02948_ ), .ZN(_05176_ ) );
INV_X2 _12900_ ( .A(_05176_ ), .ZN(_05177_ ) );
NAND3_X2 _12901_ ( .A1(_05167_ ), .A2(_05172_ ), .A3(_05177_ ), .ZN(_05178_ ) );
NAND3_X1 _12902_ ( .A1(_04782_ ), .A2(_05141_ ), .A3(_04803_ ), .ZN(_05179_ ) );
NAND2_X1 _12903_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [13] ), .ZN(_05180_ ) );
AND2_X1 _12904_ ( .A1(_05179_ ), .A2(_05180_ ), .ZN(_05181_ ) );
XNOR2_X2 _12905_ ( .A(_05181_ ), .B(_04781_ ), .ZN(_05182_ ) );
NOR2_X4 _12906_ ( .A1(_05178_ ), .A2(_05182_ ), .ZN(_05183_ ) );
OR2_X1 _12907_ ( .A1(_04852_ ), .A2(fanout_net_8 ), .ZN(_05184_ ) );
NAND2_X1 _12908_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [11] ), .ZN(_05185_ ) );
AND2_X1 _12909_ ( .A1(_05184_ ), .A2(_05185_ ), .ZN(_05186_ ) );
INV_X1 _12910_ ( .A(_04854_ ), .ZN(_05187_ ) );
NOR2_X2 _12911_ ( .A1(_05186_ ), .A2(_05187_ ), .ZN(_05188_ ) );
AND3_X1 _12912_ ( .A1(_05184_ ), .A2(_05187_ ), .A3(_05185_ ), .ZN(_05189_ ) );
NOR2_X1 _12913_ ( .A1(_05188_ ), .A2(_05189_ ), .ZN(_05190_ ) );
INV_X1 _12914_ ( .A(_05190_ ), .ZN(_05191_ ) );
NAND3_X1 _12915_ ( .A1(_04856_ ), .A2(_05142_ ), .A3(_04875_ ), .ZN(_05192_ ) );
NAND2_X1 _12916_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [10] ), .ZN(_05193_ ) );
AND2_X2 _12917_ ( .A1(_05192_ ), .A2(_05193_ ), .ZN(_05194_ ) );
XNOR2_X2 _12918_ ( .A(_05194_ ), .B(_03095_ ), .ZN(_05195_ ) );
INV_X4 _12919_ ( .A(_05195_ ), .ZN(_05196_ ) );
NAND3_X1 _12920_ ( .A1(_05183_ ), .A2(_05191_ ), .A3(_05196_ ), .ZN(_05197_ ) );
OAI21_X1 _12921_ ( .A(_05141_ ), .B1(_04921_ ), .B2(_04923_ ), .ZN(_05198_ ) );
NAND2_X1 _12922_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [9] ), .ZN(_05199_ ) );
AND2_X1 _12923_ ( .A1(_05198_ ), .A2(_05199_ ), .ZN(_05200_ ) );
INV_X2 _12924_ ( .A(_03068_ ), .ZN(_05201_ ) );
NOR2_X2 _12925_ ( .A1(_05200_ ), .A2(_05201_ ), .ZN(_05202_ ) );
AND3_X4 _12926_ ( .A1(_05201_ ), .A2(_05199_ ), .A3(_05198_ ), .ZN(_05203_ ) );
NOR2_X4 _12927_ ( .A1(_05202_ ), .A2(_05203_ ), .ZN(_05204_ ) );
NAND3_X1 _12928_ ( .A1(_04880_ ), .A2(_05142_ ), .A3(_04899_ ), .ZN(_05205_ ) );
NAND2_X1 _12929_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [8] ), .ZN(_05206_ ) );
AND2_X1 _12930_ ( .A1(_05205_ ), .A2(_05206_ ), .ZN(_05207_ ) );
XNOR2_X1 _12931_ ( .A(_05207_ ), .B(_03045_ ), .ZN(_05208_ ) );
NOR3_X2 _12932_ ( .A1(_05197_ ), .A2(_05204_ ), .A3(_05208_ ), .ZN(_05209_ ) );
NAND2_X1 _12933_ ( .A1(_05091_ ), .A2(_05142_ ), .ZN(_05210_ ) );
NAND2_X1 _12934_ ( .A1(_02921_ ), .A2(fanout_net_8 ), .ZN(_05211_ ) );
NAND2_X2 _12935_ ( .A1(_05210_ ), .A2(_05211_ ), .ZN(_05212_ ) );
INV_X4 _12936_ ( .A(_02764_ ), .ZN(_05213_ ) );
XNOR2_X2 _12937_ ( .A(_05212_ ), .B(_05213_ ), .ZN(_05214_ ) );
NAND2_X2 _12938_ ( .A1(_04998_ ), .A2(_05143_ ), .ZN(_05215_ ) );
NAND2_X1 _12939_ ( .A1(_02736_ ), .A2(fanout_net_8 ), .ZN(_05216_ ) );
NAND2_X2 _12940_ ( .A1(_05215_ ), .A2(_05216_ ), .ZN(_05217_ ) );
NOR2_X2 _12941_ ( .A1(_05217_ ), .A2(_02919_ ), .ZN(_05218_ ) );
AOI21_X2 _12942_ ( .A(_02735_ ), .B1(_05215_ ), .B2(_05216_ ), .ZN(_05219_ ) );
NOR2_X1 _12943_ ( .A1(_05218_ ), .A2(_05219_ ), .ZN(_05220_ ) );
NAND3_X1 _12944_ ( .A1(_04931_ ), .A2(_05141_ ), .A3(_04950_ ), .ZN(_05221_ ) );
NAND2_X1 _12945_ ( .A1(fanout_net_8 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_05222_ ) );
AND2_X2 _12946_ ( .A1(_05221_ ), .A2(_05222_ ), .ZN(_05223_ ) );
AND2_X4 _12947_ ( .A1(_02910_ ), .A2(_05223_ ), .ZN(_05224_ ) );
NOR2_X2 _12948_ ( .A1(_02910_ ), .A2(_05223_ ), .ZN(_05225_ ) );
NOR2_X4 _12949_ ( .A1(_05224_ ), .A2(_05225_ ), .ZN(_05226_ ) );
INV_X1 _12950_ ( .A(_02886_ ), .ZN(_05227_ ) );
NAND3_X1 _12951_ ( .A1(_05000_ ), .A2(_05019_ ), .A3(_05142_ ), .ZN(_05228_ ) );
NAND2_X1 _12952_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [2] ), .ZN(_05229_ ) );
AND2_X4 _12953_ ( .A1(_05228_ ), .A2(_05229_ ), .ZN(_05230_ ) );
INV_X2 _12954_ ( .A(_05230_ ), .ZN(_05231_ ) );
NOR3_X1 _12955_ ( .A1(_05226_ ), .A2(_05227_ ), .A3(_05231_ ), .ZN(_05232_ ) );
INV_X1 _12956_ ( .A(_05223_ ), .ZN(_05233_ ) );
AOI21_X1 _12957_ ( .A(_05232_ ), .B1(_02910_ ), .B2(_05233_ ), .ZN(_05234_ ) );
NAND2_X2 _12958_ ( .A1(_05113_ ), .A2(_05142_ ), .ZN(_05235_ ) );
NAND2_X1 _12959_ ( .A1(_02836_ ), .A2(fanout_net_8 ), .ZN(_05236_ ) );
NAND2_X4 _12960_ ( .A1(_05235_ ), .A2(_05236_ ), .ZN(_05237_ ) );
NAND2_X1 _12961_ ( .A1(_05237_ ), .A2(_02835_ ), .ZN(_05238_ ) );
XNOR2_X2 _12962_ ( .A(_05237_ ), .B(_02835_ ), .ZN(_05239_ ) );
NAND3_X2 _12963_ ( .A1(_04955_ ), .A2(_04975_ ), .A3(_05142_ ), .ZN(_05240_ ) );
OR2_X1 _12964_ ( .A1(_05141_ ), .A2(\ID_EX_imm [0] ), .ZN(_05241_ ) );
NAND2_X4 _12965_ ( .A1(_05240_ ), .A2(_05241_ ), .ZN(_05242_ ) );
NOR2_X4 _12966_ ( .A1(_05242_ ), .A2(_05116_ ), .ZN(_05243_ ) );
OAI21_X2 _12967_ ( .A(_05238_ ), .B1(_05239_ ), .B2(_05243_ ), .ZN(_05244_ ) );
XNOR2_X2 _12968_ ( .A(_05230_ ), .B(_02886_ ), .ZN(_05245_ ) );
INV_X1 _12969_ ( .A(_05245_ ), .ZN(_05246_ ) );
OAI211_X1 _12970_ ( .A(_05244_ ), .B(_05246_ ), .C1(_05224_ ), .C2(_05225_ ), .ZN(_05247_ ) );
AOI211_X1 _12971_ ( .A(_05214_ ), .B(_05220_ ), .C1(_05234_ ), .C2(_05247_ ), .ZN(_05248_ ) );
AND3_X1 _12972_ ( .A1(_05210_ ), .A2(_02764_ ), .A3(_05211_ ), .ZN(_05249_ ) );
INV_X1 _12973_ ( .A(_05217_ ), .ZN(_05250_ ) );
NOR3_X1 _12974_ ( .A1(_05214_ ), .A2(_02919_ ), .A3(_05250_ ), .ZN(_05251_ ) );
NOR3_X1 _12975_ ( .A1(_05248_ ), .A2(_05249_ ), .A3(_05251_ ), .ZN(_05252_ ) );
NAND3_X1 _12976_ ( .A1(_05025_ ), .A2(_05143_ ), .A3(_05044_ ), .ZN(_05253_ ) );
NAND2_X1 _12977_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [7] ), .ZN(_05254_ ) );
AND2_X2 _12978_ ( .A1(_05253_ ), .A2(_05254_ ), .ZN(_05255_ ) );
XNOR2_X1 _12979_ ( .A(_05255_ ), .B(_02812_ ), .ZN(_05256_ ) );
NAND2_X1 _12980_ ( .A1(_05069_ ), .A2(_05143_ ), .ZN(_05257_ ) );
OR2_X1 _12981_ ( .A1(_05143_ ), .A2(\ID_EX_imm [6] ), .ZN(_05258_ ) );
NAND2_X1 _12982_ ( .A1(_05257_ ), .A2(_05258_ ), .ZN(_05259_ ) );
XNOR2_X1 _12983_ ( .A(_05259_ ), .B(_02788_ ), .ZN(_05260_ ) );
NOR3_X2 _12984_ ( .A1(_05252_ ), .A2(_05256_ ), .A3(_05260_ ), .ZN(_05261_ ) );
INV_X1 _12985_ ( .A(_02811_ ), .ZN(_05262_ ) );
AND2_X1 _12986_ ( .A1(_05255_ ), .A2(_05262_ ), .ZN(_05263_ ) );
NOR2_X1 _12987_ ( .A1(_05255_ ), .A2(_05262_ ), .ZN(_05264_ ) );
OAI211_X1 _12988_ ( .A(_02788_ ), .B(_05259_ ), .C1(_05263_ ), .C2(_05264_ ), .ZN(_05265_ ) );
INV_X1 _12989_ ( .A(_05255_ ), .ZN(_05266_ ) );
OAI21_X1 _12990_ ( .A(_05265_ ), .B1(_05262_ ), .B2(_05266_ ), .ZN(_05267_ ) );
OAI21_X1 _12991_ ( .A(_05209_ ), .B1(_05261_ ), .B2(_05267_ ), .ZN(_05268_ ) );
NAND3_X1 _12992_ ( .A1(_05172_ ), .A2(_03020_ ), .A3(_05165_ ), .ZN(_05269_ ) );
INV_X1 _12993_ ( .A(_02948_ ), .ZN(_05270_ ) );
INV_X1 _12994_ ( .A(_05175_ ), .ZN(_05271_ ) );
NOR3_X1 _12995_ ( .A1(_05182_ ), .A2(_05270_ ), .A3(_05271_ ), .ZN(_05272_ ) );
AND4_X1 _12996_ ( .A1(_02970_ ), .A2(_05179_ ), .A3(_02950_ ), .A4(_05180_ ), .ZN(_05273_ ) );
NOR2_X1 _12997_ ( .A1(_05272_ ), .A2(_05273_ ), .ZN(_05274_ ) );
NOR3_X1 _12998_ ( .A1(_05274_ ), .A2(_05171_ ), .A3(_05166_ ), .ZN(_05275_ ) );
NAND3_X1 _12999_ ( .A1(_05191_ ), .A2(_03095_ ), .A3(_05194_ ), .ZN(_05276_ ) );
INV_X1 _13000_ ( .A(_05186_ ), .ZN(_05277_ ) );
INV_X1 _13001_ ( .A(_03045_ ), .ZN(_05278_ ) );
INV_X1 _13002_ ( .A(_05207_ ), .ZN(_05279_ ) );
NOR3_X2 _13003_ ( .A1(_05204_ ), .A2(_05278_ ), .A3(_05279_ ), .ZN(_05280_ ) );
AOI21_X1 _13004_ ( .A(_05280_ ), .B1(_03068_ ), .B2(_05200_ ), .ZN(_05281_ ) );
OAI21_X1 _13005_ ( .A(_05196_ ), .B1(_05188_ ), .B2(_05189_ ), .ZN(_05282_ ) );
OAI221_X1 _13006_ ( .A(_05276_ ), .B1(_05187_ ), .B2(_05277_ ), .C1(_05281_ ), .C2(_05282_ ), .ZN(_05283_ ) );
AOI221_X2 _13007_ ( .A(_05275_ ), .B1(_02996_ ), .B2(_05170_ ), .C1(_05283_ ), .C2(_05183_ ), .ZN(_05284_ ) );
AND3_X2 _13008_ ( .A1(_05268_ ), .A2(_05269_ ), .A3(_05284_ ), .ZN(_05285_ ) );
NAND3_X1 _13009_ ( .A1(_04355_ ), .A2(_05144_ ), .A3(_04374_ ), .ZN(_05286_ ) );
NAND2_X1 _13010_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [17] ), .ZN(_05287_ ) );
AND2_X1 _13011_ ( .A1(_05286_ ), .A2(_05287_ ), .ZN(_05288_ ) );
XNOR2_X1 _13012_ ( .A(_05288_ ), .B(_02684_ ), .ZN(_05289_ ) );
NAND2_X1 _13013_ ( .A1(_04352_ ), .A2(_05144_ ), .ZN(_05290_ ) );
NAND2_X1 _13014_ ( .A1(_02710_ ), .A2(fanout_net_8 ), .ZN(_05291_ ) );
NAND2_X1 _13015_ ( .A1(_05290_ ), .A2(_05291_ ), .ZN(_05292_ ) );
XNOR2_X1 _13016_ ( .A(_05292_ ), .B(_02709_ ), .ZN(_05293_ ) );
NAND2_X2 _13017_ ( .A1(_04454_ ), .A2(_05143_ ), .ZN(_05294_ ) );
NAND2_X1 _13018_ ( .A1(_02536_ ), .A2(fanout_net_8 ), .ZN(_05295_ ) );
NAND2_X4 _13019_ ( .A1(_05294_ ), .A2(_05295_ ), .ZN(_05296_ ) );
XNOR2_X2 _13020_ ( .A(_05296_ ), .B(_02535_ ), .ZN(_05297_ ) );
INV_X4 _13021_ ( .A(_05297_ ), .ZN(_05298_ ) );
NAND3_X1 _13022_ ( .A1(_04506_ ), .A2(_05143_ ), .A3(_04525_ ), .ZN(_05299_ ) );
NAND2_X1 _13023_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [21] ), .ZN(_05300_ ) );
AND2_X4 _13024_ ( .A1(_05299_ ), .A2(_05300_ ), .ZN(_05301_ ) );
XNOR2_X2 _13025_ ( .A(_05301_ ), .B(_04505_ ), .ZN(_05302_ ) );
INV_X2 _13026_ ( .A(_05302_ ), .ZN(_05303_ ) );
OR2_X4 _13027_ ( .A1(_04479_ ), .A2(fanout_net_8 ), .ZN(_05304_ ) );
NAND2_X1 _13028_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [23] ), .ZN(_05305_ ) );
AND2_X1 _13029_ ( .A1(_05304_ ), .A2(_05305_ ), .ZN(_05306_ ) );
INV_X2 _13030_ ( .A(_02561_ ), .ZN(_05307_ ) );
NOR2_X2 _13031_ ( .A1(_05306_ ), .A2(_05307_ ), .ZN(_05308_ ) );
AND3_X2 _13032_ ( .A1(_05304_ ), .A2(_05307_ ), .A3(_05305_ ), .ZN(_05309_ ) );
OAI211_X1 _13033_ ( .A(_05298_ ), .B(_05303_ ), .C1(_05308_ ), .C2(_05309_ ), .ZN(_05310_ ) );
NAND3_X1 _13034_ ( .A1(_04483_ ), .A2(_04502_ ), .A3(_05143_ ), .ZN(_05311_ ) );
NAND2_X1 _13035_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [20] ), .ZN(_05312_ ) );
AND2_X2 _13036_ ( .A1(_05311_ ), .A2(_05312_ ), .ZN(_05313_ ) );
XNOR2_X1 _13037_ ( .A(_05313_ ), .B(_02610_ ), .ZN(_05314_ ) );
NAND3_X2 _13038_ ( .A1(_04409_ ), .A2(_05143_ ), .A3(_04428_ ), .ZN(_05315_ ) );
NAND2_X1 _13039_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [18] ), .ZN(_05316_ ) );
AND2_X4 _13040_ ( .A1(_05315_ ), .A2(_05316_ ), .ZN(_05317_ ) );
XNOR2_X2 _13041_ ( .A(_05317_ ), .B(_02634_ ), .ZN(_05318_ ) );
INV_X4 _13042_ ( .A(_05318_ ), .ZN(_05319_ ) );
NAND3_X2 _13043_ ( .A1(_04381_ ), .A2(_05143_ ), .A3(_04405_ ), .ZN(_05320_ ) );
NAND2_X1 _13044_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [19] ), .ZN(_05321_ ) );
AND2_X4 _13045_ ( .A1(_05320_ ), .A2(_05321_ ), .ZN(_05322_ ) );
XNOR2_X2 _13046_ ( .A(_05322_ ), .B(_04380_ ), .ZN(_05323_ ) );
INV_X4 _13047_ ( .A(_05323_ ), .ZN(_05324_ ) );
NAND2_X1 _13048_ ( .A1(_05319_ ), .A2(_05324_ ), .ZN(_05325_ ) );
OR3_X2 _13049_ ( .A1(_05310_ ), .A2(_05314_ ), .A3(_05325_ ), .ZN(_05326_ ) );
OR4_X4 _13050_ ( .A1(_05285_ ), .A2(_05289_ ), .A3(_05293_ ), .A4(_05326_ ), .ZN(_05327_ ) );
NOR2_X1 _13051_ ( .A1(_05308_ ), .A2(_05309_ ), .ZN(_05328_ ) );
INV_X1 _13052_ ( .A(_05328_ ), .ZN(_05329_ ) );
NAND3_X1 _13053_ ( .A1(_05329_ ), .A2(_02535_ ), .A3(_05296_ ), .ZN(_05330_ ) );
INV_X1 _13054_ ( .A(_02610_ ), .ZN(_05331_ ) );
INV_X1 _13055_ ( .A(_05313_ ), .ZN(_05332_ ) );
NOR3_X1 _13056_ ( .A1(_05302_ ), .A2(_05331_ ), .A3(_05332_ ), .ZN(_05333_ ) );
AOI21_X1 _13057_ ( .A(_05333_ ), .B1(_04505_ ), .B2(_05301_ ), .ZN(_05334_ ) );
NOR3_X1 _13058_ ( .A1(_05334_ ), .A2(_05328_ ), .A3(_05297_ ), .ZN(_05335_ ) );
OR2_X1 _13059_ ( .A1(_05310_ ), .A2(_05314_ ), .ZN(_05336_ ) );
INV_X1 _13060_ ( .A(_02684_ ), .ZN(_05337_ ) );
AND2_X1 _13061_ ( .A1(_05288_ ), .A2(_05337_ ), .ZN(_05338_ ) );
NOR2_X1 _13062_ ( .A1(_05288_ ), .A2(_05337_ ), .ZN(_05339_ ) );
OAI211_X1 _13063_ ( .A(_02709_ ), .B(_05292_ ), .C1(_05338_ ), .C2(_05339_ ), .ZN(_05340_ ) );
NAND4_X1 _13064_ ( .A1(_05286_ ), .A2(_02683_ ), .A3(_02663_ ), .A4(_05287_ ), .ZN(_05341_ ) );
AOI21_X1 _13065_ ( .A(_05325_ ), .B1(_05340_ ), .B2(_05341_ ), .ZN(_05342_ ) );
AOI21_X1 _13066_ ( .A(_05342_ ), .B1(_04380_ ), .B2(_05322_ ), .ZN(_05343_ ) );
NAND3_X1 _13067_ ( .A1(_05324_ ), .A2(_02635_ ), .A3(_05317_ ), .ZN(_05344_ ) );
AOI21_X1 _13068_ ( .A(_05336_ ), .B1(_05343_ ), .B2(_05344_ ), .ZN(_05345_ ) );
AOI211_X1 _13069_ ( .A(_05335_ ), .B(_05345_ ), .C1(_02561_ ), .C2(_05306_ ), .ZN(_05346_ ) );
NAND3_X1 _13070_ ( .A1(_05327_ ), .A2(_05330_ ), .A3(_05346_ ), .ZN(_05347_ ) );
OR2_X1 _13071_ ( .A1(_04700_ ), .A2(\ID_EX_typ [4] ), .ZN(_05348_ ) );
NAND2_X1 _13072_ ( .A1(_03208_ ), .A2(\ID_EX_typ [4] ), .ZN(_05349_ ) );
NAND2_X1 _13073_ ( .A1(_05348_ ), .A2(_05349_ ), .ZN(_05350_ ) );
INV_X1 _13074_ ( .A(_03207_ ), .ZN(_05351_ ) );
NOR2_X1 _13075_ ( .A1(_05350_ ), .A2(_05351_ ), .ZN(_05352_ ) );
AOI21_X1 _13076_ ( .A(_03207_ ), .B1(_05348_ ), .B2(_05349_ ), .ZN(_05353_ ) );
NOR2_X1 _13077_ ( .A1(_05352_ ), .A2(_05353_ ), .ZN(_05354_ ) );
NAND3_X1 _13078_ ( .A1(_04703_ ), .A2(_05144_ ), .A3(_04721_ ), .ZN(_05355_ ) );
NAND2_X1 _13079_ ( .A1(_02488_ ), .A2(\ID_EX_typ [4] ), .ZN(_05356_ ) );
NAND2_X1 _13080_ ( .A1(_05355_ ), .A2(_05356_ ), .ZN(_05357_ ) );
XNOR2_X1 _13081_ ( .A(_05357_ ), .B(_02487_ ), .ZN(_05358_ ) );
NOR2_X1 _13082_ ( .A1(_05354_ ), .A2(_05358_ ), .ZN(_05359_ ) );
OR2_X1 _13083_ ( .A1(_04653_ ), .A2(\ID_EX_typ [4] ), .ZN(_05360_ ) );
NAND2_X1 _13084_ ( .A1(_02511_ ), .A2(\ID_EX_typ [4] ), .ZN(_05361_ ) );
NAND2_X1 _13085_ ( .A1(_05360_ ), .A2(_05361_ ), .ZN(_05362_ ) );
INV_X1 _13086_ ( .A(_02510_ ), .ZN(_05363_ ) );
NOR2_X1 _13087_ ( .A1(_05362_ ), .A2(_05363_ ), .ZN(_05364_ ) );
AOI21_X1 _13088_ ( .A(_02510_ ), .B1(_05360_ ), .B2(_05361_ ), .ZN(_05365_ ) );
NOR2_X1 _13089_ ( .A1(_05364_ ), .A2(_05365_ ), .ZN(_05366_ ) );
INV_X1 _13090_ ( .A(_05366_ ), .ZN(_05367_ ) );
NAND3_X1 _13091_ ( .A1(_04656_ ), .A2(_05144_ ), .A3(_04675_ ), .ZN(_05368_ ) );
NAND2_X1 _13092_ ( .A1(_03210_ ), .A2(\ID_EX_typ [4] ), .ZN(_05369_ ) );
NAND2_X1 _13093_ ( .A1(_05368_ ), .A2(_05369_ ), .ZN(_05370_ ) );
XNOR2_X1 _13094_ ( .A(_03184_ ), .B(_05370_ ), .ZN(_05371_ ) );
INV_X1 _13095_ ( .A(_05371_ ), .ZN(_05372_ ) );
AND3_X1 _13096_ ( .A1(_05359_ ), .A2(_05367_ ), .A3(_05372_ ), .ZN(_05373_ ) );
NAND2_X1 _13097_ ( .A1(_05347_ ), .A2(_05373_ ), .ZN(_05374_ ) );
AND3_X1 _13098_ ( .A1(_05372_ ), .A2(_02510_ ), .A3(_05362_ ), .ZN(_05375_ ) );
AOI22_X1 _13099_ ( .A1(_03163_ ), .A2(_03183_ ), .B1(_05368_ ), .B2(_05369_ ), .ZN(_05376_ ) );
OAI21_X1 _13100_ ( .A(_05359_ ), .B1(_05375_ ), .B2(_05376_ ), .ZN(_05377_ ) );
INV_X1 _13101_ ( .A(_05358_ ), .ZN(_05378_ ) );
NAND3_X1 _13102_ ( .A1(_05378_ ), .A2(_03207_ ), .A3(_05350_ ), .ZN(_05379_ ) );
NAND2_X1 _13103_ ( .A1(_05357_ ), .A2(_02487_ ), .ZN(_05380_ ) );
AND3_X1 _13104_ ( .A1(_05377_ ), .A2(_05379_ ), .A3(_05380_ ), .ZN(_05381_ ) );
AOI21_X1 _13105_ ( .A(_05162_ ), .B1(_05374_ ), .B2(_05381_ ), .ZN(_05382_ ) );
INV_X1 _13106_ ( .A(_05382_ ), .ZN(_05383_ ) );
AOI21_X1 _13107_ ( .A(_05147_ ), .B1(_02399_ ), .B2(_02400_ ), .ZN(_05384_ ) );
AND2_X1 _13108_ ( .A1(_05139_ ), .A2(_05384_ ), .ZN(_05385_ ) );
INV_X1 _13109_ ( .A(_05135_ ), .ZN(_05386_ ) );
AOI22_X1 _13110_ ( .A1(_05157_ ), .A2(_05158_ ), .B1(_02447_ ), .B2(_02428_ ), .ZN(_05387_ ) );
OAI21_X1 _13111_ ( .A(_05387_ ), .B1(_05154_ ), .B2(_05155_ ), .ZN(_05388_ ) );
INV_X1 _13112_ ( .A(_02425_ ), .ZN(_05389_ ) );
OAI21_X1 _13113_ ( .A(_05388_ ), .B1(_05389_ ), .B2(_05153_ ), .ZN(_05390_ ) );
AOI221_X4 _13114_ ( .A(_05385_ ), .B1(_05136_ ), .B2(_05386_ ), .C1(_05149_ ), .C2(_05390_ ), .ZN(_05391_ ) );
AND2_X2 _13115_ ( .A1(_05383_ ), .A2(_05391_ ), .ZN(_05392_ ) );
MUX2_X1 _13116_ ( .A(_05130_ ), .B(_05131_ ), .S(_05392_ ), .Z(_05393_ ) );
AND3_X1 _13117_ ( .A1(_05020_ ), .A2(_02884_ ), .A3(_02864_ ), .ZN(_05394_ ) );
INV_X1 _13118_ ( .A(_05394_ ), .ZN(_05395_ ) );
INV_X1 _13119_ ( .A(_02910_ ), .ZN(_05396_ ) );
AOI21_X1 _13120_ ( .A(_05119_ ), .B1(_02835_ ), .B2(_05113_ ), .ZN(_05397_ ) );
INV_X1 _13121_ ( .A(_05022_ ), .ZN(_05398_ ) );
OAI221_X1 _13122_ ( .A(_05395_ ), .B1(_05396_ ), .B2(_04951_ ), .C1(_05397_ ), .C2(_05398_ ), .ZN(_05399_ ) );
NAND3_X1 _13123_ ( .A1(_02908_ ), .A2(_02909_ ), .A3(_04951_ ), .ZN(_05400_ ) );
AND2_X1 _13124_ ( .A1(_04999_ ), .A2(_05092_ ), .ZN(_05401_ ) );
NAND4_X1 _13125_ ( .A1(_05399_ ), .A2(_05071_ ), .A3(_05400_ ), .A4(_05401_ ), .ZN(_05402_ ) );
AND3_X1 _13126_ ( .A1(_05047_ ), .A2(_02788_ ), .A3(_05069_ ), .ZN(_05403_ ) );
AND3_X1 _13127_ ( .A1(_04998_ ), .A2(_02734_ ), .A3(_02713_ ), .ZN(_05404_ ) );
NAND2_X1 _13128_ ( .A1(_05092_ ), .A2(_05404_ ), .ZN(_05405_ ) );
OAI21_X1 _13129_ ( .A(_05405_ ), .B1(_05213_ ), .B2(_05091_ ), .ZN(_05406_ ) );
AOI221_X4 _13130_ ( .A(_05403_ ), .B1(_02812_ ), .B2(_05045_ ), .C1(_05406_ ), .C2(_05071_ ), .ZN(_05407_ ) );
AND2_X1 _13131_ ( .A1(_05402_ ), .A2(_05407_ ), .ZN(_05408_ ) );
OR2_X1 _13132_ ( .A1(_05408_ ), .A2(_04930_ ), .ZN(_05409_ ) );
NAND3_X1 _13133_ ( .A1(_04779_ ), .A2(_03020_ ), .A3(_04752_ ), .ZN(_05410_ ) );
INV_X1 _13134_ ( .A(_02996_ ), .ZN(_05411_ ) );
INV_X1 _13135_ ( .A(_04829_ ), .ZN(_05412_ ) );
NAND3_X1 _13136_ ( .A1(_04855_ ), .A2(_03095_ ), .A3(_04876_ ), .ZN(_05413_ ) );
OAI21_X1 _13137_ ( .A(_05413_ ), .B1(_05187_ ), .B2(_04853_ ), .ZN(_05414_ ) );
INV_X1 _13138_ ( .A(_04925_ ), .ZN(_05415_ ) );
NAND2_X1 _13139_ ( .A1(_03045_ ), .A2(_04900_ ), .ZN(_05416_ ) );
AOI21_X1 _13140_ ( .A(_04926_ ), .B1(_05415_ ), .B2(_05416_ ), .ZN(_05417_ ) );
AOI21_X1 _13141_ ( .A(_05414_ ), .B1(_04879_ ), .B2(_05417_ ), .ZN(_05418_ ) );
OAI221_X1 _13142_ ( .A(_05410_ ), .B1(_05411_ ), .B2(_04778_ ), .C1(_05412_ ), .C2(_05418_ ), .ZN(_05419_ ) );
AND2_X1 _13143_ ( .A1(_02948_ ), .A2(_04827_ ), .ZN(_05420_ ) );
AND2_X1 _13144_ ( .A1(_04806_ ), .A2(_05420_ ), .ZN(_05421_ ) );
AOI21_X1 _13145_ ( .A(_05421_ ), .B1(_04781_ ), .B2(_04804_ ), .ZN(_05422_ ) );
INV_X1 _13146_ ( .A(_05422_ ), .ZN(_05423_ ) );
AOI21_X1 _13147_ ( .A(_05419_ ), .B1(_04780_ ), .B2(_05423_ ), .ZN(_05424_ ) );
AND2_X1 _13148_ ( .A1(_05409_ ), .A2(_05424_ ), .ZN(_05425_ ) );
INV_X1 _13149_ ( .A(_04727_ ), .ZN(_05426_ ) );
OR2_X1 _13150_ ( .A1(_05425_ ), .A2(_05426_ ), .ZN(_05427_ ) );
NAND2_X1 _13151_ ( .A1(_02709_ ), .A2(_04352_ ), .ZN(_05428_ ) );
NOR3_X1 _13152_ ( .A1(_04376_ ), .A2(_04377_ ), .A3(_05428_ ), .ZN(_05429_ ) );
OAI211_X1 _13153_ ( .A(_04431_ ), .B(_04408_ ), .C1(_05429_ ), .C2(_04376_ ), .ZN(_05430_ ) );
AND3_X1 _13154_ ( .A1(_04406_ ), .A2(_02658_ ), .A3(_02638_ ), .ZN(_05431_ ) );
INV_X1 _13155_ ( .A(_05431_ ), .ZN(_05432_ ) );
NAND3_X1 _13156_ ( .A1(_04408_ ), .A2(_02635_ ), .A3(_04429_ ), .ZN(_05433_ ) );
AND3_X1 _13157_ ( .A1(_05430_ ), .A2(_05432_ ), .A3(_05433_ ), .ZN(_05434_ ) );
NOR2_X1 _13158_ ( .A1(_05434_ ), .A2(_04530_ ), .ZN(_05435_ ) );
AND2_X1 _13159_ ( .A1(_02535_ ), .A2(_04454_ ), .ZN(_05436_ ) );
NAND2_X1 _13160_ ( .A1(_04481_ ), .A2(_05436_ ), .ZN(_05437_ ) );
OAI21_X1 _13161_ ( .A(_05437_ ), .B1(_05307_ ), .B2(_04480_ ), .ZN(_05438_ ) );
INV_X1 _13162_ ( .A(_04482_ ), .ZN(_05439_ ) );
AOI21_X1 _13163_ ( .A(_04527_ ), .B1(_02610_ ), .B2(_04503_ ), .ZN(_05440_ ) );
NOR3_X1 _13164_ ( .A1(_05439_ ), .A2(_04528_ ), .A3(_05440_ ), .ZN(_05441_ ) );
NOR3_X1 _13165_ ( .A1(_05435_ ), .A2(_05438_ ), .A3(_05441_ ), .ZN(_05442_ ) );
INV_X1 _13166_ ( .A(_04726_ ), .ZN(_05443_ ) );
NOR2_X1 _13167_ ( .A1(_05442_ ), .A2(_05443_ ), .ZN(_05444_ ) );
INV_X1 _13168_ ( .A(_04559_ ), .ZN(_05445_ ) );
AOI21_X1 _13169_ ( .A(_04583_ ), .B1(_02448_ ), .B2(_05445_ ), .ZN(_05446_ ) );
NOR2_X1 _13170_ ( .A1(_05446_ ), .A2(_04582_ ), .ZN(_05447_ ) );
AND3_X1 _13171_ ( .A1(_04607_ ), .A2(_04630_ ), .A3(_05447_ ), .ZN(_05448_ ) );
OR2_X1 _13172_ ( .A1(_05136_ ), .A2(_04629_ ), .ZN(_05449_ ) );
NOR2_X1 _13173_ ( .A1(_02401_ ), .A2(_04605_ ), .ZN(_05450_ ) );
NAND2_X1 _13174_ ( .A1(_04630_ ), .A2(_05450_ ), .ZN(_05451_ ) );
INV_X1 _13175_ ( .A(_04631_ ), .ZN(_05452_ ) );
NOR2_X1 _13176_ ( .A1(_05351_ ), .A2(_04700_ ), .ZN(_05453_ ) );
NAND2_X1 _13177_ ( .A1(_05453_ ), .A2(_04723_ ), .ZN(_05454_ ) );
INV_X1 _13178_ ( .A(_02487_ ), .ZN(_05455_ ) );
OAI21_X1 _13179_ ( .A(_05454_ ), .B1(_05455_ ), .B2(_04722_ ), .ZN(_05456_ ) );
AOI21_X1 _13180_ ( .A(_04676_ ), .B1(_03163_ ), .B2(_03183_ ), .ZN(_05457_ ) );
NOR2_X1 _13181_ ( .A1(_05363_ ), .A2(_04653_ ), .ZN(_05458_ ) );
AOI21_X1 _13182_ ( .A(_05457_ ), .B1(_04677_ ), .B2(_05458_ ), .ZN(_05459_ ) );
INV_X1 _13183_ ( .A(_05459_ ), .ZN(_05460_ ) );
AOI21_X1 _13184_ ( .A(_05456_ ), .B1(_05460_ ), .B2(_04724_ ), .ZN(_05461_ ) );
OAI211_X1 _13185_ ( .A(_05449_ ), .B(_05451_ ), .C1(_05452_ ), .C2(_05461_ ), .ZN(_05462_ ) );
NOR3_X1 _13186_ ( .A1(_05444_ ), .A2(_05448_ ), .A3(_05462_ ), .ZN(_05463_ ) );
AND2_X2 _13187_ ( .A1(_05123_ ), .A2(\ID_EX_typ [2] ), .ZN(_05464_ ) );
AND3_X1 _13188_ ( .A1(_05427_ ), .A2(_05463_ ), .A3(_05464_ ), .ZN(_05465_ ) );
AND2_X1 _13189_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_7 ), .ZN(_05466_ ) );
AND2_X2 _13190_ ( .A1(_05466_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05467_ ) );
INV_X1 _13191_ ( .A(_05467_ ), .ZN(_05468_ ) );
AOI21_X1 _13192_ ( .A(_05468_ ), .B1(_05427_ ), .B2(_05463_ ), .ZN(_05469_ ) );
NOR3_X1 _13193_ ( .A1(_05465_ ), .A2(_05469_ ), .A3(_05124_ ), .ZN(_05470_ ) );
AOI221_X4 _13194_ ( .A(_04292_ ), .B1(_05122_ ), .B2(_05124_ ), .C1(_05393_ ), .C2(_05470_ ), .ZN(_05471_ ) );
INV_X1 _13195_ ( .A(_04292_ ), .ZN(_05472_ ) );
AOI21_X1 _13196_ ( .A(_05472_ ), .B1(_04727_ ), .B2(_05121_ ), .ZN(_05473_ ) );
NOR2_X4 _13197_ ( .A1(_05471_ ), .A2(_05473_ ), .ZN(_05474_ ) );
BUF_X8 _13198_ ( .A(_05474_ ), .Z(_05475_ ) );
MUX2_X1 _13199_ ( .A(_04179_ ), .B(_04290_ ), .S(_05475_ ), .Z(_05476_ ) );
OR2_X2 _13200_ ( .A1(_05476_ ), .A2(\ID_EX_typ [3] ), .ZN(_05477_ ) );
INV_X1 _13201_ ( .A(_04145_ ), .ZN(_05478_ ) );
BUF_X4 _13202_ ( .A(_05478_ ), .Z(_05479_ ) );
BUF_X4 _13203_ ( .A(_05479_ ), .Z(_05480_ ) );
INV_X2 _13204_ ( .A(\ID_EX_typ [3] ), .ZN(_05481_ ) );
BUF_X4 _13205_ ( .A(_05481_ ), .Z(_05482_ ) );
BUF_X4 _13206_ ( .A(_05482_ ), .Z(_05483_ ) );
INV_X1 _13207_ ( .A(\ID_EX_csr [10] ), .ZN(_05484_ ) );
INV_X1 _13208_ ( .A(\ID_EX_csr [5] ), .ZN(_05485_ ) );
INV_X1 _13209_ ( .A(\ID_EX_csr [4] ), .ZN(_05486_ ) );
INV_X1 _13210_ ( .A(\ID_EX_csr [11] ), .ZN(_05487_ ) );
NAND4_X1 _13211_ ( .A1(_05484_ ), .A2(_05485_ ), .A3(_05486_ ), .A4(_05487_ ), .ZN(_05488_ ) );
AND2_X1 _13212_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_05489_ ) );
INV_X1 _13213_ ( .A(_05489_ ), .ZN(_05490_ ) );
NOR2_X1 _13214_ ( .A1(_05488_ ), .A2(_05490_ ), .ZN(_05491_ ) );
INV_X1 _13215_ ( .A(\ID_EX_csr [7] ), .ZN(_05492_ ) );
AND3_X1 _13216_ ( .A1(_05491_ ), .A2(_05492_ ), .A3(\ID_EX_csr [6] ), .ZN(_05493_ ) );
BUF_X4 _13217_ ( .A(_05493_ ), .Z(_05494_ ) );
INV_X1 _13218_ ( .A(\ID_EX_csr [0] ), .ZN(_05495_ ) );
NOR2_X1 _13219_ ( .A1(_05495_ ), .A2(\ID_EX_csr [1] ), .ZN(_05496_ ) );
NOR2_X1 _13220_ ( .A1(\ID_EX_csr [3] ), .A2(\ID_EX_csr [2] ), .ZN(_05497_ ) );
AND2_X2 _13221_ ( .A1(_05496_ ), .A2(_05497_ ), .ZN(_05498_ ) );
NAND3_X1 _13222_ ( .A1(_05494_ ), .A2(\mepc [30] ), .A3(_05498_ ), .ZN(_05499_ ) );
BUF_X4 _13223_ ( .A(_05491_ ), .Z(_05500_ ) );
NOR2_X1 _13224_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_05501_ ) );
BUF_X4 _13225_ ( .A(_05501_ ), .Z(_05502_ ) );
INV_X1 _13226_ ( .A(\ID_EX_csr [1] ), .ZN(_05503_ ) );
AND3_X1 _13227_ ( .A1(_05497_ ), .A2(_05503_ ), .A3(_05495_ ), .ZN(_05504_ ) );
BUF_X4 _13228_ ( .A(_05504_ ), .Z(_05505_ ) );
NAND4_X1 _13229_ ( .A1(_05500_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_05502_ ), .A4(_05505_ ), .ZN(_05506_ ) );
AND2_X1 _13230_ ( .A1(_05499_ ), .A2(_05506_ ), .ZN(_05507_ ) );
BUF_X4 _13231_ ( .A(_05500_ ), .Z(_05508_ ) );
INV_X1 _13232_ ( .A(\ID_EX_csr [3] ), .ZN(_05509_ ) );
AND3_X1 _13233_ ( .A1(_05496_ ), .A2(_05509_ ), .A3(\ID_EX_csr [2] ), .ZN(_05510_ ) );
BUF_X2 _13234_ ( .A(_05510_ ), .Z(_05511_ ) );
BUF_X4 _13235_ ( .A(_05502_ ), .Z(_05512_ ) );
NAND4_X1 _13236_ ( .A1(_05508_ ), .A2(_05511_ ), .A3(\mtvec [30] ), .A4(_05512_ ), .ZN(_05513_ ) );
AND4_X1 _13237_ ( .A1(\ID_EX_csr [10] ), .A2(_05485_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_05514_ ) );
AND3_X1 _13238_ ( .A1(_05514_ ), .A2(_05501_ ), .A3(_05489_ ), .ZN(_05515_ ) );
NAND2_X1 _13239_ ( .A1(_05515_ ), .A2(_05498_ ), .ZN(_05516_ ) );
BUF_X2 _13240_ ( .A(_05516_ ), .Z(_05517_ ) );
BUF_X4 _13241_ ( .A(_05493_ ), .Z(_05518_ ) );
INV_X1 _13242_ ( .A(\ID_EX_csr [2] ), .ZN(_05519_ ) );
NAND3_X1 _13243_ ( .A1(_05509_ ), .A2(_05519_ ), .A3(\ID_EX_csr [1] ), .ZN(_05520_ ) );
NOR2_X2 _13244_ ( .A1(_05520_ ), .A2(\ID_EX_csr [0] ), .ZN(_05521_ ) );
NAND3_X1 _13245_ ( .A1(_05518_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_05521_ ), .ZN(_05522_ ) );
NAND4_X1 _13246_ ( .A1(_05507_ ), .A2(_05513_ ), .A3(_05517_ ), .A4(_05522_ ), .ZN(_05523_ ) );
XNOR2_X1 _13247_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_05524_ ) );
XNOR2_X1 _13248_ ( .A(fanout_net_6 ), .B(\ID_EX_csr [0] ), .ZN(_05525_ ) );
XNOR2_X1 _13249_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .ZN(_05526_ ) );
XNOR2_X1 _13250_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_05527_ ) );
AND4_X1 _13251_ ( .A1(_05524_ ), .A2(_05525_ ), .A3(_05526_ ), .A4(_05527_ ), .ZN(_05528_ ) );
XNOR2_X1 _13252_ ( .A(\EX_LS_dest_csreg_mem [1] ), .B(\ID_EX_csr [1] ), .ZN(_05529_ ) );
XNOR2_X1 _13253_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_05530_ ) );
AND4_X2 _13254_ ( .A1(_04104_ ), .A2(_05528_ ), .A3(_05529_ ), .A4(_05530_ ), .ZN(_05531_ ) );
INV_X1 _13255_ ( .A(\ID_EX_csr [9] ), .ZN(_05532_ ) );
INV_X1 _13256_ ( .A(\ID_EX_csr [8] ), .ZN(_05533_ ) );
AOI22_X1 _13257_ ( .A1(\EX_LS_dest_csreg_mem [9] ), .A2(_05532_ ), .B1(_05533_ ), .B2(\EX_LS_dest_csreg_mem [8] ), .ZN(_05534_ ) );
XNOR2_X1 _13258_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_05535_ ) );
XNOR2_X1 _13259_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_05536_ ) );
INV_X1 _13260_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_05537_ ) );
INV_X1 _13261_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_05538_ ) );
AOI22_X1 _13262_ ( .A1(_05537_ ), .A2(\ID_EX_csr [9] ), .B1(_05538_ ), .B2(\ID_EX_csr [8] ), .ZN(_05539_ ) );
AND4_X1 _13263_ ( .A1(_05534_ ), .A2(_05535_ ), .A3(_05536_ ), .A4(_05539_ ), .ZN(_05540_ ) );
XNOR2_X1 _13264_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_05541_ ) );
XNOR2_X1 _13265_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_05542_ ) );
AND3_X2 _13266_ ( .A1(_05540_ ), .A2(_05541_ ), .A3(_05542_ ), .ZN(_05543_ ) );
AND2_X1 _13267_ ( .A1(_05531_ ), .A2(_05543_ ), .ZN(_05544_ ) );
BUF_X4 _13268_ ( .A(_05544_ ), .Z(_05545_ ) );
INV_X1 _13269_ ( .A(_05545_ ), .ZN(_05546_ ) );
NAND2_X1 _13270_ ( .A1(_05523_ ), .A2(_05546_ ), .ZN(_05547_ ) );
NAND3_X1 _13271_ ( .A1(_05531_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_05543_ ), .ZN(_05548_ ) );
AND2_X1 _13272_ ( .A1(_05547_ ), .A2(_05548_ ), .ZN(_05549_ ) );
INV_X1 _13273_ ( .A(_05549_ ), .ZN(_05550_ ) );
OAI211_X1 _13274_ ( .A(_05477_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05550_ ), .ZN(_05551_ ) );
CLKBUF_X2 _13275_ ( .A(_04145_ ), .Z(_05552_ ) );
BUF_X4 _13276_ ( .A(_05552_ ), .Z(_05553_ ) );
OAI21_X1 _13277_ ( .A(fanout_net_7 ), .B1(_03249_ ), .B2(_03221_ ), .ZN(_05554_ ) );
OAI211_X1 _13278_ ( .A(_05553_ ), .B(_05554_ ), .C1(_04290_ ), .C2(fanout_net_7 ), .ZN(_05555_ ) );
AOI21_X1 _13279_ ( .A(_04159_ ), .B1(_05551_ ), .B2(_05555_ ), .ZN(_00158_ ) );
BUF_X4 _13280_ ( .A(_05481_ ), .Z(_05556_ ) );
NAND4_X1 _13281_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_05557_ ) );
NAND2_X1 _13282_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_05558_ ) );
INV_X1 _13283_ ( .A(\ID_EX_pc [13] ), .ZN(_05559_ ) );
INV_X1 _13284_ ( .A(\ID_EX_pc [12] ), .ZN(_05560_ ) );
NOR4_X1 _13285_ ( .A1(_05557_ ), .A2(_05558_ ), .A3(_05559_ ), .A4(_05560_ ), .ZN(_05561_ ) );
AND2_X1 _13286_ ( .A1(_04166_ ), .A2(_05561_ ), .ZN(_05562_ ) );
AND4_X1 _13287_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_05563_ ) );
AND2_X1 _13288_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_05564_ ) );
AND4_X1 _13289_ ( .A1(\ID_EX_pc [21] ), .A2(_05563_ ), .A3(\ID_EX_pc [20] ), .A4(_05564_ ), .ZN(_05565_ ) );
NAND2_X1 _13290_ ( .A1(_05562_ ), .A2(_05565_ ), .ZN(_05566_ ) );
INV_X1 _13291_ ( .A(\ID_EX_pc [27] ), .ZN(_05567_ ) );
INV_X1 _13292_ ( .A(\ID_EX_pc [26] ), .ZN(_05568_ ) );
NOR3_X1 _13293_ ( .A1(_05566_ ), .A2(_05567_ ), .A3(_05568_ ), .ZN(_05569_ ) );
NAND2_X1 _13294_ ( .A1(_05569_ ), .A2(\ID_EX_pc [28] ), .ZN(_05570_ ) );
XNOR2_X1 _13295_ ( .A(_05570_ ), .B(\ID_EX_pc [29] ), .ZN(_05571_ ) );
OAI21_X1 _13296_ ( .A(_05571_ ), .B1(_05471_ ), .B2(_05473_ ), .ZN(_05572_ ) );
INV_X4 _13297_ ( .A(_05474_ ), .ZN(_05573_ ) );
BUF_X4 _13298_ ( .A(_05573_ ), .Z(_05574_ ) );
NAND2_X1 _13299_ ( .A1(_04283_ ), .A2(_04284_ ), .ZN(_05575_ ) );
XOR2_X1 _13300_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .Z(_05576_ ) );
XNOR2_X1 _13301_ ( .A(_05575_ ), .B(_05576_ ), .ZN(_05577_ ) );
OAI211_X1 _13302_ ( .A(_05556_ ), .B(_05572_ ), .C1(_05574_ ), .C2(_05577_ ), .ZN(_05578_ ) );
BUF_X4 _13303_ ( .A(_05531_ ), .Z(_05579_ ) );
BUF_X4 _13304_ ( .A(_05543_ ), .Z(_05580_ ) );
NAND3_X1 _13305_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [29] ), .A3(_05580_ ), .ZN(_05581_ ) );
BUF_X4 _13306_ ( .A(_05494_ ), .Z(_05582_ ) );
BUF_X4 _13307_ ( .A(_05498_ ), .Z(_05583_ ) );
NAND3_X1 _13308_ ( .A1(_05582_ ), .A2(\mepc [29] ), .A3(_05583_ ), .ZN(_05584_ ) );
BUF_X4 _13309_ ( .A(_05500_ ), .Z(_05585_ ) );
BUF_X4 _13310_ ( .A(_05511_ ), .Z(_05586_ ) );
BUF_X4 _13311_ ( .A(_05502_ ), .Z(_05587_ ) );
NAND4_X1 _13312_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(\mtvec [29] ), .A4(_05587_ ), .ZN(_05588_ ) );
BUF_X4 _13313_ ( .A(_05505_ ), .Z(_05589_ ) );
NAND4_X1 _13314_ ( .A1(_05585_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_05587_ ), .A4(_05589_ ), .ZN(_05590_ ) );
AND3_X1 _13315_ ( .A1(_05584_ ), .A2(_05588_ ), .A3(_05590_ ), .ZN(_05591_ ) );
BUF_X4 _13316_ ( .A(_05518_ ), .Z(_05592_ ) );
BUF_X4 _13317_ ( .A(_05521_ ), .Z(_05593_ ) );
BUF_X2 _13318_ ( .A(_05593_ ), .Z(_05594_ ) );
NAND3_X1 _13319_ ( .A1(_05592_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_05594_ ), .ZN(_05595_ ) );
AND3_X1 _13320_ ( .A1(_05591_ ), .A2(_05517_ ), .A3(_05595_ ), .ZN(_05596_ ) );
OAI21_X1 _13321_ ( .A(_05581_ ), .B1(_05596_ ), .B2(_05545_ ), .ZN(_05597_ ) );
OAI211_X1 _13322_ ( .A(_05578_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05597_ ), .ZN(_05598_ ) );
MUX2_X1 _13323_ ( .A(_05577_ ), .B(_03287_ ), .S(fanout_net_7 ), .Z(_05599_ ) );
BUF_X4 _13324_ ( .A(_05478_ ), .Z(_05600_ ) );
BUF_X2 _13325_ ( .A(_05600_ ), .Z(_05601_ ) );
OR2_X2 _13326_ ( .A1(_05599_ ), .A2(_05601_ ), .ZN(_05602_ ) );
AOI21_X1 _13327_ ( .A(_04159_ ), .B1(_05598_ ), .B2(_05602_ ), .ZN(_00159_ ) );
NAND3_X1 _13328_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_05580_ ), .ZN(_05603_ ) );
BUF_X4 _13329_ ( .A(_05494_ ), .Z(_05604_ ) );
BUF_X4 _13330_ ( .A(_05498_ ), .Z(_05605_ ) );
NAND3_X1 _13331_ ( .A1(_05604_ ), .A2(\mepc [20] ), .A3(_05605_ ), .ZN(_05606_ ) );
NAND2_X1 _13332_ ( .A1(_05515_ ), .A2(_05521_ ), .ZN(_05607_ ) );
AND2_X2 _13333_ ( .A1(_05516_ ), .A2(_05607_ ), .ZN(_05608_ ) );
NAND3_X1 _13334_ ( .A1(_05582_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_05593_ ), .ZN(_05609_ ) );
NAND4_X1 _13335_ ( .A1(_05500_ ), .A2(_05511_ ), .A3(\mtvec [20] ), .A4(_05502_ ), .ZN(_05610_ ) );
NAND4_X1 _13336_ ( .A1(_05500_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_05502_ ), .A4(_05505_ ), .ZN(_05611_ ) );
AND2_X1 _13337_ ( .A1(_05610_ ), .A2(_05611_ ), .ZN(_05612_ ) );
AND4_X1 _13338_ ( .A1(_05606_ ), .A2(_05608_ ), .A3(_05609_ ), .A4(_05612_ ), .ZN(_05613_ ) );
OAI21_X1 _13339_ ( .A(_05603_ ), .B1(_05613_ ), .B2(_05545_ ), .ZN(_05614_ ) );
NAND3_X1 _13340_ ( .A1(_04166_ ), .A2(_05561_ ), .A3(_05564_ ), .ZN(_05615_ ) );
XNOR2_X1 _13341_ ( .A(_05615_ ), .B(\ID_EX_pc [20] ), .ZN(_05616_ ) );
XOR2_X1 _13342_ ( .A(_04255_ ), .B(_04260_ ), .Z(_05617_ ) );
MUX2_X1 _13343_ ( .A(_05616_ ), .B(_05617_ ), .S(_05475_ ), .Z(_05618_ ) );
MUX2_X2 _13344_ ( .A(_05614_ ), .B(_05618_ ), .S(_05482_ ), .Z(_05619_ ) );
BUF_X4 _13345_ ( .A(_05479_ ), .Z(_05620_ ) );
NAND2_X1 _13346_ ( .A1(_05619_ ), .A2(_05620_ ), .ZN(_05621_ ) );
AND2_X2 _13347_ ( .A1(_04145_ ), .A2(fanout_net_7 ), .ZN(_05622_ ) );
AND3_X1 _13348_ ( .A1(_03255_ ), .A2(_03252_ ), .A3(_05622_ ), .ZN(_05623_ ) );
BUF_X4 _13349_ ( .A(_04147_ ), .Z(_05624_ ) );
AOI21_X1 _13350_ ( .A(_05623_ ), .B1(_05624_ ), .B2(_05617_ ), .ZN(_05625_ ) );
AOI21_X1 _13351_ ( .A(_04159_ ), .B1(_05621_ ), .B2(_05625_ ), .ZN(_00160_ ) );
BUF_X8 _13352_ ( .A(_05474_ ), .Z(_05626_ ) );
INV_X1 _13353_ ( .A(_04241_ ), .ZN(_05627_ ) );
OAI21_X1 _13354_ ( .A(_04245_ ), .B1(_04230_ ), .B2(_04238_ ), .ZN(_05628_ ) );
AOI21_X1 _13355_ ( .A(_05627_ ), .B1(_05628_ ), .B2(_04252_ ), .ZN(_05629_ ) );
NOR2_X1 _13356_ ( .A1(_05629_ ), .A2(_04247_ ), .ZN(_05630_ ) );
XNOR2_X1 _13357_ ( .A(_05630_ ), .B(_04240_ ), .ZN(_05631_ ) );
AOI21_X1 _13358_ ( .A(\ID_EX_typ [3] ), .B1(_05626_ ), .B2(_05631_ ), .ZN(_05632_ ) );
BUF_X8 _13359_ ( .A(_05626_ ), .Z(_05633_ ) );
NAND3_X1 _13360_ ( .A1(_04166_ ), .A2(\ID_EX_pc [18] ), .A3(_05561_ ), .ZN(_05634_ ) );
INV_X1 _13361_ ( .A(\ID_EX_pc [19] ), .ZN(_05635_ ) );
XNOR2_X1 _13362_ ( .A(_05634_ ), .B(_05635_ ), .ZN(_05636_ ) );
OAI21_X1 _13363_ ( .A(_05632_ ), .B1(_05633_ ), .B2(_05636_ ), .ZN(_05637_ ) );
NAND3_X1 _13364_ ( .A1(_05582_ ), .A2(\mepc [19] ), .A3(_05605_ ), .ZN(_05638_ ) );
BUF_X4 _13365_ ( .A(_05500_ ), .Z(_05639_ ) );
BUF_X4 _13366_ ( .A(_05502_ ), .Z(_05640_ ) );
NAND4_X1 _13367_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_05640_ ), .A4(_05589_ ), .ZN(_05641_ ) );
AND2_X1 _13368_ ( .A1(_05638_ ), .A2(_05641_ ), .ZN(_05642_ ) );
BUF_X4 _13369_ ( .A(_05508_ ), .Z(_05643_ ) );
BUF_X4 _13370_ ( .A(_05586_ ), .Z(_05644_ ) );
BUF_X4 _13371_ ( .A(_05512_ ), .Z(_05645_ ) );
NAND4_X1 _13372_ ( .A1(_05643_ ), .A2(_05644_ ), .A3(\mtvec [19] ), .A4(_05645_ ), .ZN(_05646_ ) );
BUF_X4 _13373_ ( .A(_05518_ ), .Z(_05647_ ) );
BUF_X4 _13374_ ( .A(_05521_ ), .Z(_05648_ ) );
NAND3_X1 _13375_ ( .A1(_05647_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_05648_ ), .ZN(_05649_ ) );
NAND4_X1 _13376_ ( .A1(_05642_ ), .A2(_05607_ ), .A3(_05646_ ), .A4(_05649_ ), .ZN(_05650_ ) );
BUF_X4 _13377_ ( .A(_05546_ ), .Z(_05651_ ) );
BUF_X4 _13378_ ( .A(_05651_ ), .Z(_05652_ ) );
NAND2_X1 _13379_ ( .A1(_05650_ ), .A2(_05652_ ), .ZN(_05653_ ) );
BUF_X2 _13380_ ( .A(_05531_ ), .Z(_05654_ ) );
BUF_X2 _13381_ ( .A(_05543_ ), .Z(_05655_ ) );
AND3_X1 _13382_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_05655_ ), .ZN(_05656_ ) );
INV_X1 _13383_ ( .A(_05656_ ), .ZN(_05657_ ) );
AND2_X1 _13384_ ( .A1(_05653_ ), .A2(_05657_ ), .ZN(_05658_ ) );
INV_X1 _13385_ ( .A(_05658_ ), .ZN(_05659_ ) );
OAI211_X1 _13386_ ( .A(_05637_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05659_ ), .ZN(_05660_ ) );
BUF_X4 _13387_ ( .A(_04146_ ), .Z(_05661_ ) );
NOR3_X1 _13388_ ( .A1(_03265_ ), .A2(_05661_ ), .A3(_05479_ ), .ZN(_05662_ ) );
AOI21_X1 _13389_ ( .A(_05662_ ), .B1(_05624_ ), .B2(_05631_ ), .ZN(_05663_ ) );
AOI21_X1 _13390_ ( .A(_04159_ ), .B1(_05660_ ), .B2(_05663_ ), .ZN(_00161_ ) );
INV_X1 _13391_ ( .A(\ID_EX_pc [18] ), .ZN(_05664_ ) );
XNOR2_X1 _13392_ ( .A(_05562_ ), .B(_05664_ ), .ZN(_05665_ ) );
AND3_X1 _13393_ ( .A1(_05628_ ), .A2(_05627_ ), .A3(_04252_ ), .ZN(_05666_ ) );
NOR2_X1 _13394_ ( .A1(_05666_ ), .A2(_05629_ ), .ZN(_05667_ ) );
MUX2_X1 _13395_ ( .A(_05665_ ), .B(_05667_ ), .S(_05475_ ), .Z(_05668_ ) );
OR2_X2 _13396_ ( .A1(_05668_ ), .A2(\ID_EX_typ [3] ), .ZN(_05669_ ) );
BUF_X4 _13397_ ( .A(_05654_ ), .Z(_05670_ ) );
BUF_X4 _13398_ ( .A(_05655_ ), .Z(_05671_ ) );
NAND3_X1 _13399_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_05671_ ), .ZN(_05672_ ) );
NAND3_X1 _13400_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_05593_ ), .ZN(_05673_ ) );
NAND3_X1 _13401_ ( .A1(_05604_ ), .A2(\mepc [18] ), .A3(_05605_ ), .ZN(_05674_ ) );
BUF_X4 _13402_ ( .A(_05505_ ), .Z(_05675_ ) );
NAND4_X1 _13403_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_05640_ ), .A4(_05675_ ), .ZN(_05676_ ) );
AND3_X1 _13404_ ( .A1(_05673_ ), .A2(_05674_ ), .A3(_05676_ ), .ZN(_05677_ ) );
BUF_X4 _13405_ ( .A(_05511_ ), .Z(_05678_ ) );
BUF_X4 _13406_ ( .A(_05678_ ), .Z(_05679_ ) );
NAND4_X1 _13407_ ( .A1(_05643_ ), .A2(_05679_ ), .A3(\mtvec [18] ), .A4(_05645_ ), .ZN(_05680_ ) );
AND3_X1 _13408_ ( .A1(_05677_ ), .A2(_05607_ ), .A3(_05680_ ), .ZN(_05681_ ) );
BUF_X4 _13409_ ( .A(_05545_ ), .Z(_05682_ ) );
OAI21_X1 _13410_ ( .A(_05672_ ), .B1(_05681_ ), .B2(_05682_ ), .ZN(_05683_ ) );
OAI211_X1 _13411_ ( .A(_05669_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05683_ ), .ZN(_05684_ ) );
BUF_X4 _13412_ ( .A(_04146_ ), .Z(_05685_ ) );
NOR4_X1 _13413_ ( .A1(_03266_ ), .A2(_03262_ ), .A3(_05685_ ), .A4(_05600_ ), .ZN(_05686_ ) );
AOI21_X1 _13414_ ( .A(_05686_ ), .B1(_05624_ ), .B2(_05667_ ), .ZN(_05687_ ) );
AOI21_X1 _13415_ ( .A(_04159_ ), .B1(_05684_ ), .B2(_05687_ ), .ZN(_00162_ ) );
AND2_X1 _13416_ ( .A1(_04239_ ), .A2(_04243_ ), .ZN(_05688_ ) );
NOR2_X1 _13417_ ( .A1(_05688_ ), .A2(_04250_ ), .ZN(_05689_ ) );
XNOR2_X1 _13418_ ( .A(_05689_ ), .B(_04244_ ), .ZN(_05690_ ) );
AOI21_X1 _13419_ ( .A(\ID_EX_typ [3] ), .B1(_05626_ ), .B2(_05690_ ), .ZN(_05691_ ) );
NAND3_X1 _13420_ ( .A1(_04170_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05692_ ) );
INV_X1 _13421_ ( .A(\ID_EX_pc [16] ), .ZN(_05693_ ) );
NOR2_X1 _13422_ ( .A1(_05692_ ), .A2(_05693_ ), .ZN(_05694_ ) );
XNOR2_X1 _13423_ ( .A(_05694_ ), .B(\ID_EX_pc [17] ), .ZN(_05695_ ) );
OAI21_X1 _13424_ ( .A(_05691_ ), .B1(_05633_ ), .B2(_05695_ ), .ZN(_05696_ ) );
NAND3_X1 _13425_ ( .A1(_05582_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_05593_ ), .ZN(_05697_ ) );
NAND4_X1 _13426_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(\mtvec [17] ), .A4(_05587_ ), .ZN(_05698_ ) );
AND2_X1 _13427_ ( .A1(_05697_ ), .A2(_05698_ ), .ZN(_05699_ ) );
BUF_X4 _13428_ ( .A(_05583_ ), .Z(_05700_ ) );
NAND3_X1 _13429_ ( .A1(_05592_ ), .A2(\mepc [17] ), .A3(_05700_ ), .ZN(_05701_ ) );
BUF_X4 _13430_ ( .A(_05589_ ), .Z(_05702_ ) );
NAND4_X1 _13431_ ( .A1(_05643_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_05645_ ), .A4(_05702_ ), .ZN(_05703_ ) );
NAND4_X1 _13432_ ( .A1(_05699_ ), .A2(_05608_ ), .A3(_05701_ ), .A4(_05703_ ), .ZN(_05704_ ) );
NAND2_X1 _13433_ ( .A1(_05704_ ), .A2(_05652_ ), .ZN(_05705_ ) );
NAND3_X1 _13434_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_05580_ ), .ZN(_05706_ ) );
AND2_X1 _13435_ ( .A1(_05705_ ), .A2(_05706_ ), .ZN(_05707_ ) );
INV_X1 _13436_ ( .A(_05707_ ), .ZN(_05708_ ) );
OAI211_X1 _13437_ ( .A(_05696_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05708_ ), .ZN(_05709_ ) );
NOR3_X1 _13438_ ( .A1(_03268_ ), .A2(_05661_ ), .A3(_05479_ ), .ZN(_05710_ ) );
AOI21_X1 _13439_ ( .A(_05710_ ), .B1(_05624_ ), .B2(_05690_ ), .ZN(_05711_ ) );
AOI21_X1 _13440_ ( .A(_04159_ ), .B1(_05709_ ), .B2(_05711_ ), .ZN(_00163_ ) );
BUF_X4 _13441_ ( .A(_05479_ ), .Z(_05712_ ) );
BUF_X4 _13442_ ( .A(_05482_ ), .Z(_05713_ ) );
NAND3_X1 _13443_ ( .A1(_05518_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_05521_ ), .ZN(_05714_ ) );
NAND3_X1 _13444_ ( .A1(_05518_ ), .A2(\mepc [16] ), .A3(_05583_ ), .ZN(_05715_ ) );
AND2_X1 _13445_ ( .A1(_05714_ ), .A2(_05715_ ), .ZN(_05716_ ) );
BUF_X4 _13446_ ( .A(_05500_ ), .Z(_05717_ ) );
BUF_X4 _13447_ ( .A(_05502_ ), .Z(_05718_ ) );
NAND4_X1 _13448_ ( .A1(_05717_ ), .A2(_05678_ ), .A3(\mtvec [16] ), .A4(_05718_ ), .ZN(_05719_ ) );
NAND4_X1 _13449_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_05718_ ), .A4(_05675_ ), .ZN(_05720_ ) );
NAND4_X1 _13450_ ( .A1(_05716_ ), .A2(_05608_ ), .A3(_05719_ ), .A4(_05720_ ), .ZN(_05721_ ) );
NAND2_X1 _13451_ ( .A1(_05721_ ), .A2(_05651_ ), .ZN(_05722_ ) );
AND3_X1 _13452_ ( .A1(_05531_ ), .A2(\EX_LS_result_csreg_mem [16] ), .A3(_05543_ ), .ZN(_05723_ ) );
INV_X1 _13453_ ( .A(_05723_ ), .ZN(_05724_ ) );
AND2_X1 _13454_ ( .A1(_05722_ ), .A2(_05724_ ), .ZN(_05725_ ) );
INV_X1 _13455_ ( .A(_05725_ ), .ZN(_05726_ ) );
XOR2_X1 _13456_ ( .A(_04239_ ), .B(_04243_ ), .Z(_05727_ ) );
AND2_X1 _13457_ ( .A1(_05633_ ), .A2(_05727_ ), .ZN(_05728_ ) );
XNOR2_X1 _13458_ ( .A(_05692_ ), .B(_05693_ ), .ZN(_05729_ ) );
OAI21_X1 _13459_ ( .A(_05482_ ), .B1(_05633_ ), .B2(_05729_ ), .ZN(_05730_ ) );
OAI221_X1 _13460_ ( .A(_05712_ ), .B1(_05713_ ), .B2(_05726_ ), .C1(_05728_ ), .C2(_05730_ ), .ZN(_05731_ ) );
BUF_X4 _13461_ ( .A(_04146_ ), .Z(_05732_ ) );
NOR4_X1 _13462_ ( .A1(_03269_ ), .A2(_03259_ ), .A3(_05732_ ), .A4(_05600_ ), .ZN(_05733_ ) );
AOI21_X1 _13463_ ( .A(_05733_ ), .B1(_05624_ ), .B2(_05727_ ), .ZN(_05734_ ) );
AOI21_X1 _13464_ ( .A(_04159_ ), .B1(_05731_ ), .B2(_05734_ ), .ZN(_00164_ ) );
INV_X1 _13465_ ( .A(_04224_ ), .ZN(_05735_ ) );
OAI21_X1 _13466_ ( .A(_04229_ ), .B1(_04213_ ), .B2(_04221_ ), .ZN(_05736_ ) );
AOI21_X1 _13467_ ( .A(_05735_ ), .B1(_05736_ ), .B2(_04237_ ), .ZN(_05737_ ) );
NOR2_X1 _13468_ ( .A1(_05737_ ), .A2(_04231_ ), .ZN(_05738_ ) );
XNOR2_X1 _13469_ ( .A(_05738_ ), .B(_04223_ ), .ZN(_05739_ ) );
AOI21_X1 _13470_ ( .A(\ID_EX_typ [3] ), .B1(_05626_ ), .B2(_05739_ ), .ZN(_05740_ ) );
AND2_X1 _13471_ ( .A1(_04170_ ), .A2(\ID_EX_pc [14] ), .ZN(_05741_ ) );
XNOR2_X1 _13472_ ( .A(_05741_ ), .B(\ID_EX_pc [15] ), .ZN(_05742_ ) );
OAI21_X1 _13473_ ( .A(_05740_ ), .B1(_05633_ ), .B2(_05742_ ), .ZN(_05743_ ) );
NAND3_X1 _13474_ ( .A1(_05582_ ), .A2(\mepc [15] ), .A3(_05605_ ), .ZN(_05744_ ) );
NAND4_X1 _13475_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_05640_ ), .A4(_05589_ ), .ZN(_05745_ ) );
AND2_X1 _13476_ ( .A1(_05744_ ), .A2(_05745_ ), .ZN(_05746_ ) );
NAND4_X1 _13477_ ( .A1(_05643_ ), .A2(_05644_ ), .A3(\mtvec [15] ), .A4(_05645_ ), .ZN(_05747_ ) );
NAND3_X1 _13478_ ( .A1(_05592_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_05648_ ), .ZN(_05748_ ) );
NAND4_X1 _13479_ ( .A1(_05746_ ), .A2(_05607_ ), .A3(_05747_ ), .A4(_05748_ ), .ZN(_05749_ ) );
NAND2_X1 _13480_ ( .A1(_05749_ ), .A2(_05651_ ), .ZN(_05750_ ) );
NAND3_X1 _13481_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_05580_ ), .ZN(_05751_ ) );
AND2_X1 _13482_ ( .A1(_05750_ ), .A2(_05751_ ), .ZN(_05752_ ) );
INV_X1 _13483_ ( .A(_05752_ ), .ZN(_05753_ ) );
OAI211_X1 _13484_ ( .A(_05743_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05753_ ), .ZN(_05754_ ) );
NOR3_X1 _13485_ ( .A1(_03277_ ), .A2(_05661_ ), .A3(_05479_ ), .ZN(_05755_ ) );
AOI21_X1 _13486_ ( .A(_05755_ ), .B1(_05624_ ), .B2(_05739_ ), .ZN(_05756_ ) );
AOI21_X1 _13487_ ( .A(_04159_ ), .B1(_05754_ ), .B2(_05756_ ), .ZN(_00165_ ) );
BUF_X4 _13488_ ( .A(_04142_ ), .Z(_05757_ ) );
NAND3_X1 _13489_ ( .A1(_05494_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_05521_ ), .ZN(_05758_ ) );
NAND3_X1 _13490_ ( .A1(_05494_ ), .A2(\mepc [14] ), .A3(_05498_ ), .ZN(_05759_ ) );
AND2_X1 _13491_ ( .A1(_05758_ ), .A2(_05759_ ), .ZN(_05760_ ) );
NAND4_X1 _13492_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(\mtvec [14] ), .A4(_05587_ ), .ZN(_05761_ ) );
NAND4_X1 _13493_ ( .A1(_05508_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_05512_ ), .A4(_05589_ ), .ZN(_05762_ ) );
NAND4_X1 _13494_ ( .A1(_05760_ ), .A2(_05608_ ), .A3(_05761_ ), .A4(_05762_ ), .ZN(_05763_ ) );
NAND2_X1 _13495_ ( .A1(_05763_ ), .A2(_05651_ ), .ZN(_05764_ ) );
AND3_X1 _13496_ ( .A1(_05531_ ), .A2(\EX_LS_result_csreg_mem [14] ), .A3(_05543_ ), .ZN(_05765_ ) );
INV_X1 _13497_ ( .A(_05765_ ), .ZN(_05766_ ) );
AND2_X1 _13498_ ( .A1(_05764_ ), .A2(_05766_ ), .ZN(_05767_ ) );
INV_X1 _13499_ ( .A(_05767_ ), .ZN(_05768_ ) );
INV_X1 _13500_ ( .A(\ID_EX_pc [14] ), .ZN(_05769_ ) );
XNOR2_X1 _13501_ ( .A(_04170_ ), .B(_05769_ ), .ZN(_05770_ ) );
AND3_X1 _13502_ ( .A1(_05736_ ), .A2(_05735_ ), .A3(_04237_ ), .ZN(_05771_ ) );
NOR2_X1 _13503_ ( .A1(_05771_ ), .A2(_05737_ ), .ZN(_05772_ ) );
MUX2_X1 _13504_ ( .A(_05770_ ), .B(_05772_ ), .S(_05475_ ), .Z(_05773_ ) );
MUX2_X2 _13505_ ( .A(_05768_ ), .B(_05773_ ), .S(_05482_ ), .Z(_05774_ ) );
NAND2_X1 _13506_ ( .A1(_05774_ ), .A2(_05620_ ), .ZN(_05775_ ) );
BUF_X4 _13507_ ( .A(_05622_ ), .Z(_05776_ ) );
BUF_X4 _13508_ ( .A(_04147_ ), .Z(_05777_ ) );
AOI22_X1 _13509_ ( .A1(_03278_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_05772_ ), .ZN(_05778_ ) );
AOI21_X1 _13510_ ( .A(_05757_ ), .B1(_05775_ ), .B2(_05778_ ), .ZN(_00166_ ) );
NAND3_X1 _13511_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [13] ), .A3(_05655_ ), .ZN(_05779_ ) );
NAND3_X1 _13512_ ( .A1(_05582_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_05593_ ), .ZN(_05780_ ) );
NAND2_X1 _13513_ ( .A1(_05780_ ), .A2(_05517_ ), .ZN(_05781_ ) );
AND3_X1 _13514_ ( .A1(_05518_ ), .A2(\mepc [13] ), .A3(_05583_ ), .ZN(_05782_ ) );
AND4_X1 _13515_ ( .A1(\mtvec [13] ), .A2(_05508_ ), .A3(_05511_ ), .A4(_05512_ ), .ZN(_05783_ ) );
AND4_X1 _13516_ ( .A1(\mycsreg.CSReg[0][13] ), .A2(_05508_ ), .A3(_05512_ ), .A4(_05589_ ), .ZN(_05784_ ) );
NOR4_X1 _13517_ ( .A1(_05781_ ), .A2(_05782_ ), .A3(_05783_ ), .A4(_05784_ ), .ZN(_05785_ ) );
OAI21_X1 _13518_ ( .A(_05779_ ), .B1(_05785_ ), .B2(_05545_ ), .ZN(_05786_ ) );
XNOR2_X1 _13519_ ( .A(_04169_ ), .B(_05559_ ), .ZN(_05787_ ) );
OAI21_X1 _13520_ ( .A(_04226_ ), .B1(_04213_ ), .B2(_04221_ ), .ZN(_05788_ ) );
NAND2_X1 _13521_ ( .A1(_05788_ ), .A2(_04235_ ), .ZN(_05789_ ) );
XNOR2_X1 _13522_ ( .A(_05789_ ), .B(_04228_ ), .ZN(_05790_ ) );
MUX2_X1 _13523_ ( .A(_05787_ ), .B(_05790_ ), .S(_05475_ ), .Z(_05791_ ) );
MUX2_X2 _13524_ ( .A(_05786_ ), .B(_05791_ ), .S(_05482_ ), .Z(_05792_ ) );
NAND2_X1 _13525_ ( .A1(_05792_ ), .A2(_05620_ ), .ZN(_05793_ ) );
NOR3_X1 _13526_ ( .A1(_03282_ ), .A2(_05661_ ), .A3(_05479_ ), .ZN(_05794_ ) );
AOI21_X1 _13527_ ( .A(_05794_ ), .B1(_05624_ ), .B2(_05790_ ), .ZN(_05795_ ) );
AOI21_X1 _13528_ ( .A(_05757_ ), .B1(_05793_ ), .B2(_05795_ ), .ZN(_00167_ ) );
XNOR2_X1 _13529_ ( .A(_04222_ ), .B(_04227_ ), .ZN(_05796_ ) );
NAND2_X1 _13530_ ( .A1(_05626_ ), .A2(_05796_ ), .ZN(_05797_ ) );
XNOR2_X1 _13531_ ( .A(_04168_ ), .B(_05560_ ), .ZN(_05798_ ) );
OAI21_X1 _13532_ ( .A(_05798_ ), .B1(_05471_ ), .B2(_05473_ ), .ZN(_05799_ ) );
NAND3_X1 _13533_ ( .A1(_05797_ ), .A2(_05556_ ), .A3(_05799_ ), .ZN(_05800_ ) );
NAND3_X1 _13534_ ( .A1(_05582_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_05593_ ), .ZN(_05801_ ) );
NAND3_X1 _13535_ ( .A1(_05582_ ), .A2(\mepc [12] ), .A3(_05583_ ), .ZN(_05802_ ) );
AND2_X1 _13536_ ( .A1(_05801_ ), .A2(_05802_ ), .ZN(_05803_ ) );
NAND4_X1 _13537_ ( .A1(_05643_ ), .A2(_05644_ ), .A3(\mtvec [12] ), .A4(_05645_ ), .ZN(_05804_ ) );
NAND4_X1 _13538_ ( .A1(_05643_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_05645_ ), .A4(_05702_ ), .ZN(_05805_ ) );
NAND4_X1 _13539_ ( .A1(_05803_ ), .A2(_05608_ ), .A3(_05804_ ), .A4(_05805_ ), .ZN(_05806_ ) );
NAND2_X1 _13540_ ( .A1(_05806_ ), .A2(_05651_ ), .ZN(_05807_ ) );
AND3_X1 _13541_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [12] ), .A3(_05655_ ), .ZN(_05808_ ) );
INV_X1 _13542_ ( .A(_05808_ ), .ZN(_05809_ ) );
AND2_X1 _13543_ ( .A1(_05807_ ), .A2(_05809_ ), .ZN(_05810_ ) );
INV_X1 _13544_ ( .A(_05810_ ), .ZN(_05811_ ) );
OAI211_X1 _13545_ ( .A(_05800_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05811_ ), .ZN(_05812_ ) );
AOI22_X1 _13546_ ( .A1(_03283_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_05796_ ), .ZN(_05813_ ) );
AOI21_X1 _13547_ ( .A(_05757_ ), .B1(_05812_ ), .B2(_05813_ ), .ZN(_00168_ ) );
XNOR2_X1 _13548_ ( .A(_04167_ ), .B(\ID_EX_pc [11] ), .ZN(_05814_ ) );
INV_X1 _13549_ ( .A(_04208_ ), .ZN(_05815_ ) );
OAI21_X1 _13550_ ( .A(_04212_ ), .B1(_04204_ ), .B2(_04205_ ), .ZN(_05816_ ) );
AOI21_X1 _13551_ ( .A(_05815_ ), .B1(_05816_ ), .B2(_04219_ ), .ZN(_05817_ ) );
OR2_X1 _13552_ ( .A1(_05817_ ), .A2(_04214_ ), .ZN(_05818_ ) );
XNOR2_X1 _13553_ ( .A(_05818_ ), .B(_04207_ ), .ZN(_05819_ ) );
MUX2_X1 _13554_ ( .A(_05814_ ), .B(_05819_ ), .S(_05626_ ), .Z(_05820_ ) );
NAND2_X1 _13555_ ( .A1(_05820_ ), .A2(_05556_ ), .ZN(_05821_ ) );
NAND3_X1 _13556_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [11] ), .A3(_05671_ ), .ZN(_05822_ ) );
NAND3_X1 _13557_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_05593_ ), .ZN(_05823_ ) );
NAND3_X1 _13558_ ( .A1(_05604_ ), .A2(\mepc [11] ), .A3(_05605_ ), .ZN(_05824_ ) );
NAND4_X1 _13559_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_05640_ ), .A4(_05675_ ), .ZN(_05825_ ) );
AND3_X1 _13560_ ( .A1(_05823_ ), .A2(_05824_ ), .A3(_05825_ ), .ZN(_05826_ ) );
NAND4_X1 _13561_ ( .A1(_05643_ ), .A2(_05679_ ), .A3(\mtvec [11] ), .A4(_05645_ ), .ZN(_05827_ ) );
AND3_X1 _13562_ ( .A1(_05826_ ), .A2(_05608_ ), .A3(_05827_ ), .ZN(_05828_ ) );
OAI21_X1 _13563_ ( .A(_05822_ ), .B1(_05828_ ), .B2(_05682_ ), .ZN(_05829_ ) );
OAI211_X1 _13564_ ( .A(_05821_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05829_ ), .ZN(_05830_ ) );
NOR2_X1 _13565_ ( .A1(_05819_ ), .A2(_04148_ ), .ZN(_05831_ ) );
AOI21_X1 _13566_ ( .A(_03128_ ), .B1(_02925_ ), .B2(_03072_ ), .ZN(_05832_ ) );
AOI21_X1 _13567_ ( .A(\ID_EX_imm [10] ), .B1(_03073_ ), .B2(_03093_ ), .ZN(_05833_ ) );
NOR3_X1 _13568_ ( .A1(_05832_ ), .A2(_03130_ ), .A3(_05833_ ), .ZN(_05834_ ) );
NOR2_X1 _13569_ ( .A1(_05834_ ), .A2(_03130_ ), .ZN(_05835_ ) );
XNOR2_X1 _13570_ ( .A(_05835_ ), .B(_03121_ ), .ZN(_05836_ ) );
AOI21_X1 _13571_ ( .A(_05831_ ), .B1(_05836_ ), .B2(_05776_ ), .ZN(_05837_ ) );
AOI21_X1 _13572_ ( .A(_05757_ ), .B1(_05830_ ), .B2(_05837_ ), .ZN(_00169_ ) );
CLKBUF_X2 _13573_ ( .A(_04145_ ), .Z(_05838_ ) );
INV_X1 _13574_ ( .A(\ID_EX_pc [28] ), .ZN(_05839_ ) );
XNOR2_X1 _13575_ ( .A(_05569_ ), .B(_05839_ ), .ZN(_05840_ ) );
AOI21_X1 _13576_ ( .A(\ID_EX_typ [3] ), .B1(_05573_ ), .B2(_05840_ ), .ZN(_05841_ ) );
AND4_X1 _13577_ ( .A1(_04104_ ), .A2(_05534_ ), .A3(_05539_ ), .A4(_05526_ ), .ZN(_05842_ ) );
AND4_X1 _13578_ ( .A1(_05535_ ), .A2(_05529_ ), .A3(_05524_ ), .A4(_05525_ ), .ZN(_05843_ ) );
NAND2_X1 _13579_ ( .A1(_05842_ ), .A2(_05843_ ), .ZN(_05844_ ) );
AND3_X1 _13580_ ( .A1(_05541_ ), .A2(_05542_ ), .A3(_05527_ ), .ZN(_05845_ ) );
NAND3_X1 _13581_ ( .A1(_05845_ ), .A2(_05536_ ), .A3(_05530_ ), .ZN(_05846_ ) );
OR3_X1 _13582_ ( .A1(_05844_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_05846_ ), .ZN(_05847_ ) );
AND3_X1 _13583_ ( .A1(_05489_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_05848_ ) );
AND3_X1 _13584_ ( .A1(_05501_ ), .A2(_05485_ ), .A3(\ID_EX_csr [4] ), .ZN(_05849_ ) );
AND2_X1 _13585_ ( .A1(_05848_ ), .A2(_05849_ ), .ZN(_05850_ ) );
AND2_X1 _13586_ ( .A1(_05850_ ), .A2(_05583_ ), .ZN(_05851_ ) );
INV_X1 _13587_ ( .A(_05851_ ), .ZN(_05852_ ) );
NAND3_X1 _13588_ ( .A1(_05494_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_05521_ ), .ZN(_05853_ ) );
NAND3_X1 _13589_ ( .A1(_05501_ ), .A2(_05485_ ), .A3(_05486_ ), .ZN(_05854_ ) );
NAND3_X1 _13590_ ( .A1(_05487_ ), .A2(\ID_EX_csr [9] ), .A3(\ID_EX_csr [8] ), .ZN(_05855_ ) );
NOR3_X1 _13591_ ( .A1(_05854_ ), .A2(\ID_EX_csr [10] ), .A3(_05855_ ), .ZN(_05856_ ) );
BUF_X4 _13592_ ( .A(_05856_ ), .Z(_05857_ ) );
NAND3_X1 _13593_ ( .A1(_05857_ ), .A2(\mtvec [28] ), .A3(_05644_ ), .ZN(_05858_ ) );
NAND3_X1 _13594_ ( .A1(_05852_ ), .A2(_05853_ ), .A3(_05858_ ), .ZN(_05859_ ) );
NAND3_X1 _13595_ ( .A1(_05494_ ), .A2(\mepc [28] ), .A3(_05583_ ), .ZN(_05860_ ) );
BUF_X4 _13596_ ( .A(_05856_ ), .Z(_05861_ ) );
NAND3_X1 _13597_ ( .A1(_05861_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_05702_ ), .ZN(_05862_ ) );
BUF_X2 _13598_ ( .A(_05844_ ), .Z(_05863_ ) );
BUF_X2 _13599_ ( .A(_05846_ ), .Z(_05864_ ) );
OAI211_X1 _13600_ ( .A(_05860_ ), .B(_05862_ ), .C1(_05863_ ), .C2(_05864_ ), .ZN(_05865_ ) );
OAI21_X1 _13601_ ( .A(_05847_ ), .B1(_05859_ ), .B2(_05865_ ), .ZN(_05866_ ) );
AOI211_X2 _13602_ ( .A(_05838_ ), .B(_05841_ ), .C1(\ID_EX_typ [3] ), .C2(_05866_ ), .ZN(_05867_ ) );
XNOR2_X1 _13603_ ( .A(_04281_ ), .B(_04282_ ), .ZN(_05868_ ) );
NAND3_X1 _13604_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_05655_ ), .ZN(_05869_ ) );
NAND4_X1 _13605_ ( .A1(_05500_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_05502_ ), .A4(_05505_ ), .ZN(_05870_ ) );
AND3_X1 _13606_ ( .A1(_05853_ ), .A2(_05860_ ), .A3(_05870_ ), .ZN(_05871_ ) );
NAND4_X1 _13607_ ( .A1(_05717_ ), .A2(_05678_ ), .A3(\mtvec [28] ), .A4(_05718_ ), .ZN(_05872_ ) );
AND3_X1 _13608_ ( .A1(_05871_ ), .A2(_05517_ ), .A3(_05872_ ), .ZN(_05873_ ) );
OAI21_X1 _13609_ ( .A(_05869_ ), .B1(_05873_ ), .B2(_05545_ ), .ZN(_05874_ ) );
OAI211_X1 _13610_ ( .A(_05626_ ), .B(_05600_ ), .C1(_05482_ ), .C2(_05874_ ), .ZN(_05875_ ) );
AOI21_X1 _13611_ ( .A(_05868_ ), .B1(_05875_ ), .B2(_04148_ ), .ZN(_05876_ ) );
NOR2_X1 _13612_ ( .A1(_05867_ ), .A2(_05876_ ), .ZN(_05877_ ) );
NAND2_X1 _13613_ ( .A1(_03288_ ), .A2(_05776_ ), .ZN(_05878_ ) );
AOI21_X1 _13614_ ( .A(_05757_ ), .B1(_05877_ ), .B2(_05878_ ), .ZN(_00170_ ) );
NAND3_X1 _13615_ ( .A1(_05494_ ), .A2(\mepc [10] ), .A3(_05498_ ), .ZN(_05879_ ) );
NAND4_X1 _13616_ ( .A1(_05500_ ), .A2(\mycsreg.CSReg[0][10] ), .A3(_05502_ ), .A4(_05505_ ), .ZN(_05880_ ) );
AND2_X1 _13617_ ( .A1(_05879_ ), .A2(_05880_ ), .ZN(_05881_ ) );
NAND4_X1 _13618_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(\mtvec [10] ), .A4(_05587_ ), .ZN(_05882_ ) );
NAND3_X1 _13619_ ( .A1(_05518_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_05593_ ), .ZN(_05883_ ) );
NAND4_X1 _13620_ ( .A1(_05881_ ), .A2(_05607_ ), .A3(_05882_ ), .A4(_05883_ ), .ZN(_05884_ ) );
NAND2_X1 _13621_ ( .A1(_05884_ ), .A2(_05651_ ), .ZN(_05885_ ) );
AND3_X1 _13622_ ( .A1(_05531_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_05543_ ), .ZN(_05886_ ) );
INV_X1 _13623_ ( .A(_05886_ ), .ZN(_05887_ ) );
AND2_X1 _13624_ ( .A1(_05885_ ), .A2(_05887_ ), .ZN(_05888_ ) );
INV_X1 _13625_ ( .A(_05888_ ), .ZN(_05889_ ) );
INV_X1 _13626_ ( .A(\ID_EX_pc [10] ), .ZN(_05890_ ) );
XNOR2_X1 _13627_ ( .A(_04166_ ), .B(_05890_ ), .ZN(_05891_ ) );
AND3_X1 _13628_ ( .A1(_05816_ ), .A2(_05815_ ), .A3(_04219_ ), .ZN(_05892_ ) );
NOR2_X1 _13629_ ( .A1(_05892_ ), .A2(_05817_ ), .ZN(_05893_ ) );
MUX2_X1 _13630_ ( .A(_05891_ ), .B(_05893_ ), .S(_05475_ ), .Z(_05894_ ) );
MUX2_X2 _13631_ ( .A(_05889_ ), .B(_05894_ ), .S(_05481_ ), .Z(_05895_ ) );
NAND2_X1 _13632_ ( .A1(_05895_ ), .A2(_05620_ ), .ZN(_05896_ ) );
XNOR2_X1 _13633_ ( .A(_05832_ ), .B(_03097_ ), .ZN(_05897_ ) );
AOI22_X1 _13634_ ( .A1(_05897_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_05893_ ), .ZN(_05898_ ) );
AOI21_X1 _13635_ ( .A(_05757_ ), .B1(_05896_ ), .B2(_05898_ ), .ZN(_00171_ ) );
INV_X1 _13636_ ( .A(\ID_EX_pc [9] ), .ZN(_05899_ ) );
XNOR2_X1 _13637_ ( .A(_04165_ ), .B(_05899_ ), .ZN(_05900_ ) );
AND2_X1 _13638_ ( .A1(_04206_ ), .A2(_04210_ ), .ZN(_05901_ ) );
NOR2_X1 _13639_ ( .A1(_05901_ ), .A2(_04217_ ), .ZN(_05902_ ) );
XNOR2_X1 _13640_ ( .A(_05902_ ), .B(_04211_ ), .ZN(_05903_ ) );
MUX2_X1 _13641_ ( .A(_05900_ ), .B(_05903_ ), .S(_05475_ ), .Z(_05904_ ) );
OR2_X2 _13642_ ( .A1(_05904_ ), .A2(\ID_EX_typ [3] ), .ZN(_05905_ ) );
NAND3_X1 _13643_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_05671_ ), .ZN(_05906_ ) );
NAND3_X1 _13644_ ( .A1(_05604_ ), .A2(\mepc [9] ), .A3(_05605_ ), .ZN(_05907_ ) );
NAND4_X1 _13645_ ( .A1(_05639_ ), .A2(_05586_ ), .A3(\mtvec [9] ), .A4(_05640_ ), .ZN(_05908_ ) );
NAND4_X1 _13646_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][9] ), .A3(_05640_ ), .A4(_05675_ ), .ZN(_05909_ ) );
AND3_X1 _13647_ ( .A1(_05907_ ), .A2(_05908_ ), .A3(_05909_ ), .ZN(_05910_ ) );
BUF_X2 _13648_ ( .A(_05582_ ), .Z(_05911_ ) );
NAND3_X1 _13649_ ( .A1(_05911_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_05594_ ), .ZN(_05912_ ) );
AND3_X1 _13650_ ( .A1(_05910_ ), .A2(_05607_ ), .A3(_05912_ ), .ZN(_05913_ ) );
OAI21_X1 _13651_ ( .A(_05906_ ), .B1(_05913_ ), .B2(_05682_ ), .ZN(_05914_ ) );
OAI211_X1 _13652_ ( .A(_05905_ ), .B(_05480_ ), .C1(_05483_ ), .C2(_05914_ ), .ZN(_05915_ ) );
NAND2_X1 _13653_ ( .A1(_02925_ ), .A2(_03046_ ), .ZN(_05916_ ) );
AND2_X1 _13654_ ( .A1(_05916_ ), .A2(_03127_ ), .ZN(_05917_ ) );
XNOR2_X1 _13655_ ( .A(_05917_ ), .B(_03126_ ), .ZN(_05918_ ) );
NOR3_X1 _13656_ ( .A1(_05918_ ), .A2(_05661_ ), .A3(_05600_ ), .ZN(_05919_ ) );
AOI21_X1 _13657_ ( .A(_05919_ ), .B1(_05624_ ), .B2(_05903_ ), .ZN(_05920_ ) );
AOI21_X1 _13658_ ( .A(_05757_ ), .B1(_05915_ ), .B2(_05920_ ), .ZN(_00172_ ) );
BUF_X4 _13659_ ( .A(_05479_ ), .Z(_05921_ ) );
NAND3_X1 _13660_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [8] ), .A3(_05671_ ), .ZN(_05922_ ) );
NAND3_X1 _13661_ ( .A1(_05582_ ), .A2(\mepc [8] ), .A3(_05583_ ), .ZN(_05923_ ) );
NAND4_X1 _13662_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(\mtvec [8] ), .A4(_05587_ ), .ZN(_05924_ ) );
NAND4_X1 _13663_ ( .A1(_05585_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_05587_ ), .A4(_05589_ ), .ZN(_05925_ ) );
AND3_X1 _13664_ ( .A1(_05923_ ), .A2(_05924_ ), .A3(_05925_ ), .ZN(_05926_ ) );
NAND3_X1 _13665_ ( .A1(_05592_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_05594_ ), .ZN(_05927_ ) );
AND3_X1 _13666_ ( .A1(_05926_ ), .A2(_05608_ ), .A3(_05927_ ), .ZN(_05928_ ) );
OAI21_X1 _13667_ ( .A(_05922_ ), .B1(_05928_ ), .B2(_05682_ ), .ZN(_05929_ ) );
XOR2_X1 _13668_ ( .A(_04206_ ), .B(_04210_ ), .Z(_05930_ ) );
AND2_X1 _13669_ ( .A1(_05633_ ), .A2(_05930_ ), .ZN(_05931_ ) );
XNOR2_X1 _13670_ ( .A(_04164_ ), .B(\ID_EX_pc [8] ), .ZN(_05932_ ) );
OAI21_X1 _13671_ ( .A(_05482_ ), .B1(_05633_ ), .B2(_05932_ ), .ZN(_05933_ ) );
OAI221_X1 _13672_ ( .A(_05921_ ), .B1(_05556_ ), .B2(_05929_ ), .C1(_05931_ ), .C2(_05933_ ), .ZN(_05934_ ) );
XOR2_X1 _13673_ ( .A(_02925_ ), .B(_03046_ ), .Z(_05935_ ) );
AOI22_X1 _13674_ ( .A1(_05935_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_05930_ ), .ZN(_05936_ ) );
AOI21_X1 _13675_ ( .A(_05757_ ), .B1(_05934_ ), .B2(_05936_ ), .ZN(_00173_ ) );
NAND3_X1 _13676_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_05580_ ), .ZN(_05937_ ) );
NAND3_X1 _13677_ ( .A1(_05604_ ), .A2(\mepc [7] ), .A3(_05605_ ), .ZN(_05938_ ) );
NAND3_X1 _13678_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_05593_ ), .ZN(_05939_ ) );
NAND4_X1 _13679_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_05640_ ), .A4(_05675_ ), .ZN(_05940_ ) );
NAND4_X1 _13680_ ( .A1(_05639_ ), .A2(_05586_ ), .A3(\mtvec [7] ), .A4(_05640_ ), .ZN(_05941_ ) );
AND4_X1 _13681_ ( .A1(_05938_ ), .A2(_05939_ ), .A3(_05940_ ), .A4(_05941_ ), .ZN(_05942_ ) );
OAI21_X1 _13682_ ( .A(_05937_ ), .B1(_05942_ ), .B2(_05545_ ), .ZN(_05943_ ) );
INV_X1 _13683_ ( .A(\ID_EX_pc [7] ), .ZN(_05944_ ) );
XNOR2_X1 _13684_ ( .A(_04163_ ), .B(_05944_ ), .ZN(_05945_ ) );
NAND2_X1 _13685_ ( .A1(_04202_ ), .A2(_04203_ ), .ZN(_05946_ ) );
XNOR2_X1 _13686_ ( .A(\ID_EX_pc [7] ), .B(\ID_EX_imm [7] ), .ZN(_05947_ ) );
XNOR2_X1 _13687_ ( .A(_05946_ ), .B(_05947_ ), .ZN(_05948_ ) );
MUX2_X1 _13688_ ( .A(_05945_ ), .B(_05948_ ), .S(_05475_ ), .Z(_05949_ ) );
MUX2_X2 _13689_ ( .A(_05943_ ), .B(_05949_ ), .S(_05481_ ), .Z(_05950_ ) );
NAND2_X1 _13690_ ( .A1(_05950_ ), .A2(_05620_ ), .ZN(_05951_ ) );
NOR2_X1 _13691_ ( .A1(_02913_ ), .A2(_02914_ ), .ZN(_05952_ ) );
NOR3_X1 _13692_ ( .A1(_05952_ ), .A2(_02765_ ), .A3(_02738_ ), .ZN(_05953_ ) );
OAI21_X1 _13693_ ( .A(_02789_ ), .B1(_05953_ ), .B2(_02923_ ), .ZN(_05954_ ) );
NAND2_X1 _13694_ ( .A1(_05954_ ), .A2(_02917_ ), .ZN(_05955_ ) );
XNOR2_X1 _13695_ ( .A(_05955_ ), .B(_02916_ ), .ZN(_05956_ ) );
AOI22_X1 _13696_ ( .A1(_05956_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_05948_ ), .ZN(_05957_ ) );
AOI21_X1 _13697_ ( .A(_05757_ ), .B1(_05951_ ), .B2(_05957_ ), .ZN(_00174_ ) );
INV_X1 _13698_ ( .A(\ID_EX_pc [6] ), .ZN(_05958_ ) );
XNOR2_X1 _13699_ ( .A(_04162_ ), .B(_05958_ ), .ZN(_05959_ ) );
XOR2_X1 _13700_ ( .A(_04200_ ), .B(_04201_ ), .Z(_05960_ ) );
MUX2_X1 _13701_ ( .A(_05959_ ), .B(_05960_ ), .S(_05475_ ), .Z(_05961_ ) );
OR2_X2 _13702_ ( .A1(_05961_ ), .A2(\ID_EX_typ [3] ), .ZN(_05962_ ) );
NAND4_X1 _13703_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(\mtvec [6] ), .A4(_05587_ ), .ZN(_05963_ ) );
AND2_X1 _13704_ ( .A1(_05517_ ), .A2(_05963_ ), .ZN(_05964_ ) );
NAND3_X1 _13705_ ( .A1(_05592_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_05648_ ), .ZN(_05965_ ) );
NAND3_X1 _13706_ ( .A1(_05647_ ), .A2(\mepc [6] ), .A3(_05700_ ), .ZN(_05966_ ) );
NAND4_X1 _13707_ ( .A1(_05643_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_05645_ ), .A4(_05702_ ), .ZN(_05967_ ) );
NAND4_X1 _13708_ ( .A1(_05964_ ), .A2(_05965_ ), .A3(_05966_ ), .A4(_05967_ ), .ZN(_05968_ ) );
NAND2_X1 _13709_ ( .A1(_05652_ ), .A2(_05968_ ), .ZN(_05969_ ) );
AND3_X1 _13710_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [6] ), .A3(_05655_ ), .ZN(_05970_ ) );
INV_X1 _13711_ ( .A(_05970_ ), .ZN(_05971_ ) );
AND2_X1 _13712_ ( .A1(_05969_ ), .A2(_05971_ ), .ZN(_05972_ ) );
INV_X1 _13713_ ( .A(_05972_ ), .ZN(_05973_ ) );
OAI211_X1 _13714_ ( .A(_05962_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_05973_ ), .ZN(_05974_ ) );
OR3_X1 _13715_ ( .A1(_05953_ ), .A2(_02923_ ), .A3(_02789_ ), .ZN(_05975_ ) );
AND2_X1 _13716_ ( .A1(_05975_ ), .A2(_05954_ ), .ZN(_05976_ ) );
AOI22_X1 _13717_ ( .A1(_05976_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_05960_ ), .ZN(_05977_ ) );
AOI21_X1 _13718_ ( .A(_05757_ ), .B1(_05974_ ), .B2(_05977_ ), .ZN(_00175_ ) );
BUF_X4 _13719_ ( .A(_04142_ ), .Z(_05978_ ) );
NAND3_X1 _13720_ ( .A1(_05647_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_05648_ ), .ZN(_05979_ ) );
NAND4_X1 _13721_ ( .A1(_05717_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_05718_ ), .A4(_05675_ ), .ZN(_05980_ ) );
NAND4_X1 _13722_ ( .A1(_05717_ ), .A2(_05678_ ), .A3(\mtvec [5] ), .A4(_05718_ ), .ZN(_05981_ ) );
NAND3_X1 _13723_ ( .A1(_05979_ ), .A2(_05980_ ), .A3(_05981_ ), .ZN(_05982_ ) );
NAND3_X1 _13724_ ( .A1(_05647_ ), .A2(\mepc [5] ), .A3(_05605_ ), .ZN(_05983_ ) );
NAND2_X1 _13725_ ( .A1(_05983_ ), .A2(_05517_ ), .ZN(_05984_ ) );
OAI21_X1 _13726_ ( .A(_05651_ ), .B1(_05982_ ), .B2(_05984_ ), .ZN(_05985_ ) );
NAND3_X1 _13727_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [5] ), .A3(_05580_ ), .ZN(_05986_ ) );
AND2_X1 _13728_ ( .A1(_05985_ ), .A2(_05986_ ), .ZN(_05987_ ) );
INV_X1 _13729_ ( .A(_05987_ ), .ZN(_05988_ ) );
XNOR2_X1 _13730_ ( .A(\ID_EX_pc [5] ), .B(\ID_EX_imm [5] ), .ZN(_05989_ ) );
XNOR2_X1 _13731_ ( .A(_04196_ ), .B(_05989_ ), .ZN(_05990_ ) );
AND2_X1 _13732_ ( .A1(_05626_ ), .A2(_05990_ ), .ZN(_05991_ ) );
XNOR2_X1 _13733_ ( .A(_04161_ ), .B(\ID_EX_pc [5] ), .ZN(_05992_ ) );
OAI21_X1 _13734_ ( .A(_05482_ ), .B1(_05633_ ), .B2(_05992_ ), .ZN(_05993_ ) );
OAI221_X1 _13735_ ( .A(_05921_ ), .B1(_05556_ ), .B2(_05988_ ), .C1(_05991_ ), .C2(_05993_ ), .ZN(_05994_ ) );
NOR2_X1 _13736_ ( .A1(_05952_ ), .A2(_02738_ ), .ZN(_05995_ ) );
AOI21_X1 _13737_ ( .A(_05995_ ), .B1(\ID_EX_imm [4] ), .B2(_02735_ ), .ZN(_05996_ ) );
XOR2_X1 _13738_ ( .A(_05996_ ), .B(_02765_ ), .Z(_05997_ ) );
AOI22_X1 _13739_ ( .A1(_05997_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_05990_ ), .ZN(_05998_ ) );
AOI21_X1 _13740_ ( .A(_05978_ ), .B1(_05994_ ), .B2(_05998_ ), .ZN(_00176_ ) );
XNOR2_X1 _13741_ ( .A(_04160_ ), .B(\ID_EX_pc [4] ), .ZN(_05999_ ) );
OR2_X1 _13742_ ( .A1(_04192_ ), .A2(_04193_ ), .ZN(_06000_ ) );
XOR2_X1 _13743_ ( .A(_06000_ ), .B(_04183_ ), .Z(_06001_ ) );
INV_X1 _13744_ ( .A(_06001_ ), .ZN(_06002_ ) );
MUX2_X1 _13745_ ( .A(_05999_ ), .B(_06002_ ), .S(_05626_ ), .Z(_06003_ ) );
NAND2_X1 _13746_ ( .A1(_06003_ ), .A2(_05556_ ), .ZN(_06004_ ) );
NAND3_X1 _13747_ ( .A1(_05647_ ), .A2(\mepc [4] ), .A3(_05700_ ), .ZN(_06005_ ) );
NAND4_X1 _13748_ ( .A1(_05717_ ), .A2(_05678_ ), .A3(\mtvec [4] ), .A4(_05718_ ), .ZN(_06006_ ) );
NAND4_X1 _13749_ ( .A1(_05717_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_05718_ ), .A4(_05702_ ), .ZN(_06007_ ) );
NAND3_X1 _13750_ ( .A1(_06005_ ), .A2(_06006_ ), .A3(_06007_ ), .ZN(_06008_ ) );
NAND3_X1 _13751_ ( .A1(_05647_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_05648_ ), .ZN(_06009_ ) );
NAND2_X1 _13752_ ( .A1(_06009_ ), .A2(_05517_ ), .ZN(_06010_ ) );
OAI21_X1 _13753_ ( .A(_05651_ ), .B1(_06008_ ), .B2(_06010_ ), .ZN(_06011_ ) );
NAND3_X1 _13754_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [4] ), .A3(_05580_ ), .ZN(_06012_ ) );
AND2_X1 _13755_ ( .A1(_06011_ ), .A2(_06012_ ), .ZN(_06013_ ) );
INV_X1 _13756_ ( .A(_06013_ ), .ZN(_06014_ ) );
OAI211_X1 _13757_ ( .A(_06004_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06014_ ), .ZN(_06015_ ) );
XNOR2_X1 _13758_ ( .A(_05952_ ), .B(_02737_ ), .ZN(_06016_ ) );
AOI22_X1 _13759_ ( .A1(_06016_ ), .A2(_05776_ ), .B1(_05777_ ), .B2(_06001_ ), .ZN(_06017_ ) );
AOI21_X1 _13760_ ( .A(_05978_ ), .B1(_06015_ ), .B2(_06017_ ), .ZN(_00177_ ) );
NAND3_X1 _13761_ ( .A1(_05647_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_05648_ ), .ZN(_06018_ ) );
NAND4_X1 _13762_ ( .A1(_05717_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_05718_ ), .A4(_05675_ ), .ZN(_06019_ ) );
NAND4_X1 _13763_ ( .A1(_05717_ ), .A2(_05678_ ), .A3(\mtvec [3] ), .A4(_05640_ ), .ZN(_06020_ ) );
NAND3_X1 _13764_ ( .A1(_06018_ ), .A2(_06019_ ), .A3(_06020_ ), .ZN(_06021_ ) );
NAND3_X1 _13765_ ( .A1(_05647_ ), .A2(\mepc [3] ), .A3(_05605_ ), .ZN(_06022_ ) );
NAND2_X1 _13766_ ( .A1(_06022_ ), .A2(_05517_ ), .ZN(_06023_ ) );
OAI21_X1 _13767_ ( .A(_05651_ ), .B1(_06021_ ), .B2(_06023_ ), .ZN(_06024_ ) );
NAND3_X1 _13768_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [3] ), .A3(_05655_ ), .ZN(_06025_ ) );
AND2_X1 _13769_ ( .A1(_06024_ ), .A2(_06025_ ), .ZN(_06026_ ) );
INV_X1 _13770_ ( .A(_06026_ ), .ZN(_06027_ ) );
NAND2_X1 _13771_ ( .A1(_04189_ ), .A2(_04190_ ), .ZN(_06028_ ) );
XOR2_X1 _13772_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_imm [3] ), .Z(_06029_ ) );
XOR2_X1 _13773_ ( .A(_06028_ ), .B(_06029_ ), .Z(_06030_ ) );
INV_X1 _13774_ ( .A(_06030_ ), .ZN(_06031_ ) );
OAI21_X1 _13775_ ( .A(_05556_ ), .B1(_05574_ ), .B2(_06031_ ), .ZN(_06032_ ) );
XNOR2_X1 _13776_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .ZN(_06033_ ) );
NOR2_X1 _13777_ ( .A1(_05633_ ), .A2(_06033_ ), .ZN(_06034_ ) );
OAI221_X1 _13778_ ( .A(_05921_ ), .B1(_05556_ ), .B2(_06027_ ), .C1(_06032_ ), .C2(_06034_ ), .ZN(_06035_ ) );
XOR2_X1 _13779_ ( .A(_02890_ ), .B(_02912_ ), .Z(_06036_ ) );
AOI22_X1 _13780_ ( .A1(_06036_ ), .A2(_05622_ ), .B1(_05777_ ), .B2(_06030_ ), .ZN(_06037_ ) );
AOI21_X1 _13781_ ( .A(_05978_ ), .B1(_06035_ ), .B2(_06037_ ), .ZN(_00178_ ) );
NAND3_X1 _13782_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_05580_ ), .ZN(_06038_ ) );
NAND3_X1 _13783_ ( .A1(_05518_ ), .A2(\mycsreg.CSReg[3][2] ), .A3(_05521_ ), .ZN(_06039_ ) );
NAND4_X1 _13784_ ( .A1(_05508_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_05512_ ), .A4(_05589_ ), .ZN(_06040_ ) );
NAND4_X1 _13785_ ( .A1(_05508_ ), .A2(_05511_ ), .A3(\mtvec [2] ), .A4(_05512_ ), .ZN(_06041_ ) );
AND3_X1 _13786_ ( .A1(_06039_ ), .A2(_06040_ ), .A3(_06041_ ), .ZN(_06042_ ) );
NAND3_X1 _13787_ ( .A1(_05647_ ), .A2(\mepc [2] ), .A3(_05700_ ), .ZN(_06043_ ) );
AND3_X1 _13788_ ( .A1(_06042_ ), .A2(_05607_ ), .A3(_06043_ ), .ZN(_06044_ ) );
OAI21_X1 _13789_ ( .A(_06038_ ), .B1(_06044_ ), .B2(_05545_ ), .ZN(_06045_ ) );
OR3_X1 _13790_ ( .A1(_04187_ ), .A2(_04188_ ), .A3(_04184_ ), .ZN(_06046_ ) );
AND2_X1 _13791_ ( .A1(_06046_ ), .A2(_04189_ ), .ZN(_06047_ ) );
MUX2_X1 _13792_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B(_06047_ ), .S(_05474_ ), .Z(_06048_ ) );
MUX2_X2 _13793_ ( .A(_06045_ ), .B(_06048_ ), .S(_05481_ ), .Z(_06049_ ) );
NAND2_X1 _13794_ ( .A1(_06049_ ), .A2(_05620_ ), .ZN(_06050_ ) );
XOR2_X1 _13795_ ( .A(_02863_ ), .B(_02887_ ), .Z(_06051_ ) );
AOI22_X1 _13796_ ( .A1(_06051_ ), .A2(_05622_ ), .B1(_04147_ ), .B2(_06047_ ), .ZN(_06052_ ) );
AOI21_X1 _13797_ ( .A(_05978_ ), .B1(_06050_ ), .B2(_06052_ ), .ZN(_00179_ ) );
XOR2_X1 _13798_ ( .A(_04185_ ), .B(_04186_ ), .Z(_06053_ ) );
AOI21_X1 _13799_ ( .A(\ID_EX_typ [3] ), .B1(_05626_ ), .B2(_06053_ ), .ZN(_06054_ ) );
INV_X1 _13800_ ( .A(\ID_EX_pc [1] ), .ZN(_06055_ ) );
OAI21_X1 _13801_ ( .A(_06054_ ), .B1(_06055_ ), .B2(_05633_ ), .ZN(_06056_ ) );
NAND3_X1 _13802_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_05671_ ), .ZN(_06057_ ) );
NAND3_X1 _13803_ ( .A1(_05911_ ), .A2(\mepc [1] ), .A3(_05700_ ), .ZN(_06058_ ) );
NAND3_X1 _13804_ ( .A1(_05911_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_05594_ ), .ZN(_06059_ ) );
BUF_X4 _13805_ ( .A(_05717_ ), .Z(_06060_ ) );
BUF_X4 _13806_ ( .A(_05718_ ), .Z(_06061_ ) );
NAND4_X1 _13807_ ( .A1(_06060_ ), .A2(_05679_ ), .A3(\mtvec [1] ), .A4(_06061_ ), .ZN(_06062_ ) );
BUF_X4 _13808_ ( .A(_05589_ ), .Z(_06063_ ) );
NAND4_X1 _13809_ ( .A1(_06060_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_06061_ ), .A4(_06063_ ), .ZN(_06064_ ) );
AND4_X1 _13810_ ( .A1(_06058_ ), .A2(_06059_ ), .A3(_06062_ ), .A4(_06064_ ), .ZN(_06065_ ) );
OAI21_X1 _13811_ ( .A(_06057_ ), .B1(_06065_ ), .B2(_05682_ ), .ZN(_06066_ ) );
OAI211_X1 _13812_ ( .A(_06056_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06066_ ), .ZN(_06067_ ) );
XOR2_X1 _13813_ ( .A(_02837_ ), .B(_02860_ ), .Z(_06068_ ) );
AOI22_X1 _13814_ ( .A1(_06068_ ), .A2(_05622_ ), .B1(_04147_ ), .B2(_06053_ ), .ZN(_06069_ ) );
AOI21_X1 _13815_ ( .A(_05978_ ), .B1(_06067_ ), .B2(_06069_ ), .ZN(_00180_ ) );
NAND3_X1 _13816_ ( .A1(_05562_ ), .A2(\ID_EX_pc [26] ), .A3(_05565_ ), .ZN(_06070_ ) );
XNOR2_X1 _13817_ ( .A(_06070_ ), .B(\ID_EX_pc [27] ), .ZN(_06071_ ) );
OAI21_X1 _13818_ ( .A(_06071_ ), .B1(_05471_ ), .B2(_05473_ ), .ZN(_06072_ ) );
NAND2_X1 _13819_ ( .A1(_04275_ ), .A2(_04277_ ), .ZN(_06073_ ) );
NAND2_X1 _13820_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_06074_ ) );
NAND2_X1 _13821_ ( .A1(_06073_ ), .A2(_06074_ ), .ZN(_06075_ ) );
XNOR2_X1 _13822_ ( .A(_06075_ ), .B(_04276_ ), .ZN(_06076_ ) );
OAI211_X1 _13823_ ( .A(_05556_ ), .B(_06072_ ), .C1(_05574_ ), .C2(_06076_ ), .ZN(_06077_ ) );
NAND3_X1 _13824_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_05671_ ), .ZN(_06078_ ) );
NAND4_X1 _13825_ ( .A1(_05643_ ), .A2(_05644_ ), .A3(\mtvec [27] ), .A4(_05645_ ), .ZN(_06079_ ) );
AND2_X1 _13826_ ( .A1(_05517_ ), .A2(_06079_ ), .ZN(_06080_ ) );
NAND4_X1 _13827_ ( .A1(_06060_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_06061_ ), .A4(_06063_ ), .ZN(_06081_ ) );
NAND3_X1 _13828_ ( .A1(_05911_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_05594_ ), .ZN(_06082_ ) );
NAND3_X1 _13829_ ( .A1(_05592_ ), .A2(\mepc [27] ), .A3(_05700_ ), .ZN(_06083_ ) );
AND4_X1 _13830_ ( .A1(_06080_ ), .A2(_06081_ ), .A3(_06082_ ), .A4(_06083_ ), .ZN(_06084_ ) );
OAI21_X1 _13831_ ( .A(_06078_ ), .B1(_06084_ ), .B2(_05682_ ), .ZN(_06085_ ) );
OAI211_X1 _13832_ ( .A(_06077_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06085_ ), .ZN(_06086_ ) );
MUX2_X1 _13833_ ( .A(_06076_ ), .B(_03291_ ), .S(fanout_net_7 ), .Z(_06087_ ) );
OR2_X1 _13834_ ( .A1(_06087_ ), .A2(_05601_ ), .ZN(_06088_ ) );
AOI21_X1 _13835_ ( .A(_05978_ ), .B1(_06086_ ), .B2(_06088_ ), .ZN(_00181_ ) );
NAND3_X1 _13836_ ( .A1(_05494_ ), .A2(\mepc [0] ), .A3(_05498_ ), .ZN(_06089_ ) );
NAND4_X1 _13837_ ( .A1(_05500_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_05502_ ), .A4(_05505_ ), .ZN(_06090_ ) );
AND2_X1 _13838_ ( .A1(_06089_ ), .A2(_06090_ ), .ZN(_06091_ ) );
NAND4_X1 _13839_ ( .A1(_05508_ ), .A2(_05511_ ), .A3(\mtvec [0] ), .A4(_05512_ ), .ZN(_06092_ ) );
NAND3_X1 _13840_ ( .A1(_05518_ ), .A2(\mycsreg.CSReg[3][0] ), .A3(_05593_ ), .ZN(_06093_ ) );
NAND4_X1 _13841_ ( .A1(_06091_ ), .A2(_05607_ ), .A3(_06092_ ), .A4(_06093_ ), .ZN(_06094_ ) );
NAND2_X1 _13842_ ( .A1(_06094_ ), .A2(_05546_ ), .ZN(_06095_ ) );
NAND3_X1 _13843_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_05655_ ), .ZN(_06096_ ) );
AND2_X1 _13844_ ( .A1(_06095_ ), .A2(_06096_ ), .ZN(_06097_ ) );
INV_X1 _13845_ ( .A(_06097_ ), .ZN(_06098_ ) );
XOR2_X1 _13846_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_06099_ ) );
MUX2_X1 _13847_ ( .A(\ID_EX_pc [0] ), .B(_06099_ ), .S(_05474_ ), .Z(_06100_ ) );
MUX2_X2 _13848_ ( .A(_06098_ ), .B(_06100_ ), .S(_05481_ ), .Z(_06101_ ) );
AOI22_X1 _13849_ ( .A1(_06101_ ), .A2(_05620_ ), .B1(_05777_ ), .B2(_06099_ ), .ZN(_06102_ ) );
NOR2_X1 _13850_ ( .A1(_06102_ ), .A2(_04159_ ), .ZN(_00182_ ) );
XNOR2_X1 _13851_ ( .A(_05566_ ), .B(\ID_EX_pc [26] ), .ZN(_06103_ ) );
AOI21_X1 _13852_ ( .A(\ID_EX_typ [3] ), .B1(_05574_ ), .B2(_06103_ ), .ZN(_06104_ ) );
XOR2_X1 _13853_ ( .A(_04275_ ), .B(_04277_ ), .Z(_06105_ ) );
INV_X1 _13854_ ( .A(_06105_ ), .ZN(_06106_ ) );
OAI21_X1 _13855_ ( .A(_06104_ ), .B1(_05574_ ), .B2(_06106_ ), .ZN(_06107_ ) );
NAND3_X1 _13856_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_05671_ ), .ZN(_06108_ ) );
NAND3_X1 _13857_ ( .A1(_05911_ ), .A2(\mepc [26] ), .A3(_05700_ ), .ZN(_06109_ ) );
NAND3_X1 _13858_ ( .A1(_05911_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_05594_ ), .ZN(_06110_ ) );
NAND4_X1 _13859_ ( .A1(_06060_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_06061_ ), .A4(_06063_ ), .ZN(_06111_ ) );
NAND4_X1 _13860_ ( .A1(_06060_ ), .A2(_05679_ ), .A3(\mtvec [26] ), .A4(_05645_ ), .ZN(_06112_ ) );
AND4_X1 _13861_ ( .A1(_06109_ ), .A2(_06110_ ), .A3(_06111_ ), .A4(_06112_ ), .ZN(_06113_ ) );
OAI21_X1 _13862_ ( .A(_06108_ ), .B1(_06113_ ), .B2(_05682_ ), .ZN(_06114_ ) );
OAI211_X1 _13863_ ( .A(_06107_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06114_ ), .ZN(_06115_ ) );
NOR4_X1 _13864_ ( .A1(_03289_ ), .A2(_03292_ ), .A3(_05732_ ), .A4(_05600_ ), .ZN(_06116_ ) );
AOI21_X1 _13865_ ( .A(_06116_ ), .B1(_05624_ ), .B2(_06105_ ), .ZN(_06117_ ) );
AOI21_X1 _13866_ ( .A(_05978_ ), .B1(_06115_ ), .B2(_06117_ ), .ZN(_00183_ ) );
AND3_X1 _13867_ ( .A1(_05564_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_06118_ ) );
AND2_X1 _13868_ ( .A1(_05562_ ), .A2(_06118_ ), .ZN(_06119_ ) );
NAND3_X1 _13869_ ( .A1(_06119_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_06120_ ) );
INV_X1 _13870_ ( .A(\ID_EX_pc [24] ), .ZN(_06121_ ) );
NOR2_X1 _13871_ ( .A1(_06120_ ), .A2(_06121_ ), .ZN(_06122_ ) );
INV_X1 _13872_ ( .A(\ID_EX_pc [25] ), .ZN(_06123_ ) );
XNOR2_X1 _13873_ ( .A(_06122_ ), .B(_06123_ ), .ZN(_06124_ ) );
AOI21_X1 _13874_ ( .A(\ID_EX_typ [3] ), .B1(_05574_ ), .B2(_06124_ ), .ZN(_06125_ ) );
OR2_X1 _13875_ ( .A1(_04262_ ), .A2(_04270_ ), .ZN(_06126_ ) );
AND2_X1 _13876_ ( .A1(_06126_ ), .A2(_04181_ ), .ZN(_06127_ ) );
OR2_X1 _13877_ ( .A1(_06127_ ), .A2(_04272_ ), .ZN(_06128_ ) );
XNOR2_X1 _13878_ ( .A(_06128_ ), .B(_04180_ ), .ZN(_06129_ ) );
OAI21_X1 _13879_ ( .A(_06125_ ), .B1(_05574_ ), .B2(_06129_ ), .ZN(_06130_ ) );
NAND3_X1 _13880_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_05671_ ), .ZN(_06131_ ) );
NAND3_X1 _13881_ ( .A1(_05911_ ), .A2(\mepc [25] ), .A3(_05700_ ), .ZN(_06132_ ) );
NAND3_X1 _13882_ ( .A1(_05911_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_05594_ ), .ZN(_06133_ ) );
NAND4_X1 _13883_ ( .A1(_06060_ ), .A2(_05679_ ), .A3(\mtvec [25] ), .A4(_06061_ ), .ZN(_06134_ ) );
NAND4_X1 _13884_ ( .A1(_06060_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_06061_ ), .A4(_06063_ ), .ZN(_06135_ ) );
AND4_X1 _13885_ ( .A1(_06132_ ), .A2(_06133_ ), .A3(_06134_ ), .A4(_06135_ ), .ZN(_06136_ ) );
OAI21_X1 _13886_ ( .A(_06131_ ), .B1(_06136_ ), .B2(_05682_ ), .ZN(_06137_ ) );
OAI211_X1 _13887_ ( .A(_06130_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06137_ ), .ZN(_06138_ ) );
NOR2_X1 _13888_ ( .A1(_06129_ ), .A2(_04148_ ), .ZN(_06139_ ) );
BUF_X4 _13889_ ( .A(_04146_ ), .Z(_06140_ ) );
BUF_X4 _13890_ ( .A(_05600_ ), .Z(_06141_ ) );
NOR3_X1 _13891_ ( .A1(_03294_ ), .A2(_06140_ ), .A3(_06141_ ), .ZN(_06142_ ) );
NOR2_X1 _13892_ ( .A1(_06139_ ), .A2(_06142_ ), .ZN(_06143_ ) );
AOI21_X1 _13893_ ( .A(_05978_ ), .B1(_06138_ ), .B2(_06143_ ), .ZN(_00184_ ) );
XNOR2_X1 _13894_ ( .A(_06120_ ), .B(\ID_EX_pc [24] ), .ZN(_06144_ ) );
AOI21_X1 _13895_ ( .A(\ID_EX_typ [3] ), .B1(_05573_ ), .B2(_06144_ ), .ZN(_06145_ ) );
XOR2_X1 _13896_ ( .A(_06126_ ), .B(_04181_ ), .Z(_06146_ ) );
INV_X1 _13897_ ( .A(_06146_ ), .ZN(_06147_ ) );
OAI21_X1 _13898_ ( .A(_06145_ ), .B1(_05574_ ), .B2(_06147_ ), .ZN(_06148_ ) );
NAND3_X1 _13899_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_05580_ ), .ZN(_06149_ ) );
NAND3_X1 _13900_ ( .A1(_05518_ ), .A2(\mepc [24] ), .A3(_05583_ ), .ZN(_06150_ ) );
NAND4_X1 _13901_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(\mtvec [24] ), .A4(_05587_ ), .ZN(_06151_ ) );
NAND4_X1 _13902_ ( .A1(_05585_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_05587_ ), .A4(_05589_ ), .ZN(_06152_ ) );
AND3_X1 _13903_ ( .A1(_06150_ ), .A2(_06151_ ), .A3(_06152_ ), .ZN(_06153_ ) );
NAND3_X1 _13904_ ( .A1(_05592_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_05648_ ), .ZN(_06154_ ) );
AND3_X1 _13905_ ( .A1(_06153_ ), .A2(_05608_ ), .A3(_06154_ ), .ZN(_06155_ ) );
OAI21_X1 _13906_ ( .A(_06149_ ), .B1(_06155_ ), .B2(_05545_ ), .ZN(_06156_ ) );
OAI211_X1 _13907_ ( .A(_06148_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06156_ ), .ZN(_06157_ ) );
NOR4_X1 _13908_ ( .A1(_03295_ ), .A2(_03160_ ), .A3(_05732_ ), .A4(_05600_ ), .ZN(_06158_ ) );
AOI21_X1 _13909_ ( .A(_06158_ ), .B1(_05624_ ), .B2(_06146_ ), .ZN(_06159_ ) );
AOI21_X1 _13910_ ( .A(_05978_ ), .B1(_06157_ ), .B2(_06159_ ), .ZN(_00185_ ) );
NAND3_X1 _13911_ ( .A1(_05562_ ), .A2(\ID_EX_pc [22] ), .A3(_06118_ ), .ZN(_06160_ ) );
XNOR2_X1 _13912_ ( .A(_06160_ ), .B(\ID_EX_pc [23] ), .ZN(_06161_ ) );
OAI21_X1 _13913_ ( .A(_06161_ ), .B1(_05471_ ), .B2(_05473_ ), .ZN(_06162_ ) );
INV_X1 _13914_ ( .A(_04257_ ), .ZN(_06163_ ) );
OAI21_X1 _13915_ ( .A(_04261_ ), .B1(_04246_ ), .B2(_04254_ ), .ZN(_06164_ ) );
AOI21_X1 _13916_ ( .A(_06163_ ), .B1(_06164_ ), .B2(_04268_ ), .ZN(_06165_ ) );
OR2_X1 _13917_ ( .A1(_06165_ ), .A2(_04263_ ), .ZN(_06166_ ) );
XNOR2_X1 _13918_ ( .A(_06166_ ), .B(_04256_ ), .ZN(_06167_ ) );
OAI211_X1 _13919_ ( .A(_05556_ ), .B(_06162_ ), .C1(_05574_ ), .C2(_06167_ ), .ZN(_06168_ ) );
NAND3_X1 _13920_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_05671_ ), .ZN(_06169_ ) );
NAND3_X1 _13921_ ( .A1(_05911_ ), .A2(\mepc [23] ), .A3(_05700_ ), .ZN(_06170_ ) );
NAND3_X1 _13922_ ( .A1(_05592_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_05594_ ), .ZN(_06171_ ) );
NAND4_X1 _13923_ ( .A1(_06060_ ), .A2(_05679_ ), .A3(\mtvec [23] ), .A4(_06061_ ), .ZN(_06172_ ) );
NAND4_X1 _13924_ ( .A1(_05643_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_06061_ ), .A4(_06063_ ), .ZN(_06173_ ) );
AND4_X1 _13925_ ( .A1(_06170_ ), .A2(_06171_ ), .A3(_06172_ ), .A4(_06173_ ), .ZN(_06174_ ) );
OAI21_X1 _13926_ ( .A(_06169_ ), .B1(_06174_ ), .B2(_05682_ ), .ZN(_06175_ ) );
OAI211_X1 _13927_ ( .A(_06168_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06175_ ), .ZN(_06176_ ) );
MUX2_X1 _13928_ ( .A(_06167_ ), .B(_03302_ ), .S(fanout_net_7 ), .Z(_06177_ ) );
OR2_X1 _13929_ ( .A1(_06177_ ), .A2(_05601_ ), .ZN(_06178_ ) );
AOI21_X1 _13930_ ( .A(_05978_ ), .B1(_06176_ ), .B2(_06178_ ), .ZN(_00186_ ) );
NAND3_X1 _13931_ ( .A1(_05579_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_05580_ ), .ZN(_06179_ ) );
NAND3_X1 _13932_ ( .A1(_05494_ ), .A2(\mepc [22] ), .A3(_05583_ ), .ZN(_06180_ ) );
NAND4_X1 _13933_ ( .A1(_05508_ ), .A2(_05511_ ), .A3(\mtvec [22] ), .A4(_05512_ ), .ZN(_06181_ ) );
NAND4_X1 _13934_ ( .A1(_05508_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_05512_ ), .A4(_05505_ ), .ZN(_06182_ ) );
AND3_X1 _13935_ ( .A1(_06180_ ), .A2(_06181_ ), .A3(_06182_ ), .ZN(_06183_ ) );
NAND3_X1 _13936_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_05648_ ), .ZN(_06184_ ) );
AND3_X1 _13937_ ( .A1(_06183_ ), .A2(_05608_ ), .A3(_06184_ ), .ZN(_06185_ ) );
OAI21_X1 _13938_ ( .A(_06179_ ), .B1(_06185_ ), .B2(_05545_ ), .ZN(_06186_ ) );
INV_X1 _13939_ ( .A(\ID_EX_pc [22] ), .ZN(_06187_ ) );
XNOR2_X1 _13940_ ( .A(_06119_ ), .B(_06187_ ), .ZN(_06188_ ) );
AND3_X1 _13941_ ( .A1(_06164_ ), .A2(_06163_ ), .A3(_04268_ ), .ZN(_06189_ ) );
NOR2_X1 _13942_ ( .A1(_06189_ ), .A2(_06165_ ), .ZN(_06190_ ) );
MUX2_X1 _13943_ ( .A(_06188_ ), .B(_06190_ ), .S(_05474_ ), .Z(_06191_ ) );
MUX2_X2 _13944_ ( .A(_06186_ ), .B(_06191_ ), .S(_05481_ ), .Z(_06192_ ) );
NAND2_X1 _13945_ ( .A1(_06192_ ), .A2(_05620_ ), .ZN(_06193_ ) );
AOI22_X1 _13946_ ( .A1(_03303_ ), .A2(_05622_ ), .B1(_04147_ ), .B2(_06190_ ), .ZN(_06194_ ) );
AOI21_X1 _13947_ ( .A(_04142_ ), .B1(_06193_ ), .B2(_06194_ ), .ZN(_00187_ ) );
INV_X1 _13948_ ( .A(\ID_EX_pc [20] ), .ZN(_06195_ ) );
NOR2_X1 _13949_ ( .A1(_05615_ ), .A2(_06195_ ), .ZN(_06196_ ) );
INV_X1 _13950_ ( .A(\ID_EX_pc [21] ), .ZN(_06197_ ) );
XNOR2_X1 _13951_ ( .A(_06196_ ), .B(_06197_ ), .ZN(_06198_ ) );
AOI21_X1 _13952_ ( .A(\ID_EX_typ [3] ), .B1(_05573_ ), .B2(_06198_ ), .ZN(_06199_ ) );
AND2_X1 _13953_ ( .A1(_04255_ ), .A2(_04260_ ), .ZN(_06200_ ) );
OR2_X1 _13954_ ( .A1(_06200_ ), .A2(_04266_ ), .ZN(_06201_ ) );
XNOR2_X1 _13955_ ( .A(_06201_ ), .B(_04259_ ), .ZN(_06202_ ) );
OAI21_X1 _13956_ ( .A(_06199_ ), .B1(_05574_ ), .B2(_06202_ ), .ZN(_06203_ ) );
NAND3_X1 _13957_ ( .A1(_05647_ ), .A2(\mepc [21] ), .A3(_05605_ ), .ZN(_06204_ ) );
NAND4_X1 _13958_ ( .A1(_05717_ ), .A2(_05678_ ), .A3(\mtvec [21] ), .A4(_05640_ ), .ZN(_06205_ ) );
NAND4_X1 _13959_ ( .A1(_05639_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_05718_ ), .A4(_05675_ ), .ZN(_06206_ ) );
NAND3_X1 _13960_ ( .A1(_06204_ ), .A2(_06205_ ), .A3(_06206_ ), .ZN(_06207_ ) );
NAND3_X1 _13961_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_05648_ ), .ZN(_06208_ ) );
NAND2_X1 _13962_ ( .A1(_06208_ ), .A2(_05517_ ), .ZN(_06209_ ) );
OAI21_X1 _13963_ ( .A(_05651_ ), .B1(_06207_ ), .B2(_06209_ ), .ZN(_06210_ ) );
NAND3_X1 _13964_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [21] ), .A3(_05655_ ), .ZN(_06211_ ) );
AND2_X1 _13965_ ( .A1(_06210_ ), .A2(_06211_ ), .ZN(_06212_ ) );
INV_X1 _13966_ ( .A(_06212_ ), .ZN(_06213_ ) );
OAI211_X1 _13967_ ( .A(_06203_ ), .B(_05712_ ), .C1(_05713_ ), .C2(_06213_ ), .ZN(_06214_ ) );
BUF_X4 _13968_ ( .A(_04146_ ), .Z(_06215_ ) );
NOR3_X1 _13969_ ( .A1(_03254_ ), .A2(_06215_ ), .A3(_06141_ ), .ZN(_06216_ ) );
NOR2_X1 _13970_ ( .A1(_06202_ ), .A2(_04148_ ), .ZN(_06217_ ) );
NOR2_X1 _13971_ ( .A1(_06216_ ), .A2(_06217_ ), .ZN(_06218_ ) );
AOI21_X1 _13972_ ( .A(_04142_ ), .B1(_06214_ ), .B2(_06218_ ), .ZN(_00188_ ) );
OAI21_X1 _13973_ ( .A(_04289_ ), .B1(_04286_ ), .B2(_04287_ ), .ZN(_06219_ ) );
NAND2_X1 _13974_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_06220_ ) );
AND2_X1 _13975_ ( .A1(_06219_ ), .A2(_06220_ ), .ZN(_06221_ ) );
XNOR2_X1 _13976_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_06222_ ) );
XNOR2_X1 _13977_ ( .A(_06221_ ), .B(_06222_ ), .ZN(_06223_ ) );
MUX2_X1 _13978_ ( .A(_06223_ ), .B(_03245_ ), .S(fanout_net_7 ), .Z(_06224_ ) );
OR2_X1 _13979_ ( .A1(_06224_ ), .A2(_06141_ ), .ZN(_06225_ ) );
OR3_X1 _13980_ ( .A1(_05844_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_05846_ ), .ZN(_06226_ ) );
NAND3_X1 _13981_ ( .A1(_05856_ ), .A2(\mtvec [31] ), .A3(_05678_ ), .ZN(_06227_ ) );
NAND3_X1 _13982_ ( .A1(_05856_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_05675_ ), .ZN(_06228_ ) );
AND2_X1 _13983_ ( .A1(_06227_ ), .A2(_06228_ ), .ZN(_06229_ ) );
NAND3_X1 _13984_ ( .A1(_05592_ ), .A2(\mepc [31] ), .A3(_05700_ ), .ZN(_06230_ ) );
NAND3_X1 _13985_ ( .A1(_05592_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_05594_ ), .ZN(_06231_ ) );
NAND3_X1 _13986_ ( .A1(_06229_ ), .A2(_06230_ ), .A3(_06231_ ), .ZN(_06232_ ) );
NOR2_X1 _13987_ ( .A1(_05844_ ), .A2(_05846_ ), .ZN(_06233_ ) );
OAI21_X1 _13988_ ( .A(_06226_ ), .B1(_06232_ ), .B2(_06233_ ), .ZN(_06234_ ) );
INV_X1 _13989_ ( .A(\ID_EX_pc [30] ), .ZN(_06235_ ) );
NOR2_X1 _13990_ ( .A1(_04178_ ), .A2(_06235_ ), .ZN(_06236_ ) );
XNOR2_X1 _13991_ ( .A(_06236_ ), .B(\ID_EX_pc [31] ), .ZN(_06237_ ) );
MUX2_X1 _13992_ ( .A(_06237_ ), .B(_06223_ ), .S(_05475_ ), .Z(_06238_ ) );
MUX2_X2 _13993_ ( .A(_06234_ ), .B(_06238_ ), .S(_05482_ ), .Z(_06239_ ) );
OAI211_X1 _13994_ ( .A(_04158_ ), .B(_06225_ ), .C1(_06239_ ), .C2(_05553_ ), .ZN(_00189_ ) );
INV_X1 _13995_ ( .A(\ID_EX_pc [31] ), .ZN(_06240_ ) );
NOR3_X1 _13996_ ( .A1(_06240_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00190_ ) );
NOR3_X1 _13997_ ( .A1(_06235_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00191_ ) );
NOR3_X1 _13998_ ( .A1(_06197_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00192_ ) );
NOR3_X1 _13999_ ( .A1(_06195_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00193_ ) );
NOR3_X1 _14000_ ( .A1(_05635_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00194_ ) );
NOR3_X1 _14001_ ( .A1(_05664_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00195_ ) );
INV_X1 _14002_ ( .A(\ID_EX_pc [17] ), .ZN(_06241_ ) );
NOR3_X1 _14003_ ( .A1(_06241_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00196_ ) );
NOR3_X1 _14004_ ( .A1(_05693_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00197_ ) );
INV_X1 _14005_ ( .A(\ID_EX_pc [15] ), .ZN(_06242_ ) );
NOR3_X1 _14006_ ( .A1(_06242_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00198_ ) );
NOR3_X1 _14007_ ( .A1(_05769_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00199_ ) );
NOR3_X1 _14008_ ( .A1(_05559_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00200_ ) );
NOR3_X1 _14009_ ( .A1(_05560_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00201_ ) );
NOR3_X1 _14010_ ( .A1(_04285_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00202_ ) );
INV_X1 _14011_ ( .A(\ID_EX_pc [11] ), .ZN(_06243_ ) );
NOR3_X1 _14012_ ( .A1(_06243_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00203_ ) );
NOR3_X1 _14013_ ( .A1(_05890_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00204_ ) );
NOR3_X1 _14014_ ( .A1(_05899_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00205_ ) );
INV_X1 _14015_ ( .A(\ID_EX_pc [8] ), .ZN(_06244_ ) );
NOR3_X1 _14016_ ( .A1(_06244_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00206_ ) );
NOR3_X1 _14017_ ( .A1(_05944_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00207_ ) );
NOR3_X1 _14018_ ( .A1(_05958_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00208_ ) );
AND2_X1 _14019_ ( .A1(_04158_ ), .A2(\ID_EX_pc [5] ), .ZN(_00209_ ) );
INV_X1 _14020_ ( .A(\ID_EX_pc [4] ), .ZN(_06245_ ) );
NOR3_X1 _14021_ ( .A1(_06245_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00210_ ) );
NOR3_X1 _14022_ ( .A1(_04191_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00211_ ) );
INV_X1 _14023_ ( .A(\ID_EX_pc [2] ), .ZN(_06246_ ) );
NOR3_X1 _14024_ ( .A1(_06246_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00212_ ) );
NOR3_X1 _14025_ ( .A1(_05839_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00213_ ) );
NOR3_X1 _14026_ ( .A1(_06055_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00214_ ) );
AND2_X1 _14027_ ( .A1(_04158_ ), .A2(\ID_EX_pc [0] ), .ZN(_00215_ ) );
NOR3_X1 _14028_ ( .A1(_05567_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00216_ ) );
NOR3_X1 _14029_ ( .A1(_05568_ ), .A2(fanout_net_5 ), .A3(fanout_net_17 ), .ZN(_00217_ ) );
NOR3_X1 _14030_ ( .A1(_06123_ ), .A2(reset ), .A3(fanout_net_17 ), .ZN(_00218_ ) );
NOR3_X1 _14031_ ( .A1(_06121_ ), .A2(reset ), .A3(fanout_net_17 ), .ZN(_00219_ ) );
INV_X1 _14032_ ( .A(\ID_EX_pc [23] ), .ZN(_06247_ ) );
NOR3_X1 _14033_ ( .A1(_06247_ ), .A2(reset ), .A3(fanout_net_17 ), .ZN(_00220_ ) );
NOR3_X1 _14034_ ( .A1(_06187_ ), .A2(reset ), .A3(excp_written ), .ZN(_00221_ ) );
NOR3_X1 _14035_ ( .A1(_03605_ ), .A2(reset ), .A3(excp_written ), .ZN(_00222_ ) );
INV_X1 _14036_ ( .A(io_master_awready ), .ZN(_06248_ ) );
NAND3_X1 _14037_ ( .A1(_02255_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A3(_06248_ ), .ZN(_06249_ ) );
OAI21_X1 _14038_ ( .A(_06249_ ), .B1(\mylsu.state [4] ), .B2(\mylsu.state [0] ), .ZN(_06250_ ) );
NAND4_X1 _14039_ ( .A1(_02170_ ), .A2(_02184_ ), .A3(\myclint.rvalid ), .A4(_02224_ ), .ZN(_06251_ ) );
AND4_X1 _14040_ ( .A1(_02193_ ), .A2(_02211_ ), .A3(_02201_ ), .A4(_02219_ ), .ZN(_06252_ ) );
NAND2_X1 _14041_ ( .A1(_04074_ ), .A2(_06252_ ), .ZN(_06253_ ) );
AND4_X1 _14042_ ( .A1(_02158_ ), .A2(_02174_ ), .A3(_02162_ ), .A4(_02178_ ), .ZN(_06254_ ) );
AND4_X1 _14043_ ( .A1(_02197_ ), .A2(_02215_ ), .A3(_02206_ ), .A4(\io_master_araddr [25] ), .ZN(_06255_ ) );
NAND2_X1 _14044_ ( .A1(_06254_ ), .A2(_06255_ ), .ZN(_06256_ ) );
NOR2_X1 _14045_ ( .A1(_06253_ ), .A2(_06256_ ), .ZN(_06257_ ) );
OAI21_X1 _14046_ ( .A(_06251_ ), .B1(_06257_ ), .B2(io_master_arready ), .ZN(_06258_ ) );
INV_X1 _14047_ ( .A(_02220_ ), .ZN(_06259_ ) );
BUF_X4 _14048_ ( .A(_06259_ ), .Z(_06260_ ) );
OR2_X1 _14049_ ( .A1(_06258_ ), .A2(_06260_ ), .ZN(_06261_ ) );
AOI21_X1 _14050_ ( .A(_06250_ ), .B1(_06261_ ), .B2(_04112_ ), .ZN(_06262_ ) );
AND2_X1 _14051_ ( .A1(_03320_ ), .A2(EXU_valid_LSU ), .ZN(_06263_ ) );
INV_X1 _14052_ ( .A(_06263_ ), .ZN(_06264_ ) );
OAI22_X1 _14053_ ( .A1(_06262_ ), .A2(_06264_ ), .B1(_04142_ ), .B2(_04143_ ), .ZN(_00223_ ) );
NOR3_X1 _14054_ ( .A1(_04155_ ), .A2(reset ), .A3(excp_written ), .ZN(_00224_ ) );
NOR3_X1 _14055_ ( .A1(_04150_ ), .A2(reset ), .A3(excp_written ), .ZN(_00225_ ) );
NOR3_X1 _14056_ ( .A1(_05144_ ), .A2(reset ), .A3(excp_written ), .ZN(_00226_ ) );
NOR3_X1 _14057_ ( .A1(_05483_ ), .A2(reset ), .A3(excp_written ), .ZN(_00227_ ) );
BUF_X4 _14058_ ( .A(_05127_ ), .Z(_06265_ ) );
BUF_X4 _14059_ ( .A(_06265_ ), .Z(_06266_ ) );
NOR3_X1 _14060_ ( .A1(_06266_ ), .A2(reset ), .A3(excp_written ), .ZN(_00228_ ) );
NOR3_X1 _14061_ ( .A1(_05125_ ), .A2(reset ), .A3(excp_written ), .ZN(_00229_ ) );
NOR3_X1 _14062_ ( .A1(_06215_ ), .A2(reset ), .A3(excp_written ), .ZN(_00230_ ) );
AND2_X1 _14063_ ( .A1(_02268_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_06267_ ) );
CLKBUF_X2 _14064_ ( .A(_06267_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _14065_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .ZN(_06268_ ) );
BUF_X2 _14066_ ( .A(_06268_ ), .Z(_06269_ ) );
AND3_X1 _14067_ ( .A1(_02268_ ), .A2(_06269_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00278_ ) );
AND3_X1 _14068_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_04014_ ), .A3(fanout_net_9 ), .ZN(_00279_ ) );
AND3_X1 _14069_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_13 ), .A3(_04021_ ), .ZN(_00280_ ) );
INV_X1 _14070_ ( .A(\EX_LS_pc [2] ), .ZN(_06270_ ) );
NOR3_X1 _14071_ ( .A1(_06270_ ), .A2(reset ), .A3(excp_written ), .ZN(_00318_ ) );
INV_X1 _14072_ ( .A(\mylsu.state [3] ), .ZN(_06271_ ) );
BUF_X2 _14073_ ( .A(_06271_ ), .Z(_06272_ ) );
BUF_X4 _14074_ ( .A(_06272_ ), .Z(_06273_ ) );
NOR3_X1 _14075_ ( .A1(_06273_ ), .A2(reset ), .A3(excp_written ), .ZN(_00319_ ) );
NOR2_X1 _14076_ ( .A1(\mylsu.state [3] ), .A2(\mylsu.state [1] ), .ZN(_06274_ ) );
AND2_X1 _14077_ ( .A1(_03338_ ), .A2(_06274_ ), .ZN(_06275_ ) );
INV_X1 _14078_ ( .A(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06276_ ) );
NAND2_X1 _14079_ ( .A1(_06275_ ), .A2(_06276_ ), .ZN(_06277_ ) );
INV_X1 _14080_ ( .A(_02253_ ), .ZN(_06278_ ) );
BUF_X4 _14081_ ( .A(_04101_ ), .Z(_06279_ ) );
NOR2_X1 _14082_ ( .A1(_06278_ ), .A2(_06279_ ), .ZN(_06280_ ) );
OAI21_X1 _14083_ ( .A(_02254_ ), .B1(_02318_ ), .B2(_02319_ ), .ZN(_06281_ ) );
OR2_X1 _14084_ ( .A1(_06281_ ), .A2(_02322_ ), .ZN(_06282_ ) );
AOI21_X1 _14085_ ( .A(_04109_ ), .B1(_06282_ ), .B2(\EX_LS_flag [2] ), .ZN(_06283_ ) );
AOI21_X1 _14086_ ( .A(_06277_ ), .B1(_06280_ ), .B2(_06283_ ), .ZN(_00332_ ) );
NOR2_X1 _14087_ ( .A1(_02255_ ), .A2(_02145_ ), .ZN(_06284_ ) );
AOI21_X1 _14088_ ( .A(_06278_ ), .B1(_06282_ ), .B2(_06284_ ), .ZN(_06285_ ) );
AOI21_X1 _14089_ ( .A(_06277_ ), .B1(_06285_ ), .B2(_04113_ ), .ZN(_00333_ ) );
NAND3_X1 _14090_ ( .A1(_02323_ ), .A2(\EX_LS_flag [2] ), .A3(_02243_ ), .ZN(_06286_ ) );
NOR2_X1 _14091_ ( .A1(_06286_ ), .A2(_06277_ ), .ZN(_00334_ ) );
AOI21_X1 _14092_ ( .A(_06277_ ), .B1(_04103_ ), .B2(_02253_ ), .ZN(_00335_ ) );
AOI21_X1 _14093_ ( .A(_06277_ ), .B1(_04113_ ), .B2(_06286_ ), .ZN(_00336_ ) );
INV_X1 _14094_ ( .A(_02264_ ), .ZN(_06287_ ) );
INV_X1 _14095_ ( .A(_02247_ ), .ZN(_06288_ ) );
AND2_X1 _14096_ ( .A1(_06288_ ), .A2(_02252_ ), .ZN(_06289_ ) );
AND3_X1 _14097_ ( .A1(_06281_ ), .A2(_02321_ ), .A3(_06284_ ), .ZN(_06290_ ) );
OR3_X1 _14098_ ( .A1(_06289_ ), .A2(_02257_ ), .A3(_06290_ ), .ZN(_06291_ ) );
INV_X1 _14099_ ( .A(_04109_ ), .ZN(_06292_ ) );
AND3_X1 _14100_ ( .A1(_03338_ ), .A2(_06274_ ), .A3(EXU_valid_LSU ), .ZN(_06293_ ) );
AND4_X1 _14101_ ( .A1(_06287_ ), .A2(_06291_ ), .A3(_06292_ ), .A4(_06293_ ), .ZN(_00337_ ) );
INV_X1 _14102_ ( .A(_00319_ ), .ZN(_06294_ ) );
BUF_X4 _14103_ ( .A(_04105_ ), .Z(_06295_ ) );
OAI21_X1 _14104_ ( .A(_06293_ ), .B1(_06295_ ), .B2(_02374_ ), .ZN(_06296_ ) );
OAI21_X1 _14105_ ( .A(_06294_ ), .B1(_02257_ ), .B2(_06296_ ), .ZN(_00338_ ) );
CLKBUF_X2 _14106_ ( .A(_02232_ ), .Z(_06297_ ) );
CLKBUF_X2 _14107_ ( .A(_06297_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _14108_ ( .A(_02186_ ), .Z(_06298_ ) );
NOR3_X1 _14109_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(_04156_ ), .ZN(_06299_ ) );
BUF_X4 _14110_ ( .A(_06260_ ), .Z(_06300_ ) );
BUF_X4 _14111_ ( .A(_06300_ ), .Z(_06301_ ) );
BUF_X4 _14112_ ( .A(_06301_ ), .Z(_06302_ ) );
INV_X1 _14113_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06303_ ) );
BUF_X4 _14114_ ( .A(_02189_ ), .Z(_06304_ ) );
INV_X1 _14115_ ( .A(_06304_ ), .ZN(_06305_ ) );
AOI211_X1 _14116_ ( .A(_06299_ ), .B(_06302_ ), .C1(_06303_ ), .C2(_06305_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _14117_ ( .A1(_06298_ ), .A2(fanout_net_6 ), .A3(_04156_ ), .ZN(_06306_ ) );
INV_X1 _14118_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06307_ ) );
AOI211_X1 _14119_ ( .A(_06306_ ), .B(_06301_ ), .C1(_06307_ ), .C2(_06305_ ), .ZN(\io_master_araddr [0] ) );
OR3_X1 _14120_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(_04156_ ), .ZN(_06308_ ) );
OAI21_X1 _14121_ ( .A(_06308_ ), .B1(_06304_ ), .B2(\mylsu.araddr_tmp [15] ), .ZN(_06309_ ) );
BUF_X4 _14122_ ( .A(_02167_ ), .Z(_06310_ ) );
BUF_X4 _14123_ ( .A(_06310_ ), .Z(_06311_ ) );
BUF_X4 _14124_ ( .A(_06311_ ), .Z(_06312_ ) );
OAI22_X1 _14125_ ( .A1(_06302_ ), .A2(_06309_ ), .B1(_01993_ ), .B2(_06312_ ), .ZN(\io_master_araddr [15] ) );
AND2_X2 _14126_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ) );
AND4_X1 _14127_ ( .A1(\EX_LS_dest_csreg_mem [14] ), .A2(_02243_ ), .A3(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .A4(_02145_ ), .ZN(_06313_ ) );
AOI21_X1 _14128_ ( .A(_06313_ ), .B1(_06305_ ), .B2(\mylsu.araddr_tmp [14] ), .ZN(_06314_ ) );
OAI22_X1 _14129_ ( .A1(_06302_ ), .A2(_06314_ ), .B1(_02024_ ), .B2(_06312_ ), .ZN(\io_master_araddr [14] ) );
OR3_X1 _14130_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(_04156_ ), .ZN(_06315_ ) );
OAI21_X1 _14131_ ( .A(_06315_ ), .B1(_06304_ ), .B2(\mylsu.araddr_tmp [5] ), .ZN(_06316_ ) );
OAI22_X1 _14132_ ( .A1(_06302_ ), .A2(_06316_ ), .B1(_03782_ ), .B2(_06312_ ), .ZN(\io_master_araddr [5] ) );
OR3_X1 _14133_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(_04156_ ), .ZN(_06317_ ) );
OAI21_X1 _14134_ ( .A(_06317_ ), .B1(_06304_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_06318_ ) );
OAI22_X1 _14135_ ( .A1(_06302_ ), .A2(_06318_ ), .B1(_04014_ ), .B2(_06312_ ), .ZN(\io_master_araddr [4] ) );
OAI221_X1 _14136_ ( .A(fanout_net_9 ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_06319_ ) );
OR3_X1 _14137_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(_04156_ ), .ZN(_06320_ ) );
OAI211_X1 _14138_ ( .A(_02202_ ), .B(_06320_ ), .C1(\mylsu.araddr_tmp [3] ), .C2(_06304_ ), .ZN(_06321_ ) );
OAI21_X1 _14139_ ( .A(_06319_ ), .B1(\io_master_arburst [0] ), .B2(_06321_ ), .ZN(\io_master_araddr [3] ) );
INV_X1 _14140_ ( .A(_02193_ ), .ZN(\io_master_araddr [31] ) );
INV_X1 _14141_ ( .A(_02206_ ), .ZN(\io_master_araddr [30] ) );
INV_X1 _14142_ ( .A(_02197_ ), .ZN(\io_master_araddr [29] ) );
INV_X1 _14143_ ( .A(_02201_ ), .ZN(\io_master_araddr [28] ) );
INV_X1 _14144_ ( .A(_02215_ ), .ZN(\io_master_araddr [27] ) );
INV_X1 _14145_ ( .A(_02219_ ), .ZN(\io_master_araddr [26] ) );
INV_X1 _14146_ ( .A(_02211_ ), .ZN(\io_master_araddr [24] ) );
AND4_X1 _14147_ ( .A1(\EX_LS_dest_csreg_mem [13] ), .A2(_02243_ ), .A3(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .A4(_02145_ ), .ZN(_06322_ ) );
AOI21_X1 _14148_ ( .A(_06322_ ), .B1(_06305_ ), .B2(\mylsu.araddr_tmp [13] ), .ZN(_06323_ ) );
OAI22_X1 _14149_ ( .A1(_06302_ ), .A2(_06323_ ), .B1(_03743_ ), .B2(_06312_ ), .ZN(\io_master_araddr [13] ) );
NOR2_X1 _14150_ ( .A1(_02189_ ), .A2(\mylsu.araddr_tmp [12] ), .ZN(_06324_ ) );
NOR3_X1 _14151_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(_02187_ ), .ZN(_06325_ ) );
NOR3_X1 _14152_ ( .A1(_02150_ ), .A2(_06324_ ), .A3(_06325_ ), .ZN(_06326_ ) );
MUX2_X1 _14153_ ( .A(_06326_ ), .B(\IF_ID_pc [12] ), .S(_06297_ ), .Z(\io_master_araddr [12] ) );
OR3_X1 _14154_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [11] ), .A3(_04156_ ), .ZN(_06327_ ) );
OAI21_X1 _14155_ ( .A(_06327_ ), .B1(_06304_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_06328_ ) );
OAI22_X1 _14156_ ( .A1(_06302_ ), .A2(_06328_ ), .B1(_02092_ ), .B2(_06312_ ), .ZN(\io_master_araddr [11] ) );
OAI221_X1 _14157_ ( .A(\IF_ID_pc [10] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02156_ ), .C2(_02191_ ), .ZN(_06329_ ) );
OR3_X1 _14158_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(_02187_ ), .ZN(_06330_ ) );
OAI211_X1 _14159_ ( .A(_02202_ ), .B(_06330_ ), .C1(\mylsu.araddr_tmp [10] ), .C2(_06304_ ), .ZN(_06331_ ) );
OAI21_X1 _14160_ ( .A(_06329_ ), .B1(\io_master_arburst [0] ), .B2(_06331_ ), .ZN(\io_master_araddr [10] ) );
NAND4_X1 _14161_ ( .A1(_02243_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .A3(_05537_ ), .A4(_04117_ ), .ZN(_06332_ ) );
OAI21_X1 _14162_ ( .A(_06332_ ), .B1(_06304_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06333_ ) );
OAI22_X1 _14163_ ( .A1(_06302_ ), .A2(_06333_ ), .B1(_01960_ ), .B2(_06312_ ), .ZN(\io_master_araddr [9] ) );
NAND4_X1 _14164_ ( .A1(_02243_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .A3(_05538_ ), .A4(_04117_ ), .ZN(_06334_ ) );
OAI21_X1 _14165_ ( .A(_06334_ ), .B1(_06304_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_06335_ ) );
OAI22_X1 _14166_ ( .A1(_06302_ ), .A2(_06335_ ), .B1(_01983_ ), .B2(_06312_ ), .ZN(\io_master_araddr [8] ) );
NOR2_X1 _14167_ ( .A1(_02189_ ), .A2(\mylsu.araddr_tmp [7] ), .ZN(_06336_ ) );
NOR3_X1 _14168_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(_02187_ ), .ZN(_06337_ ) );
NOR3_X1 _14169_ ( .A1(_02150_ ), .A2(_06336_ ), .A3(_06337_ ), .ZN(_06338_ ) );
MUX2_X1 _14170_ ( .A(_06338_ ), .B(\IF_ID_pc [7] ), .S(_06297_ ), .Z(\io_master_araddr [7] ) );
OR3_X1 _14171_ ( .A1(_06298_ ), .A2(\EX_LS_dest_csreg_mem [6] ), .A3(_04156_ ), .ZN(_06339_ ) );
OAI21_X1 _14172_ ( .A(_06339_ ), .B1(_06304_ ), .B2(\mylsu.araddr_tmp [6] ), .ZN(_06340_ ) );
OAI22_X1 _14173_ ( .A1(_06302_ ), .A2(_06340_ ), .B1(_02133_ ), .B2(_06312_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _14174_ ( .A1(_02186_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(_02187_ ), .ZN(_06341_ ) );
OAI211_X1 _14175_ ( .A(_02202_ ), .B(_06341_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_02189_ ), .ZN(_06342_ ) );
NOR2_X1 _14176_ ( .A1(_02205_ ), .A2(_06342_ ), .ZN(_06343_ ) );
BUF_X4 _14177_ ( .A(_06343_ ), .Z(_06344_ ) );
BUF_X2 _14178_ ( .A(_06344_ ), .Z(\io_master_araddr [2] ) );
BUF_X2 _14179_ ( .A(_02220_ ), .Z(\io_master_arid [1] ) );
BUF_X2 _14180_ ( .A(_06310_ ), .Z(_06345_ ) );
AND3_X1 _14181_ ( .A1(_06345_ ), .A2(\EX_LS_typ [3] ), .A3(_02202_ ), .ZN(\io_master_arsize [2] ) );
AND3_X1 _14182_ ( .A1(_06345_ ), .A2(\EX_LS_typ [1] ), .A3(_02202_ ), .ZN(\io_master_arsize [0] ) );
OAI22_X1 _14183_ ( .A1(_02142_ ), .A2(_02143_ ), .B1(_02235_ ), .B2(_02150_ ), .ZN(\io_master_arsize [1] ) );
NOR3_X1 _14184_ ( .A1(_04080_ ), .A2(_02273_ ), .A3(_02274_ ), .ZN(io_master_arvalid ) );
AND2_X1 _14185_ ( .A1(_02256_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_06346_ ) );
BUF_X4 _14186_ ( .A(_06346_ ), .Z(_06347_ ) );
BUF_X4 _14187_ ( .A(_06347_ ), .Z(_06348_ ) );
MUX2_X1 _14188_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06348_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _14189_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06348_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _14190_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06348_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _14191_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06348_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _14192_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06348_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _14193_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06348_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _14194_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06348_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _14195_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06348_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _14196_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06348_ ), .Z(\io_master_awaddr [15] ) );
BUF_X4 _14197_ ( .A(_06347_ ), .Z(_06349_ ) );
MUX2_X1 _14198_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06349_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _14199_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06349_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _14200_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06349_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _14201_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06349_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _14202_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06349_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _14203_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06349_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _14204_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06349_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _14205_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06349_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _14206_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06349_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _14207_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06349_ ), .Z(\io_master_awaddr [6] ) );
BUF_X4 _14208_ ( .A(_06347_ ), .Z(_06350_ ) );
MUX2_X1 _14209_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06350_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _14210_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06350_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _14211_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06350_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _14212_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06350_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _14213_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06350_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _14214_ ( .A(\mylsu.awaddr_tmp [1] ), .B(\EX_LS_dest_csreg_mem [1] ), .S(_06350_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _14215_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_6 ), .S(_06350_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _14216_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06350_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _14217_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06350_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _14218_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06350_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _14219_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06347_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _14220_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06347_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _14221_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06347_ ), .Z(\io_master_awaddr [22] ) );
AND3_X1 _14222_ ( .A1(_02259_ ), .A2(\EX_LS_typ [1] ), .A3(_02238_ ), .ZN(\io_master_awsize [0] ) );
NAND2_X1 _14223_ ( .A1(_02259_ ), .A2(_02238_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _14224_ ( .A1(_02253_ ), .A2(_02265_ ), .A3(_06348_ ), .ZN(_06351_ ) );
INV_X1 _14225_ ( .A(\mylsu.state [4] ), .ZN(_06352_ ) );
NAND2_X1 _14226_ ( .A1(_06351_ ), .A2(_06352_ ), .ZN(io_master_awvalid ) );
INV_X1 _14227_ ( .A(\mylsu.state [2] ), .ZN(_06353_ ) );
INV_X1 _14228_ ( .A(\mylsu.state [1] ), .ZN(_06354_ ) );
NAND4_X1 _14229_ ( .A1(_06351_ ), .A2(_06353_ ), .A3(_06352_ ), .A4(_06354_ ), .ZN(io_master_bready ) );
NOR2_X1 _14230_ ( .A1(_04084_ ), .A2(\io_master_rid [0] ), .ZN(_06355_ ) );
NAND4_X1 _14231_ ( .A1(_06355_ ), .A2(io_master_rlast ), .A3(_04082_ ), .A4(_04083_ ), .ZN(_06356_ ) );
AOI21_X1 _14232_ ( .A(_06260_ ), .B1(_04081_ ), .B2(_06356_ ), .ZN(_06357_ ) );
AOI21_X1 _14233_ ( .A(_06273_ ), .B1(_06357_ ), .B2(_04089_ ), .ZN(_06358_ ) );
NOR3_X1 _14234_ ( .A1(_02149_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_06359_ ) );
NAND2_X1 _14235_ ( .A1(\io_master_bid [1] ), .A2(\io_master_bid [0] ), .ZN(_06360_ ) );
OR3_X1 _14236_ ( .A1(_06360_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bid [2] ), .ZN(_06361_ ) );
NOR2_X1 _14237_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_06362_ ) );
NAND2_X1 _14238_ ( .A1(_06362_ ), .A2(io_master_bvalid ), .ZN(_06363_ ) );
NOR2_X1 _14239_ ( .A1(_06361_ ), .A2(_06363_ ), .ZN(_06364_ ) );
NOR2_X1 _14240_ ( .A1(_06364_ ), .A2(_06354_ ), .ZN(_06365_ ) );
NOR3_X1 _14241_ ( .A1(_06358_ ), .A2(_06359_ ), .A3(_06365_ ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
NOR3_X1 _14242_ ( .A1(_04080_ ), .A2(_02267_ ), .A3(_02270_ ), .ZN(io_master_rready ) );
MUX2_X1 _14243_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_6 ), .Z(_06366_ ) );
INV_X1 _14244_ ( .A(\EX_LS_dest_csreg_mem [1] ), .ZN(_06367_ ) );
CLKBUF_X2 _14245_ ( .A(_06367_ ), .Z(_06368_ ) );
AND2_X1 _14246_ ( .A1(_06366_ ), .A2(_06368_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _14247_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_6 ), .Z(_06369_ ) );
AND2_X1 _14248_ ( .A1(_06369_ ), .A2(_06368_ ), .ZN(\io_master_wdata [14] ) );
INV_X1 _14249_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_06370_ ) );
NOR3_X1 _14250_ ( .A1(_06370_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [5] ) );
INV_X1 _14251_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_06371_ ) );
NOR3_X1 _14252_ ( .A1(_06371_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [4] ) );
INV_X1 _14253_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_06372_ ) );
NOR3_X1 _14254_ ( .A1(_06372_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14255_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_06373_ ) );
NOR3_X1 _14256_ ( .A1(_06373_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14257_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06374_ ) );
NOR3_X1 _14258_ ( .A1(_06374_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14259_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06375_ ) );
NOR3_X1 _14260_ ( .A1(_06375_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14261_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_6 ), .Z(_06376_ ) );
AND2_X1 _14262_ ( .A1(_06376_ ), .A2(_06368_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14263_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_6 ), .Z(_06377_ ) );
AND2_X1 _14264_ ( .A1(_06377_ ), .A2(_06368_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14265_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_6 ), .Z(_06378_ ) );
AND2_X1 _14266_ ( .A1(_06378_ ), .A2(_06368_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14267_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_6 ), .Z(_06379_ ) );
AND2_X1 _14268_ ( .A1(_06379_ ), .A2(_06368_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14269_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_6 ), .Z(_06380_ ) );
AND2_X1 _14270_ ( .A1(_06380_ ), .A2(_06368_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14271_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_6 ), .Z(_06381_ ) );
AND2_X1 _14272_ ( .A1(_06381_ ), .A2(_06368_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14273_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06382_ ) );
NOR3_X1 _14274_ ( .A1(_06382_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [7] ) );
INV_X1 _14275_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_06383_ ) );
NOR3_X1 _14276_ ( .A1(_06383_ ), .A2(fanout_net_6 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14277_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_6 ), .Z(_06384_ ) );
MUX2_X1 _14278_ ( .A(_06384_ ), .B(_06366_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14279_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_6 ), .Z(_06385_ ) );
MUX2_X1 _14280_ ( .A(_06385_ ), .B(_06369_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [30] ) );
NOR2_X1 _14281_ ( .A1(_06367_ ), .A2(fanout_net_6 ), .ZN(_06386_ ) );
INV_X1 _14282_ ( .A(_06386_ ), .ZN(_06387_ ) );
INV_X1 _14283_ ( .A(fanout_net_6 ), .ZN(_06388_ ) );
OAI21_X1 _14284_ ( .A(_06367_ ), .B1(_06388_ ), .B2(\EX_LS_result_csreg_mem [13] ), .ZN(_06389_ ) );
NOR2_X1 _14285_ ( .A1(fanout_net_6 ), .A2(\EX_LS_result_csreg_mem [21] ), .ZN(_06390_ ) );
OAI22_X1 _14286_ ( .A1(_06387_ ), .A2(_06370_ ), .B1(_06389_ ), .B2(_06390_ ), .ZN(\io_master_wdata [21] ) );
OAI21_X1 _14287_ ( .A(_06367_ ), .B1(_06388_ ), .B2(\EX_LS_result_csreg_mem [12] ), .ZN(_06391_ ) );
NOR2_X1 _14288_ ( .A1(fanout_net_6 ), .A2(\EX_LS_result_csreg_mem [20] ), .ZN(_06392_ ) );
OAI22_X1 _14289_ ( .A1(_06387_ ), .A2(_06371_ ), .B1(_06391_ ), .B2(_06392_ ), .ZN(\io_master_wdata [20] ) );
OAI21_X1 _14290_ ( .A(_06367_ ), .B1(_06388_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_06393_ ) );
NOR2_X1 _14291_ ( .A1(fanout_net_6 ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_06394_ ) );
OAI22_X1 _14292_ ( .A1(_06387_ ), .A2(_06372_ ), .B1(_06393_ ), .B2(_06394_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _14293_ ( .A(_06367_ ), .B1(_06388_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_06395_ ) );
NOR2_X1 _14294_ ( .A1(fanout_net_6 ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_06396_ ) );
OAI22_X1 _14295_ ( .A1(_06387_ ), .A2(_06373_ ), .B1(_06395_ ), .B2(_06396_ ), .ZN(\io_master_wdata [18] ) );
INV_X1 _14296_ ( .A(\EX_LS_result_csreg_mem [17] ), .ZN(_06397_ ) );
INV_X1 _14297_ ( .A(\EX_LS_result_csreg_mem [9] ), .ZN(_06398_ ) );
MUX2_X1 _14298_ ( .A(_06397_ ), .B(_06398_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06399_ ) );
OAI22_X1 _14299_ ( .A1(_06399_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06387_ ), .B2(_06374_ ), .ZN(\io_master_wdata [17] ) );
OAI21_X1 _14300_ ( .A(_06367_ ), .B1(_06388_ ), .B2(\EX_LS_result_csreg_mem [8] ), .ZN(_06400_ ) );
NOR2_X1 _14301_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [16] ), .ZN(_06401_ ) );
OAI22_X1 _14302_ ( .A1(_06387_ ), .A2(_06375_ ), .B1(_06400_ ), .B2(_06401_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14303_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06402_ ) );
MUX2_X1 _14304_ ( .A(_06402_ ), .B(_06376_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14305_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06403_ ) );
MUX2_X1 _14306_ ( .A(_06403_ ), .B(_06377_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14307_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06404_ ) );
MUX2_X1 _14308_ ( .A(_06404_ ), .B(_06378_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14309_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06405_ ) );
MUX2_X1 _14310_ ( .A(_06405_ ), .B(_06379_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14311_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06406_ ) );
MUX2_X1 _14312_ ( .A(_06406_ ), .B(_06380_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14313_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06407_ ) );
MUX2_X1 _14314_ ( .A(_06407_ ), .B(_06381_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [24] ) );
INV_X1 _14315_ ( .A(\EX_LS_result_csreg_mem [23] ), .ZN(_06408_ ) );
INV_X1 _14316_ ( .A(\EX_LS_result_csreg_mem [15] ), .ZN(_06409_ ) );
MUX2_X1 _14317_ ( .A(_06408_ ), .B(_06409_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06410_ ) );
OAI22_X1 _14318_ ( .A1(_06410_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06387_ ), .B2(_06382_ ), .ZN(\io_master_wdata [23] ) );
OAI21_X1 _14319_ ( .A(_06367_ ), .B1(_06388_ ), .B2(\EX_LS_result_csreg_mem [14] ), .ZN(_06411_ ) );
NOR2_X1 _14320_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [22] ), .ZN(_06412_ ) );
OAI22_X1 _14321_ ( .A1(_06387_ ), .A2(_06383_ ), .B1(_06411_ ), .B2(_06412_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14322_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06413_ ) );
AND2_X1 _14323_ ( .A1(_06413_ ), .A2(_06368_ ), .ZN(\io_master_wstrb [1] ) );
NOR3_X1 _14324_ ( .A1(_02233_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14325_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06414_ ) );
MUX2_X1 _14326_ ( .A(_06414_ ), .B(_06413_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14327_ ( .A1(_06368_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_06415_ ) );
OAI221_X1 _14328_ ( .A(_06415_ ), .B1(_02261_ ), .B2(_02235_ ), .C1(_06387_ ), .C2(_02233_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _14329_ ( .A1(_06351_ ), .A2(_06353_ ), .ZN(io_master_wvalid ) );
AND2_X1 _14330_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06416_ ) );
NOR2_X1 _14331_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06417_ ) );
AND2_X1 _14332_ ( .A1(_06416_ ), .A2(_06417_ ), .ZN(_06418_ ) );
NOR4_X1 _14333_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .A3(\LS_WB_waddr_csreg [5] ), .A4(\LS_WB_waddr_csreg [4] ), .ZN(_06419_ ) );
NAND2_X1 _14334_ ( .A1(_06418_ ), .A2(_06419_ ), .ZN(_06420_ ) );
INV_X1 _14335_ ( .A(\LS_WB_wen_csreg [7] ), .ZN(_06421_ ) );
NOR2_X1 _14336_ ( .A1(_06421_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_06422_ ) );
INV_X1 _14337_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_06423_ ) );
INV_X1 _14338_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_06424_ ) );
INV_X1 _14339_ ( .A(\LS_WB_waddr_csreg [2] ), .ZN(_06425_ ) );
NAND4_X1 _14340_ ( .A1(_06422_ ), .A2(_06423_ ), .A3(_06424_ ), .A4(_06425_ ), .ZN(_06426_ ) );
NOR2_X1 _14341_ ( .A1(_06420_ ), .A2(_06426_ ), .ZN(\mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _14342_ ( .A1(_06422_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(_06424_ ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_06427_ ) );
NOR2_X1 _14343_ ( .A1(_06420_ ), .A2(_06427_ ), .ZN(\mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _14344_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06428_ ) );
NAND2_X1 _14345_ ( .A1(_06428_ ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06429_ ) );
NOR2_X1 _14346_ ( .A1(_06429_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06430_ ) );
AND4_X1 _14347_ ( .A1(\LS_WB_waddr_csreg [0] ), .A2(_06430_ ), .A3(_06424_ ), .A4(_06422_ ), .ZN(_06431_ ) );
AND3_X1 _14348_ ( .A1(_06431_ ), .A2(_06425_ ), .A3(_06418_ ), .ZN(\mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14349_ ( .A(_06430_ ), .ZN(_06432_ ) );
NOR4_X1 _14350_ ( .A1(_06432_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(_06424_ ), .A4(\LS_WB_waddr_csreg [3] ), .ZN(_06433_ ) );
NAND3_X1 _14351_ ( .A1(_06433_ ), .A2(_06425_ ), .A3(_06418_ ), .ZN(_06434_ ) );
AOI21_X1 _14352_ ( .A(_06421_ ), .B1(_06434_ ), .B2(_02307_ ), .ZN(\mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _14353_ ( .A(_02316_ ), .B1(_02320_ ), .B2(_02322_ ), .ZN(_06435_ ) );
NAND2_X1 _14354_ ( .A1(_02266_ ), .A2(_06435_ ), .ZN(_06436_ ) );
BUF_X4 _14355_ ( .A(_06436_ ), .Z(_06437_ ) );
MUX2_X1 _14356_ ( .A(\ID_EX_pc [21] ), .B(\EX_LS_pc [21] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14357_ ( .A(\ID_EX_pc [20] ), .B(\EX_LS_pc [20] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14358_ ( .A(\ID_EX_pc [19] ), .B(\EX_LS_pc [19] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14359_ ( .A(\ID_EX_pc [18] ), .B(\EX_LS_pc [18] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14360_ ( .A(\ID_EX_pc [17] ), .B(\EX_LS_pc [17] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14361_ ( .A(\ID_EX_pc [16] ), .B(\EX_LS_pc [16] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14362_ ( .A(\ID_EX_pc [15] ), .B(\EX_LS_pc [15] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14363_ ( .A(\ID_EX_pc [14] ), .B(\EX_LS_pc [14] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14364_ ( .A(\ID_EX_pc [13] ), .B(\EX_LS_pc [13] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14365_ ( .A(\ID_EX_pc [12] ), .B(\EX_LS_pc [12] ), .S(_06437_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14366_ ( .A(_06436_ ), .Z(_06438_ ) );
MUX2_X1 _14367_ ( .A(\ID_EX_pc [30] ), .B(\EX_LS_pc [30] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14368_ ( .A(\ID_EX_pc [11] ), .B(\EX_LS_pc [11] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14369_ ( .A(\ID_EX_pc [10] ), .B(\EX_LS_pc [10] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14370_ ( .A(\ID_EX_pc [9] ), .B(\EX_LS_pc [9] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14371_ ( .A(\ID_EX_pc [8] ), .B(\EX_LS_pc [8] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14372_ ( .A(\ID_EX_pc [7] ), .B(\EX_LS_pc [7] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14373_ ( .A(\ID_EX_pc [6] ), .B(\EX_LS_pc [6] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14374_ ( .A(\ID_EX_pc [5] ), .B(\EX_LS_pc [5] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14375_ ( .A(\ID_EX_pc [4] ), .B(\EX_LS_pc [4] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14376_ ( .A(\ID_EX_pc [3] ), .B(\EX_LS_pc [3] ), .S(_06438_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14377_ ( .A(_06436_ ), .Z(_06439_ ) );
MUX2_X1 _14378_ ( .A(\ID_EX_pc [2] ), .B(\EX_LS_pc [2] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14379_ ( .A(\ID_EX_pc [29] ), .B(\EX_LS_pc [29] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14380_ ( .A(\ID_EX_pc [1] ), .B(\EX_LS_pc [1] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14381_ ( .A(\ID_EX_pc [0] ), .B(\EX_LS_pc [0] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14382_ ( .A(\ID_EX_pc [28] ), .B(\EX_LS_pc [28] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14383_ ( .A(\ID_EX_pc [27] ), .B(\EX_LS_pc [27] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14384_ ( .A(\ID_EX_pc [26] ), .B(\EX_LS_pc [26] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14385_ ( .A(\ID_EX_pc [25] ), .B(\EX_LS_pc [25] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14386_ ( .A(\ID_EX_pc [24] ), .B(\EX_LS_pc [24] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14387_ ( .A(\ID_EX_pc [23] ), .B(\EX_LS_pc [23] ), .S(_06439_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14388_ ( .A(\ID_EX_pc [22] ), .B(\EX_LS_pc [22] ), .S(_06436_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14389_ ( .A(\ID_EX_pc [31] ), .B(\EX_LS_pc [31] ), .S(_06436_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
AOI21_X1 _14390_ ( .A(_02314_ ), .B1(_02253_ ), .B2(_02265_ ), .ZN(_06440_ ) );
AOI21_X1 _14391_ ( .A(_02314_ ), .B1(_02323_ ), .B2(_02316_ ), .ZN(_06441_ ) );
OR2_X1 _14392_ ( .A1(_06440_ ), .A2(_06441_ ), .ZN(\myec.state_$_NOR__A_Y_$_ANDNOT__A_Y ) );
NAND4_X1 _14393_ ( .A1(_02266_ ), .A2(_02316_ ), .A3(_02323_ ), .A4(_02312_ ), .ZN(_06442_ ) );
XNOR2_X1 _14394_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06443_ ) );
XNOR2_X1 _14395_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06444_ ) );
XNOR2_X1 _14396_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06445_ ) );
XNOR2_X1 _14397_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06446_ ) );
AND4_X1 _14398_ ( .A1(_06443_ ), .A2(_06444_ ), .A3(_06445_ ), .A4(_06446_ ), .ZN(_06447_ ) );
XNOR2_X1 _14399_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06448_ ) );
XNOR2_X1 _14400_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06449_ ) );
XNOR2_X1 _14401_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06450_ ) );
XNOR2_X1 _14402_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06451_ ) );
AND4_X1 _14403_ ( .A1(_06448_ ), .A2(_06449_ ), .A3(_06450_ ), .A4(_06451_ ), .ZN(_06452_ ) );
XNOR2_X1 _14404_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_06453_ ) );
XNOR2_X1 _14405_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_06454_ ) );
XNOR2_X1 _14406_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_06455_ ) );
XNOR2_X1 _14407_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_06456_ ) );
AND4_X1 _14408_ ( .A1(_06453_ ), .A2(_06454_ ), .A3(_06455_ ), .A4(_06456_ ), .ZN(_06457_ ) );
XNOR2_X1 _14409_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06458_ ) );
XNOR2_X1 _14410_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06459_ ) );
XNOR2_X1 _14411_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06460_ ) );
XNOR2_X1 _14412_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06461_ ) );
AND4_X1 _14413_ ( .A1(_06458_ ), .A2(_06459_ ), .A3(_06460_ ), .A4(_06461_ ), .ZN(_06462_ ) );
AND4_X1 _14414_ ( .A1(_06447_ ), .A2(_06452_ ), .A3(_06457_ ), .A4(_06462_ ), .ZN(_06463_ ) );
XNOR2_X1 _14415_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06464_ ) );
XNOR2_X1 _14416_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06465_ ) );
XNOR2_X1 _14417_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06466_ ) );
XNOR2_X1 _14418_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06467_ ) );
AND4_X1 _14419_ ( .A1(_06464_ ), .A2(_06465_ ), .A3(_06466_ ), .A4(_06467_ ), .ZN(_06468_ ) );
XNOR2_X1 _14420_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06469_ ) );
XNOR2_X1 _14421_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06470_ ) );
XNOR2_X1 _14422_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06471_ ) );
XNOR2_X1 _14423_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06472_ ) );
AND4_X1 _14424_ ( .A1(_06469_ ), .A2(_06470_ ), .A3(_06471_ ), .A4(_06472_ ), .ZN(_06473_ ) );
XNOR2_X1 _14425_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06474_ ) );
XNOR2_X1 _14426_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06475_ ) );
XNOR2_X1 _14427_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06476_ ) );
XNOR2_X1 _14428_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06477_ ) );
AND4_X1 _14429_ ( .A1(_06474_ ), .A2(_06475_ ), .A3(_06476_ ), .A4(_06477_ ), .ZN(_06478_ ) );
XNOR2_X1 _14430_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06479_ ) );
XNOR2_X1 _14431_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06480_ ) );
XNOR2_X1 _14432_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06481_ ) );
XNOR2_X1 _14433_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06482_ ) );
AND4_X1 _14434_ ( .A1(_06479_ ), .A2(_06480_ ), .A3(_06481_ ), .A4(_06482_ ), .ZN(_06483_ ) );
AND4_X1 _14435_ ( .A1(_06468_ ), .A2(_06473_ ), .A3(_06478_ ), .A4(_06483_ ), .ZN(_06484_ ) );
NAND3_X1 _14436_ ( .A1(_06463_ ), .A2(_06484_ ), .A3(excp_written ), .ZN(_06485_ ) );
OAI21_X1 _14437_ ( .A(_06485_ ), .B1(\myec.state [1] ), .B2(\myec.state [0] ), .ZN(_06486_ ) );
AND2_X1 _14438_ ( .A1(_06442_ ), .A2(_06486_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14439_ ( .A1(_06068_ ), .A2(_03257_ ), .ZN(_06487_ ) );
AND2_X1 _14440_ ( .A1(_03246_ ), .A2(_04150_ ), .ZN(_06488_ ) );
BUF_X4 _14441_ ( .A(_06488_ ), .Z(_06489_ ) );
INV_X1 _14442_ ( .A(_06489_ ), .ZN(_06490_ ) );
BUF_X4 _14443_ ( .A(_06490_ ), .Z(_06491_ ) );
BUF_X4 _14444_ ( .A(_06491_ ), .Z(_06492_ ) );
OAI21_X1 _14445_ ( .A(_06487_ ), .B1(_05503_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _14446_ ( .A(_05116_ ), .B(\ID_EX_imm [0] ), .ZN(_06493_ ) );
BUF_X4 _14447_ ( .A(_06489_ ), .Z(_06494_ ) );
AOI22_X1 _14448_ ( .A1(_06493_ ), .A2(_03257_ ), .B1(_05495_ ), .B2(_06494_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
NAND2_X1 _14449_ ( .A1(_05897_ ), .A2(_03257_ ), .ZN(_06495_ ) );
OAI21_X1 _14450_ ( .A(_06495_ ), .B1(_05484_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
AOI22_X1 _14451_ ( .A1(_05918_ ), .A2(_03257_ ), .B1(_05532_ ), .B2(_06494_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
NOR2_X1 _14452_ ( .A1(_05935_ ), .A2(_03247_ ), .ZN(_06496_ ) );
BUF_X4 _14453_ ( .A(_06489_ ), .Z(_06497_ ) );
BUF_X4 _14454_ ( .A(_06497_ ), .Z(_06498_ ) );
AOI21_X1 _14455_ ( .A(_06496_ ), .B1(_05533_ ), .B2(_06498_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _14456_ ( .A1(_05956_ ), .A2(_03257_ ), .ZN(_06499_ ) );
OAI21_X1 _14457_ ( .A(_06499_ ), .B1(_05492_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
AND2_X1 _14458_ ( .A1(_03604_ ), .A2(\ID_EX_typ [7] ), .ZN(_06500_ ) );
OR2_X1 _14459_ ( .A1(_05976_ ), .A2(_06500_ ), .ZN(_06501_ ) );
BUF_X2 _14460_ ( .A(_06490_ ), .Z(_06502_ ) );
MUX2_X1 _14461_ ( .A(\ID_EX_csr [6] ), .B(_06501_ ), .S(_06502_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14462_ ( .A1(_05997_ ), .A2(_03256_ ), .ZN(_06503_ ) );
OAI21_X1 _14463_ ( .A(_06503_ ), .B1(_05485_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _14464_ ( .A1(_06016_ ), .A2(_03256_ ), .ZN(_06504_ ) );
OAI21_X1 _14465_ ( .A(_06504_ ), .B1(_05486_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _14466_ ( .A1(_06036_ ), .A2(_03256_ ), .ZN(_06505_ ) );
OAI21_X1 _14467_ ( .A(_06505_ ), .B1(_05509_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _14468_ ( .A1(_06051_ ), .A2(_03256_ ), .ZN(_06506_ ) );
OAI21_X1 _14469_ ( .A(_06506_ ), .B1(_05519_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
NAND2_X1 _14470_ ( .A1(_05836_ ), .A2(_03256_ ), .ZN(_06507_ ) );
OAI21_X1 _14471_ ( .A(_06507_ ), .B1(_05487_ ), .B2(_06492_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X4 _14472_ ( .A(_06489_ ), .Z(_06508_ ) );
AND3_X1 _14473_ ( .A1(_06210_ ), .A2(\ID_EX_typ [2] ), .A3(_06211_ ), .ZN(_06509_ ) );
NAND3_X1 _14474_ ( .A1(_02565_ ), .A2(_05661_ ), .A3(_02585_ ), .ZN(_06510_ ) );
NAND2_X1 _14475_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [21] ), .ZN(_06511_ ) );
AOI21_X1 _14476_ ( .A(_06509_ ), .B1(_06510_ ), .B2(_06511_ ), .ZN(_06512_ ) );
NOR2_X1 _14477_ ( .A1(_05125_ ), .A2(\ID_EX_typ [2] ), .ZN(_06513_ ) );
INV_X1 _14478_ ( .A(_06513_ ), .ZN(_06514_ ) );
BUF_X4 _14479_ ( .A(_06514_ ), .Z(_06515_ ) );
AOI21_X1 _14480_ ( .A(_06515_ ), .B1(_06210_ ), .B2(_06211_ ), .ZN(_06516_ ) );
OAI21_X1 _14481_ ( .A(_06508_ ), .B1(_06512_ ), .B2(_06516_ ), .ZN(_06517_ ) );
BUF_X4 _14482_ ( .A(_06497_ ), .Z(_06518_ ) );
INV_X1 _14483_ ( .A(_06500_ ), .ZN(_06519_ ) );
BUF_X4 _14484_ ( .A(_06519_ ), .Z(_06520_ ) );
MUX2_X1 _14485_ ( .A(_06197_ ), .B(_04526_ ), .S(_06520_ ), .Z(_06521_ ) );
OAI21_X1 _14486_ ( .A(_06517_ ), .B1(_06518_ ), .B2(_06521_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
OAI211_X1 _14487_ ( .A(_03247_ ), .B(_04150_ ), .C1(_05732_ ), .C2(\ID_EX_imm [20] ), .ZN(_06522_ ) );
AOI21_X1 _14488_ ( .A(_06522_ ), .B1(_05331_ ), .B2(_06215_ ), .ZN(_06523_ ) );
OAI21_X1 _14489_ ( .A(_06523_ ), .B1(_06266_ ), .B2(_05614_ ), .ZN(_06524_ ) );
BUF_X4 _14490_ ( .A(_06513_ ), .Z(_06525_ ) );
BUF_X4 _14491_ ( .A(_06489_ ), .Z(_06526_ ) );
NAND3_X1 _14492_ ( .A1(_05614_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(_06527_ ) );
BUF_X4 _14493_ ( .A(_06519_ ), .Z(_06528_ ) );
MUX2_X1 _14494_ ( .A(_06195_ ), .B(_04503_ ), .S(_06528_ ), .Z(_06529_ ) );
OAI211_X1 _14495_ ( .A(_06524_ ), .B(_06527_ ), .C1(_06498_ ), .C2(_06529_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
AOI211_X1 _14496_ ( .A(_06265_ ), .B(_05656_ ), .C1(_05650_ ), .C2(_05652_ ), .ZN(_06530_ ) );
AOI21_X1 _14497_ ( .A(fanout_net_7 ), .B1(_02638_ ), .B2(_02658_ ), .ZN(_06531_ ) );
NOR2_X1 _14498_ ( .A1(_05685_ ), .A2(\ID_EX_imm [19] ), .ZN(_06532_ ) );
NOR3_X1 _14499_ ( .A1(_06530_ ), .A2(_06531_ ), .A3(_06532_ ), .ZN(_06533_ ) );
AOI21_X1 _14500_ ( .A(_06515_ ), .B1(_05653_ ), .B2(_05657_ ), .ZN(_06534_ ) );
OAI21_X1 _14501_ ( .A(_06508_ ), .B1(_06533_ ), .B2(_06534_ ), .ZN(_06535_ ) );
MUX2_X1 _14502_ ( .A(_05635_ ), .B(_04406_ ), .S(_06520_ ), .Z(_06536_ ) );
OAI21_X1 _14503_ ( .A(_06535_ ), .B1(_06518_ ), .B2(_06536_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
OAI211_X1 _14504_ ( .A(_03247_ ), .B(_04150_ ), .C1(_05732_ ), .C2(\ID_EX_imm [18] ), .ZN(_06537_ ) );
INV_X1 _14505_ ( .A(_02635_ ), .ZN(_06538_ ) );
AOI21_X1 _14506_ ( .A(_06537_ ), .B1(_06538_ ), .B2(_06215_ ), .ZN(_06539_ ) );
OAI21_X1 _14507_ ( .A(_06539_ ), .B1(_06266_ ), .B2(_05683_ ), .ZN(_06540_ ) );
NAND3_X1 _14508_ ( .A1(_05683_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(_06541_ ) );
MUX2_X1 _14509_ ( .A(_05664_ ), .B(_04429_ ), .S(_06528_ ), .Z(_06542_ ) );
OAI211_X1 _14510_ ( .A(_06540_ ), .B(_06541_ ), .C1(_06498_ ), .C2(_06542_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
AND3_X1 _14511_ ( .A1(_05654_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_05655_ ), .ZN(_06543_ ) );
AOI211_X1 _14512_ ( .A(_06265_ ), .B(_06543_ ), .C1(_05704_ ), .C2(_05652_ ), .ZN(_06544_ ) );
AOI21_X1 _14513_ ( .A(fanout_net_7 ), .B1(_02663_ ), .B2(_02683_ ), .ZN(_06545_ ) );
NOR2_X1 _14514_ ( .A1(_05685_ ), .A2(\ID_EX_imm [17] ), .ZN(_06546_ ) );
NOR3_X1 _14515_ ( .A1(_06544_ ), .A2(_06545_ ), .A3(_06546_ ), .ZN(_06547_ ) );
AOI21_X1 _14516_ ( .A(_06515_ ), .B1(_05705_ ), .B2(_05706_ ), .ZN(_06548_ ) );
OAI21_X1 _14517_ ( .A(_06508_ ), .B1(_06547_ ), .B2(_06548_ ), .ZN(_06549_ ) );
MUX2_X1 _14518_ ( .A(_06241_ ), .B(_04375_ ), .S(_06520_ ), .Z(_06550_ ) );
OAI21_X1 _14519_ ( .A(_06549_ ), .B1(_06518_ ), .B2(_06550_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
AOI211_X1 _14520_ ( .A(_06265_ ), .B(_05723_ ), .C1(_05721_ ), .C2(_05652_ ), .ZN(_06551_ ) );
NAND3_X1 _14521_ ( .A1(_02687_ ), .A2(_05661_ ), .A3(_02707_ ), .ZN(_06552_ ) );
NAND2_X1 _14522_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [16] ), .ZN(_06553_ ) );
AOI21_X1 _14523_ ( .A(_06551_ ), .B1(_06552_ ), .B2(_06553_ ), .ZN(_06554_ ) );
AOI21_X1 _14524_ ( .A(_06515_ ), .B1(_05722_ ), .B2(_05724_ ), .ZN(_06555_ ) );
OAI21_X1 _14525_ ( .A(_06508_ ), .B1(_06554_ ), .B2(_06555_ ), .ZN(_06556_ ) );
MUX2_X1 _14526_ ( .A(_05693_ ), .B(_04352_ ), .S(_06520_ ), .Z(_06557_ ) );
OAI21_X1 _14527_ ( .A(_06556_ ), .B1(_06518_ ), .B2(_06557_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
NAND3_X1 _14528_ ( .A1(_02975_ ), .A2(_05685_ ), .A3(_02995_ ), .ZN(_06558_ ) );
NAND2_X1 _14529_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [15] ), .ZN(_06559_ ) );
NAND2_X1 _14530_ ( .A1(_06558_ ), .A2(_06559_ ), .ZN(_06560_ ) );
AOI21_X1 _14531_ ( .A(_06514_ ), .B1(_05750_ ), .B2(_05751_ ), .ZN(_06561_ ) );
OAI221_X1 _14532_ ( .A(_06508_ ), .B1(_06560_ ), .B2(_06561_ ), .C1(_05753_ ), .C2(_06266_ ), .ZN(_06562_ ) );
BUF_X4 _14533_ ( .A(_06491_ ), .Z(_06563_ ) );
NAND4_X1 _14534_ ( .A1(_06242_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06564_ ) );
OAI211_X1 _14535_ ( .A(_06563_ ), .B(_06564_ ), .C1(_04778_ ), .C2(_06500_ ), .ZN(_06565_ ) );
NAND2_X1 _14536_ ( .A1(_06562_ ), .A2(_06565_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
AOI211_X1 _14537_ ( .A(_06265_ ), .B(_05765_ ), .C1(_05763_ ), .C2(_05652_ ), .ZN(_06566_ ) );
AOI21_X1 _14538_ ( .A(fanout_net_7 ), .B1(_02998_ ), .B2(_03018_ ), .ZN(_06567_ ) );
NOR2_X1 _14539_ ( .A1(_05685_ ), .A2(\ID_EX_imm [14] ), .ZN(_06568_ ) );
NOR3_X1 _14540_ ( .A1(_06566_ ), .A2(_06567_ ), .A3(_06568_ ), .ZN(_06569_ ) );
AOI21_X1 _14541_ ( .A(_06515_ ), .B1(_05764_ ), .B2(_05766_ ), .ZN(_06570_ ) );
OAI21_X1 _14542_ ( .A(_06508_ ), .B1(_06569_ ), .B2(_06570_ ), .ZN(_06571_ ) );
MUX2_X1 _14543_ ( .A(_05769_ ), .B(_04752_ ), .S(_06520_ ), .Z(_06572_ ) );
OAI21_X1 _14544_ ( .A(_06571_ ), .B1(_06518_ ), .B2(_06572_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OAI211_X1 _14545_ ( .A(_03247_ ), .B(_04150_ ), .C1(_05732_ ), .C2(\ID_EX_imm [13] ), .ZN(_06573_ ) );
INV_X1 _14546_ ( .A(_04781_ ), .ZN(_06574_ ) );
AOI21_X1 _14547_ ( .A(_06573_ ), .B1(_06574_ ), .B2(_06140_ ), .ZN(_06575_ ) );
OAI21_X1 _14548_ ( .A(_06575_ ), .B1(_06266_ ), .B2(_05786_ ), .ZN(_06576_ ) );
NAND3_X1 _14549_ ( .A1(_05786_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(_06577_ ) );
MUX2_X1 _14550_ ( .A(_05559_ ), .B(_04804_ ), .S(_06528_ ), .Z(_06578_ ) );
OAI211_X1 _14551_ ( .A(_06576_ ), .B(_06577_ ), .C1(_06498_ ), .C2(_06578_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AOI211_X1 _14552_ ( .A(_06265_ ), .B(_05808_ ), .C1(_05806_ ), .C2(_05652_ ), .ZN(_06579_ ) );
NAND3_X1 _14553_ ( .A1(_02926_ ), .A2(_05661_ ), .A3(_02946_ ), .ZN(_06580_ ) );
NAND2_X1 _14554_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [12] ), .ZN(_06581_ ) );
AOI21_X1 _14555_ ( .A(_06579_ ), .B1(_06580_ ), .B2(_06581_ ), .ZN(_06582_ ) );
AOI21_X1 _14556_ ( .A(_06515_ ), .B1(_05807_ ), .B2(_05809_ ), .ZN(_06583_ ) );
OAI21_X1 _14557_ ( .A(_06508_ ), .B1(_06582_ ), .B2(_06583_ ), .ZN(_06584_ ) );
MUX2_X1 _14558_ ( .A(_05560_ ), .B(_04827_ ), .S(_06520_ ), .Z(_06585_ ) );
OAI21_X1 _14559_ ( .A(_06584_ ), .B1(_06518_ ), .B2(_06585_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
OAI211_X1 _14560_ ( .A(_02400_ ), .B(_04146_ ), .C1(_02373_ ), .C2(_02398_ ), .ZN(_06586_ ) );
NAND2_X1 _14561_ ( .A1(_02402_ ), .A2(fanout_net_7 ), .ZN(_06587_ ) );
NAND3_X1 _14562_ ( .A1(_05547_ ), .A2(\ID_EX_typ [2] ), .A3(_05548_ ), .ZN(_06588_ ) );
NAND3_X1 _14563_ ( .A1(_06586_ ), .A2(_06587_ ), .A3(_06588_ ), .ZN(_06589_ ) );
OR2_X1 _14564_ ( .A1(_05549_ ), .A2(_06514_ ), .ZN(_06590_ ) );
AND3_X1 _14565_ ( .A1(_06589_ ), .A2(_06489_ ), .A3(_06590_ ), .ZN(_06591_ ) );
BUF_X4 _14566_ ( .A(_06519_ ), .Z(_06592_ ) );
MUX2_X1 _14567_ ( .A(_06235_ ), .B(_04606_ ), .S(_06592_ ), .Z(_06593_ ) );
AOI21_X1 _14568_ ( .A(_06591_ ), .B1(_06492_ ), .B2(_06593_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
OAI211_X1 _14569_ ( .A(_03246_ ), .B(_04150_ ), .C1(_05732_ ), .C2(\ID_EX_imm [11] ), .ZN(_06594_ ) );
AOI21_X1 _14570_ ( .A(_06594_ ), .B1(_05187_ ), .B2(_06140_ ), .ZN(_06595_ ) );
OAI21_X1 _14571_ ( .A(_06595_ ), .B1(_06266_ ), .B2(_05829_ ), .ZN(_06596_ ) );
NAND3_X1 _14572_ ( .A1(_05829_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(_06597_ ) );
MUX2_X1 _14573_ ( .A(_06243_ ), .B(_04852_ ), .S(_06528_ ), .Z(_06598_ ) );
OAI211_X1 _14574_ ( .A(_06596_ ), .B(_06597_ ), .C1(_06498_ ), .C2(_06598_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI211_X1 _14575_ ( .A(_05127_ ), .B(_05886_ ), .C1(_05884_ ), .C2(_05652_ ), .ZN(_06599_ ) );
NAND3_X1 _14576_ ( .A1(_03073_ ), .A2(_05685_ ), .A3(_03093_ ), .ZN(_06600_ ) );
NAND2_X1 _14577_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [10] ), .ZN(_06601_ ) );
AOI21_X1 _14578_ ( .A(_06599_ ), .B1(_06600_ ), .B2(_06601_ ), .ZN(_06602_ ) );
AOI21_X1 _14579_ ( .A(_06515_ ), .B1(_05885_ ), .B2(_05887_ ), .ZN(_06603_ ) );
OAI21_X1 _14580_ ( .A(_06508_ ), .B1(_06602_ ), .B2(_06603_ ), .ZN(_06604_ ) );
MUX2_X1 _14581_ ( .A(_05890_ ), .B(_04876_ ), .S(_06520_ ), .Z(_06605_ ) );
OAI21_X1 _14582_ ( .A(_06604_ ), .B1(_06518_ ), .B2(_06605_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
OAI211_X1 _14583_ ( .A(_03246_ ), .B(_04150_ ), .C1(_05732_ ), .C2(\ID_EX_imm [9] ), .ZN(_06606_ ) );
AOI21_X1 _14584_ ( .A(_06606_ ), .B1(_05201_ ), .B2(_06140_ ), .ZN(_06607_ ) );
OAI21_X1 _14585_ ( .A(_06607_ ), .B1(_06266_ ), .B2(_05914_ ), .ZN(_06608_ ) );
NAND3_X1 _14586_ ( .A1(_05914_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(_06609_ ) );
MUX2_X1 _14587_ ( .A(_05899_ ), .B(_04924_ ), .S(_06528_ ), .Z(_06610_ ) );
OAI211_X1 _14588_ ( .A(_06608_ ), .B(_06609_ ), .C1(_06498_ ), .C2(_06610_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
OAI211_X1 _14589_ ( .A(_03246_ ), .B(_04150_ ), .C1(_05732_ ), .C2(\ID_EX_imm [8] ), .ZN(_06611_ ) );
AOI21_X1 _14590_ ( .A(_06611_ ), .B1(_05278_ ), .B2(_06140_ ), .ZN(_06612_ ) );
OAI21_X1 _14591_ ( .A(_06612_ ), .B1(_06266_ ), .B2(_05929_ ), .ZN(_06613_ ) );
NAND3_X1 _14592_ ( .A1(_05929_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(_06614_ ) );
MUX2_X1 _14593_ ( .A(_06244_ ), .B(_04900_ ), .S(_06528_ ), .Z(_06615_ ) );
OAI211_X1 _14594_ ( .A(_06613_ ), .B(_06614_ ), .C1(_06498_ ), .C2(_06615_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
OAI211_X1 _14595_ ( .A(_03246_ ), .B(_04150_ ), .C1(_05732_ ), .C2(\ID_EX_imm [7] ), .ZN(_06616_ ) );
OR3_X1 _14596_ ( .A1(_05863_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_05864_ ), .ZN(_06617_ ) );
NAND3_X1 _14597_ ( .A1(_05861_ ), .A2(\mtvec [7] ), .A3(_05644_ ), .ZN(_06618_ ) );
NAND3_X1 _14598_ ( .A1(_05861_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_05702_ ), .ZN(_06619_ ) );
AND2_X1 _14599_ ( .A1(_06618_ ), .A2(_06619_ ), .ZN(_06620_ ) );
NAND3_X1 _14600_ ( .A1(_06620_ ), .A2(_05938_ ), .A3(_05939_ ), .ZN(_06621_ ) );
OAI21_X1 _14601_ ( .A(_06617_ ), .B1(_06621_ ), .B2(_06233_ ), .ZN(_06622_ ) );
AOI21_X1 _14602_ ( .A(_06616_ ), .B1(_06622_ ), .B2(\ID_EX_typ [2] ), .ZN(_06623_ ) );
OAI21_X1 _14603_ ( .A(_06623_ ), .B1(_02812_ ), .B2(fanout_net_7 ), .ZN(_06624_ ) );
NAND3_X1 _14604_ ( .A1(_05943_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(_06625_ ) );
MUX2_X1 _14605_ ( .A(_05944_ ), .B(_05045_ ), .S(_06520_ ), .Z(_06626_ ) );
BUF_X4 _14606_ ( .A(_06489_ ), .Z(_06627_ ) );
BUF_X4 _14607_ ( .A(_06627_ ), .Z(_06628_ ) );
OAI211_X1 _14608_ ( .A(_06624_ ), .B(_06625_ ), .C1(_06626_ ), .C2(_06628_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
AOI211_X1 _14609_ ( .A(_06265_ ), .B(_05970_ ), .C1(_05652_ ), .C2(_05968_ ), .ZN(_06629_ ) );
AOI21_X1 _14610_ ( .A(fanout_net_7 ), .B1(_02785_ ), .B2(_02786_ ), .ZN(_06630_ ) );
NOR2_X1 _14611_ ( .A1(_05685_ ), .A2(\ID_EX_imm [6] ), .ZN(_06631_ ) );
NOR3_X1 _14612_ ( .A1(_06629_ ), .A2(_06630_ ), .A3(_06631_ ), .ZN(_06632_ ) );
AOI21_X1 _14613_ ( .A(_06515_ ), .B1(_05969_ ), .B2(_05971_ ), .ZN(_06633_ ) );
OAI21_X1 _14614_ ( .A(_06526_ ), .B1(_06632_ ), .B2(_06633_ ), .ZN(_06634_ ) );
MUX2_X1 _14615_ ( .A(_05958_ ), .B(_05069_ ), .S(_06520_ ), .Z(_06635_ ) );
OAI21_X1 _14616_ ( .A(_06634_ ), .B1(_06518_ ), .B2(_06635_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
AND3_X1 _14617_ ( .A1(_05985_ ), .A2(\ID_EX_typ [2] ), .A3(_05986_ ), .ZN(_06636_ ) );
NOR2_X1 _14618_ ( .A1(_05685_ ), .A2(\ID_EX_imm [5] ), .ZN(_06637_ ) );
AOI21_X1 _14619_ ( .A(fanout_net_7 ), .B1(_02739_ ), .B2(_02762_ ), .ZN(_06638_ ) );
NOR3_X1 _14620_ ( .A1(_06636_ ), .A2(_06637_ ), .A3(_06638_ ), .ZN(_06639_ ) );
AOI21_X1 _14621_ ( .A(_06515_ ), .B1(_05985_ ), .B2(_05986_ ), .ZN(_06640_ ) );
OAI21_X1 _14622_ ( .A(_06526_ ), .B1(_06639_ ), .B2(_06640_ ), .ZN(_06641_ ) );
AND4_X1 _14623_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06642_ ) );
AOI21_X1 _14624_ ( .A(_06642_ ), .B1(_05091_ ), .B2(_06592_ ), .ZN(_06643_ ) );
OAI21_X1 _14625_ ( .A(_06641_ ), .B1(_06518_ ), .B2(_06643_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
AND3_X1 _14626_ ( .A1(_06011_ ), .A2(\ID_EX_typ [2] ), .A3(_06012_ ), .ZN(_06644_ ) );
NOR2_X1 _14627_ ( .A1(_05685_ ), .A2(\ID_EX_imm [4] ), .ZN(_06645_ ) );
AOI21_X1 _14628_ ( .A(fanout_net_7 ), .B1(_02713_ ), .B2(_02734_ ), .ZN(_06646_ ) );
NOR3_X1 _14629_ ( .A1(_06644_ ), .A2(_06645_ ), .A3(_06646_ ), .ZN(_06647_ ) );
AOI21_X1 _14630_ ( .A(_06514_ ), .B1(_06011_ ), .B2(_06012_ ), .ZN(_06648_ ) );
OAI21_X1 _14631_ ( .A(_06526_ ), .B1(_06647_ ), .B2(_06648_ ), .ZN(_06649_ ) );
MUX2_X1 _14632_ ( .A(_06245_ ), .B(_04998_ ), .S(_06520_ ), .Z(_06650_ ) );
OAI21_X1 _14633_ ( .A(_06649_ ), .B1(_06518_ ), .B2(_06650_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _14634_ ( .A1(_02910_ ), .A2(_06140_ ), .ZN(_06651_ ) );
NAND2_X1 _14635_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [3] ), .ZN(_06652_ ) );
NAND2_X1 _14636_ ( .A1(_06651_ ), .A2(_06652_ ), .ZN(_06653_ ) );
AOI21_X1 _14637_ ( .A(_06515_ ), .B1(_06024_ ), .B2(_06025_ ), .ZN(_06654_ ) );
OAI221_X1 _14638_ ( .A(_06508_ ), .B1(_06266_ ), .B2(_06027_ ), .C1(_06653_ ), .C2(_06654_ ), .ZN(_06655_ ) );
NAND4_X1 _14639_ ( .A1(_04191_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06656_ ) );
OAI211_X1 _14640_ ( .A(_06563_ ), .B(_06656_ ), .C1(_04951_ ), .C2(_06500_ ), .ZN(_06657_ ) );
NAND2_X1 _14641_ ( .A1(_06655_ ), .A2(_06657_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
OR3_X1 _14642_ ( .A1(_05844_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_05846_ ), .ZN(_06658_ ) );
NAND2_X1 _14643_ ( .A1(_05850_ ), .A2(_05648_ ), .ZN(_06659_ ) );
NAND3_X1 _14644_ ( .A1(_05857_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_06063_ ), .ZN(_06660_ ) );
NAND4_X1 _14645_ ( .A1(_06043_ ), .A2(_06039_ ), .A3(_06659_ ), .A4(_06660_ ), .ZN(_06661_ ) );
NAND3_X1 _14646_ ( .A1(_05857_ ), .A2(\mtvec [2] ), .A3(_05644_ ), .ZN(_06662_ ) );
OAI21_X1 _14647_ ( .A(_06662_ ), .B1(_05863_ ), .B2(_05864_ ), .ZN(_06663_ ) );
OAI21_X1 _14648_ ( .A(_06658_ ), .B1(_06661_ ), .B2(_06663_ ), .ZN(_06664_ ) );
AOI22_X1 _14649_ ( .A1(_05227_ ), .A2(_06140_ ), .B1(\ID_EX_typ [2] ), .B2(_06664_ ), .ZN(_06665_ ) );
OAI211_X1 _14650_ ( .A(_06665_ ), .B(_06497_ ), .C1(_06215_ ), .C2(\ID_EX_imm [2] ), .ZN(_06666_ ) );
OR3_X1 _14651_ ( .A1(_06664_ ), .A2(_06514_ ), .A3(_06490_ ), .ZN(_06667_ ) );
MUX2_X1 _14652_ ( .A(_06246_ ), .B(_05020_ ), .S(_06528_ ), .Z(_06668_ ) );
OAI211_X1 _14653_ ( .A(_06666_ ), .B(_06667_ ), .C1(_06498_ ), .C2(_06668_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
AOI21_X1 _14654_ ( .A(fanout_net_7 ), .B1(_02423_ ), .B2(_02424_ ), .ZN(_06669_ ) );
AND2_X1 _14655_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [29] ), .ZN(_06670_ ) );
OAI221_X1 _14656_ ( .A(_06627_ ), .B1(_06265_ ), .B2(_05597_ ), .C1(_06669_ ), .C2(_06670_ ), .ZN(_06671_ ) );
AND3_X1 _14657_ ( .A1(_05911_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_05594_ ), .ZN(_06672_ ) );
NOR2_X1 _14658_ ( .A1(_06672_ ), .A2(_05851_ ), .ZN(_06673_ ) );
INV_X1 _14659_ ( .A(_06233_ ), .ZN(_06674_ ) );
NAND3_X1 _14660_ ( .A1(_05857_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_06063_ ), .ZN(_06675_ ) );
AND2_X1 _14661_ ( .A1(_05584_ ), .A2(_06675_ ), .ZN(_06676_ ) );
NAND3_X1 _14662_ ( .A1(_05857_ ), .A2(\mtvec [29] ), .A3(_05679_ ), .ZN(_06677_ ) );
NAND4_X1 _14663_ ( .A1(_06673_ ), .A2(_06674_ ), .A3(_06676_ ), .A4(_06677_ ), .ZN(_06678_ ) );
OR3_X1 _14664_ ( .A1(_05863_ ), .A2(\EX_LS_result_csreg_mem [29] ), .A3(_05864_ ), .ZN(_06679_ ) );
NAND4_X1 _14665_ ( .A1(_06678_ ), .A2(_06525_ ), .A3(_06679_ ), .A4(_06627_ ), .ZN(_06680_ ) );
AND3_X1 _14666_ ( .A1(_03604_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_typ [7] ), .ZN(_06681_ ) );
AOI21_X1 _14667_ ( .A(_06681_ ), .B1(_04581_ ), .B2(_06592_ ), .ZN(_06682_ ) );
OAI211_X1 _14668_ ( .A(_06671_ ), .B(_06680_ ), .C1(_06498_ ), .C2(_06682_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR3_X1 _14669_ ( .A1(_05863_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_05864_ ), .ZN(_06683_ ) );
NAND3_X1 _14670_ ( .A1(_05861_ ), .A2(\mtvec [1] ), .A3(_05644_ ), .ZN(_06684_ ) );
NAND3_X1 _14671_ ( .A1(_05861_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_05702_ ), .ZN(_06685_ ) );
AND2_X1 _14672_ ( .A1(_06684_ ), .A2(_06685_ ), .ZN(_06686_ ) );
NAND3_X1 _14673_ ( .A1(_06686_ ), .A2(_06058_ ), .A3(_06059_ ), .ZN(_06687_ ) );
OAI21_X1 _14674_ ( .A(_06683_ ), .B1(_06687_ ), .B2(_06233_ ), .ZN(_06688_ ) );
AOI22_X1 _14675_ ( .A1(_06688_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02836_ ), .ZN(_06689_ ) );
OAI211_X1 _14676_ ( .A(_06497_ ), .B(_06689_ ), .C1(_02835_ ), .C2(fanout_net_7 ), .ZN(_06690_ ) );
AND2_X1 _14677_ ( .A1(_06058_ ), .A2(_06059_ ), .ZN(_06691_ ) );
NAND3_X1 _14678_ ( .A1(_06674_ ), .A2(_06691_ ), .A3(_06686_ ), .ZN(_06692_ ) );
NAND4_X1 _14679_ ( .A1(_06692_ ), .A2(_06525_ ), .A3(_06683_ ), .A4(_06627_ ), .ZN(_06693_ ) );
MUX2_X1 _14680_ ( .A(_06055_ ), .B(_05113_ ), .S(_06528_ ), .Z(_06694_ ) );
OAI211_X1 _14681_ ( .A(_06690_ ), .B(_06693_ ), .C1(_06498_ ), .C2(_06694_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
NAND3_X1 _14682_ ( .A1(_02838_ ), .A2(_05685_ ), .A3(_02859_ ), .ZN(_06695_ ) );
NAND2_X1 _14683_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [0] ), .ZN(_06696_ ) );
NAND2_X1 _14684_ ( .A1(_06695_ ), .A2(_06696_ ), .ZN(_06697_ ) );
AOI21_X1 _14685_ ( .A(_06514_ ), .B1(_06095_ ), .B2(_06096_ ), .ZN(_06698_ ) );
OAI221_X1 _14686_ ( .A(_06508_ ), .B1(_06697_ ), .B2(_06698_ ), .C1(_06098_ ), .C2(_06266_ ), .ZN(_06699_ ) );
NAND3_X1 _14687_ ( .A1(_04955_ ), .A2(_04975_ ), .A3(_06592_ ), .ZN(_06700_ ) );
OAI211_X1 _14688_ ( .A(_06700_ ), .B(_06563_ ), .C1(\ID_EX_pc [0] ), .C2(_06592_ ), .ZN(_06701_ ) );
NAND2_X1 _14689_ ( .A1(_06699_ ), .A2(_06701_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
AOI22_X1 _14690_ ( .A1(_05160_ ), .A2(_06140_ ), .B1(\ID_EX_typ [2] ), .B2(_05866_ ), .ZN(_06702_ ) );
OAI211_X1 _14691_ ( .A(_06702_ ), .B(_06497_ ), .C1(_06215_ ), .C2(\ID_EX_imm [28] ), .ZN(_06703_ ) );
OR3_X1 _14692_ ( .A1(_05866_ ), .A2(_06514_ ), .A3(_06490_ ), .ZN(_06704_ ) );
MUX2_X1 _14693_ ( .A(_05839_ ), .B(_05445_ ), .S(_06528_ ), .Z(_06705_ ) );
OAI211_X1 _14694_ ( .A(_06703_ ), .B(_06704_ ), .C1(_06628_ ), .C2(_06705_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
OR3_X1 _14695_ ( .A1(_05844_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_05846_ ), .ZN(_06706_ ) );
NAND3_X1 _14696_ ( .A1(_05857_ ), .A2(\mtvec [27] ), .A3(_05644_ ), .ZN(_06707_ ) );
NAND3_X1 _14697_ ( .A1(_05852_ ), .A2(_06082_ ), .A3(_06707_ ), .ZN(_06708_ ) );
NAND3_X1 _14698_ ( .A1(_05861_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_05702_ ), .ZN(_06709_ ) );
OAI211_X1 _14699_ ( .A(_06083_ ), .B(_06709_ ), .C1(_05863_ ), .C2(_05864_ ), .ZN(_06710_ ) );
OAI21_X1 _14700_ ( .A(_06706_ ), .B1(_06708_ ), .B2(_06710_ ), .ZN(_06711_ ) );
AOI22_X1 _14701_ ( .A1(_05455_ ), .A2(_06140_ ), .B1(\ID_EX_typ [2] ), .B2(_06711_ ), .ZN(_06712_ ) );
OAI211_X1 _14702_ ( .A(_06712_ ), .B(_06497_ ), .C1(_06215_ ), .C2(\ID_EX_imm [27] ), .ZN(_06713_ ) );
OR3_X1 _14703_ ( .A1(_06711_ ), .A2(_06514_ ), .A3(_06490_ ), .ZN(_06714_ ) );
AND3_X1 _14704_ ( .A1(_03604_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_06715_ ) );
AOI21_X1 _14705_ ( .A(_06715_ ), .B1(_04722_ ), .B2(_06592_ ), .ZN(_06716_ ) );
OAI211_X1 _14706_ ( .A(_06713_ ), .B(_06714_ ), .C1(_06628_ ), .C2(_06716_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
OR3_X1 _14707_ ( .A1(_05844_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_05846_ ), .ZN(_06717_ ) );
NAND3_X1 _14708_ ( .A1(_05861_ ), .A2(\mtvec [26] ), .A3(_05678_ ), .ZN(_06718_ ) );
NAND3_X1 _14709_ ( .A1(_05856_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_05675_ ), .ZN(_06719_ ) );
AND2_X1 _14710_ ( .A1(_06718_ ), .A2(_06719_ ), .ZN(_06720_ ) );
NAND3_X1 _14711_ ( .A1(_06720_ ), .A2(_06109_ ), .A3(_06110_ ), .ZN(_06721_ ) );
OAI21_X1 _14712_ ( .A(_06717_ ), .B1(_06721_ ), .B2(_06233_ ), .ZN(_06722_ ) );
AOI22_X1 _14713_ ( .A1(_05351_ ), .A2(_06140_ ), .B1(\ID_EX_typ [2] ), .B2(_06722_ ), .ZN(_06723_ ) );
OAI211_X1 _14714_ ( .A(_06723_ ), .B(_06497_ ), .C1(_06215_ ), .C2(\ID_EX_imm [26] ), .ZN(_06724_ ) );
AND2_X1 _14715_ ( .A1(_06109_ ), .A2(_06110_ ), .ZN(_06725_ ) );
NAND3_X1 _14716_ ( .A1(_06674_ ), .A2(_06725_ ), .A3(_06720_ ), .ZN(_06726_ ) );
NAND4_X1 _14717_ ( .A1(_06726_ ), .A2(_06525_ ), .A3(_06717_ ), .A4(_06627_ ), .ZN(_06727_ ) );
AND3_X1 _14718_ ( .A1(_03604_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_06728_ ) );
AOI21_X1 _14719_ ( .A(_06728_ ), .B1(_04700_ ), .B2(_06592_ ), .ZN(_06729_ ) );
OAI211_X1 _14720_ ( .A(_06724_ ), .B(_06727_ ), .C1(_06628_ ), .C2(_06729_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
OR3_X1 _14721_ ( .A1(_05844_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_05846_ ), .ZN(_06730_ ) );
NAND3_X1 _14722_ ( .A1(_05861_ ), .A2(\mtvec [25] ), .A3(_05644_ ), .ZN(_06731_ ) );
NAND3_X1 _14723_ ( .A1(_05861_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_05702_ ), .ZN(_06732_ ) );
AND2_X1 _14724_ ( .A1(_06731_ ), .A2(_06732_ ), .ZN(_06733_ ) );
NAND3_X1 _14725_ ( .A1(_06733_ ), .A2(_06132_ ), .A3(_06133_ ), .ZN(_06734_ ) );
OAI21_X1 _14726_ ( .A(_06730_ ), .B1(_06734_ ), .B2(_06233_ ), .ZN(_06735_ ) );
AOI22_X1 _14727_ ( .A1(_06735_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_03210_ ), .ZN(_06736_ ) );
OAI211_X1 _14728_ ( .A(_06497_ ), .B(_06736_ ), .C1(_03184_ ), .C2(\ID_EX_typ [0] ), .ZN(_06737_ ) );
AND2_X1 _14729_ ( .A1(_06132_ ), .A2(_06133_ ), .ZN(_06738_ ) );
NAND3_X1 _14730_ ( .A1(_06674_ ), .A2(_06738_ ), .A3(_06733_ ), .ZN(_06739_ ) );
NAND4_X1 _14731_ ( .A1(_06739_ ), .A2(_06513_ ), .A3(_06730_ ), .A4(_06627_ ), .ZN(_06740_ ) );
AND3_X1 _14732_ ( .A1(_03604_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06741_ ) );
AOI21_X1 _14733_ ( .A(_06741_ ), .B1(_04676_ ), .B2(_06592_ ), .ZN(_06742_ ) );
OAI211_X1 _14734_ ( .A(_06737_ ), .B(_06740_ ), .C1(_06628_ ), .C2(_06742_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _14735_ ( .A(\ID_EX_typ [0] ), .B1(_02490_ ), .B2(_02509_ ), .ZN(_06743_ ) );
AND2_X1 _14736_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [24] ), .ZN(_06744_ ) );
OAI221_X1 _14737_ ( .A(_06627_ ), .B1(_06265_ ), .B2(_06156_ ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_06745_ ) );
NAND3_X1 _14738_ ( .A1(_05857_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_06063_ ), .ZN(_06746_ ) );
AND2_X1 _14739_ ( .A1(_06150_ ), .A2(_06746_ ), .ZN(_06747_ ) );
NAND4_X1 _14740_ ( .A1(_06747_ ), .A2(_05852_ ), .A3(_06659_ ), .A4(_06154_ ), .ZN(_06748_ ) );
NAND3_X1 _14741_ ( .A1(_05857_ ), .A2(\mtvec [24] ), .A3(_05679_ ), .ZN(_06749_ ) );
OAI21_X1 _14742_ ( .A(_06749_ ), .B1(_05863_ ), .B2(_05864_ ), .ZN(_06750_ ) );
OR2_X1 _14743_ ( .A1(_06748_ ), .A2(_06750_ ), .ZN(_06751_ ) );
OR3_X1 _14744_ ( .A1(_05863_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_05864_ ), .ZN(_06752_ ) );
NAND4_X1 _14745_ ( .A1(_06751_ ), .A2(_06513_ ), .A3(_06752_ ), .A4(_06627_ ), .ZN(_06753_ ) );
AND3_X1 _14746_ ( .A1(_03604_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_typ [7] ), .ZN(_06754_ ) );
AOI21_X1 _14747_ ( .A(_06754_ ), .B1(_04653_ ), .B2(_06592_ ), .ZN(_06755_ ) );
OAI211_X1 _14748_ ( .A(_06745_ ), .B(_06753_ ), .C1(_06628_ ), .C2(_06755_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
OR3_X1 _14749_ ( .A1(_05844_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_05846_ ), .ZN(_06756_ ) );
NAND3_X1 _14750_ ( .A1(_05861_ ), .A2(\mtvec [23] ), .A3(_05678_ ), .ZN(_06757_ ) );
NAND3_X1 _14751_ ( .A1(_05856_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_05702_ ), .ZN(_06758_ ) );
AND2_X1 _14752_ ( .A1(_06757_ ), .A2(_06758_ ), .ZN(_06759_ ) );
NAND3_X1 _14753_ ( .A1(_06759_ ), .A2(_06170_ ), .A3(_06171_ ), .ZN(_06760_ ) );
OAI21_X1 _14754_ ( .A(_06756_ ), .B1(_06760_ ), .B2(_06233_ ), .ZN(_06761_ ) );
AOI22_X1 _14755_ ( .A1(_05307_ ), .A2(_05661_ ), .B1(\ID_EX_typ [2] ), .B2(_06761_ ), .ZN(_06762_ ) );
OAI211_X1 _14756_ ( .A(_06762_ ), .B(_06497_ ), .C1(_06215_ ), .C2(\ID_EX_imm [23] ), .ZN(_06763_ ) );
OR3_X1 _14757_ ( .A1(_06761_ ), .A2(_06514_ ), .A3(_06490_ ), .ZN(_06764_ ) );
MUX2_X1 _14758_ ( .A(_06247_ ), .B(_04479_ ), .S(_06528_ ), .Z(_06765_ ) );
OAI211_X1 _14759_ ( .A(_06763_ ), .B(_06764_ ), .C1(_06628_ ), .C2(_06765_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
AOI21_X1 _14760_ ( .A(\ID_EX_typ [0] ), .B1(_02514_ ), .B2(_02534_ ), .ZN(_06766_ ) );
AND2_X1 _14761_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [22] ), .ZN(_06767_ ) );
OAI221_X1 _14762_ ( .A(_06627_ ), .B1(_06265_ ), .B2(_06186_ ), .C1(_06766_ ), .C2(_06767_ ), .ZN(_06768_ ) );
NAND3_X1 _14763_ ( .A1(_05857_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_06063_ ), .ZN(_06769_ ) );
AND2_X1 _14764_ ( .A1(_06180_ ), .A2(_06769_ ), .ZN(_06770_ ) );
NAND4_X1 _14765_ ( .A1(_06770_ ), .A2(_05852_ ), .A3(_06659_ ), .A4(_06184_ ), .ZN(_06771_ ) );
NAND3_X1 _14766_ ( .A1(_05857_ ), .A2(\mtvec [22] ), .A3(_05679_ ), .ZN(_06772_ ) );
OAI21_X1 _14767_ ( .A(_06772_ ), .B1(_05863_ ), .B2(_05864_ ), .ZN(_06773_ ) );
OR2_X1 _14768_ ( .A1(_06771_ ), .A2(_06773_ ), .ZN(_06774_ ) );
OR3_X1 _14769_ ( .A1(_05863_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_05864_ ), .ZN(_06775_ ) );
NAND4_X1 _14770_ ( .A1(_06774_ ), .A2(_06513_ ), .A3(_06775_ ), .A4(_06627_ ), .ZN(_06776_ ) );
MUX2_X1 _14771_ ( .A(_06187_ ), .B(_04454_ ), .S(_06519_ ), .Z(_06777_ ) );
OAI211_X1 _14772_ ( .A(_06768_ ), .B(_06776_ ), .C1(_06628_ ), .C2(_06777_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
AOI22_X1 _14773_ ( .A1(_05136_ ), .A2(_05661_ ), .B1(\ID_EX_typ [2] ), .B2(_06234_ ), .ZN(_06778_ ) );
OAI211_X1 _14774_ ( .A(_06778_ ), .B(_06497_ ), .C1(_06215_ ), .C2(\ID_EX_imm [31] ), .ZN(_06779_ ) );
OR3_X1 _14775_ ( .A1(_06234_ ), .A2(_06514_ ), .A3(_06490_ ), .ZN(_06780_ ) );
AND3_X1 _14776_ ( .A1(_03604_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06781_ ) );
AOI21_X1 _14777_ ( .A(_06781_ ), .B1(_04629_ ), .B2(_06592_ ), .ZN(_06782_ ) );
OAI211_X1 _14778_ ( .A(_06779_ ), .B(_06780_ ), .C1(_06628_ ), .C2(_06782_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
OR2_X1 _14779_ ( .A1(_06212_ ), .A2(_06502_ ), .ZN(_06783_ ) );
NOR3_X1 _14780_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06784_ ) );
AND2_X2 _14781_ ( .A1(\ID_EX_typ [3] ), .A2(\ID_EX_typ [2] ), .ZN(_06785_ ) );
AND2_X1 _14782_ ( .A1(_06784_ ), .A2(_06785_ ), .ZN(_06786_ ) );
INV_X1 _14783_ ( .A(_06786_ ), .ZN(_06787_ ) );
BUF_X4 _14784_ ( .A(_06787_ ), .Z(_06788_ ) );
NOR2_X1 _14785_ ( .A1(_06202_ ), .A2(_06788_ ), .ZN(_06789_ ) );
AND2_X1 _14786_ ( .A1(_02610_ ), .A2(_04503_ ), .ZN(_06790_ ) );
OAI21_X1 _14787_ ( .A(_05434_ ), .B1(_05425_ ), .B2(_04433_ ), .ZN(_06791_ ) );
AOI21_X1 _14788_ ( .A(_06790_ ), .B1(_06791_ ), .B2(_04504_ ), .ZN(_06792_ ) );
XNOR2_X1 _14789_ ( .A(_06792_ ), .B(_04529_ ), .ZN(_06793_ ) );
AND3_X1 _14790_ ( .A1(_04291_ ), .A2(\ID_EX_typ [3] ), .A3(_05127_ ), .ZN(_06794_ ) );
AND2_X2 _14791_ ( .A1(_06794_ ), .A2(_05144_ ), .ZN(_06795_ ) );
AND2_X1 _14792_ ( .A1(_06793_ ), .A2(_06795_ ), .ZN(_06796_ ) );
NOR3_X1 _14793_ ( .A1(_05125_ ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06797_ ) );
AND3_X1 _14794_ ( .A1(_06797_ ), .A2(\ID_EX_imm [21] ), .A3(_06785_ ), .ZN(_06798_ ) );
NOR3_X1 _14795_ ( .A1(_06789_ ), .A2(_06796_ ), .A3(_06798_ ), .ZN(_06799_ ) );
NOR2_X1 _14796_ ( .A1(_04149_ ), .A2(\ID_EX_typ [6] ), .ZN(_06800_ ) );
AND2_X1 _14797_ ( .A1(_06800_ ), .A2(_03605_ ), .ZN(_06801_ ) );
INV_X1 _14798_ ( .A(_06801_ ), .ZN(_06802_ ) );
BUF_X4 _14799_ ( .A(_06802_ ), .Z(_06803_ ) );
OAI21_X1 _14800_ ( .A(_06141_ ), .B1(_06799_ ), .B2(_06803_ ), .ZN(_06804_ ) );
INV_X1 _14801_ ( .A(_05116_ ), .ZN(_06805_ ) );
NOR2_X1 _14802_ ( .A1(_06805_ ), .A2(_05242_ ), .ZN(_06806_ ) );
INV_X1 _14803_ ( .A(_06806_ ), .ZN(_06807_ ) );
AND3_X1 _14804_ ( .A1(_02835_ ), .A2(_05235_ ), .A3(_05236_ ), .ZN(_06808_ ) );
AOI21_X1 _14805_ ( .A(_02835_ ), .B1(_05235_ ), .B2(_05236_ ), .ZN(_06809_ ) );
NOR3_X1 _14806_ ( .A1(_06807_ ), .A2(_06808_ ), .A3(_06809_ ), .ZN(_06810_ ) );
NOR2_X1 _14807_ ( .A1(_06810_ ), .A2(_06808_ ), .ZN(_06811_ ) );
NOR2_X1 _14808_ ( .A1(_06811_ ), .A2(_05246_ ), .ZN(_06812_ ) );
NOR2_X1 _14809_ ( .A1(_05230_ ), .A2(_05227_ ), .ZN(_06813_ ) );
OR3_X1 _14810_ ( .A1(_06812_ ), .A2(_05224_ ), .A3(_06813_ ), .ZN(_06814_ ) );
INV_X1 _14811_ ( .A(_05225_ ), .ZN(_06815_ ) );
AND4_X1 _14812_ ( .A1(_05256_ ), .A2(_05214_ ), .A3(_05260_ ), .A4(_05220_ ), .ZN(_06816_ ) );
NAND3_X1 _14813_ ( .A1(_06814_ ), .A2(_06815_ ), .A3(_06816_ ), .ZN(_06817_ ) );
INV_X1 _14814_ ( .A(_02788_ ), .ZN(_06818_ ) );
NOR2_X1 _14815_ ( .A1(_05259_ ), .A2(_06818_ ), .ZN(_06819_ ) );
AND2_X1 _14816_ ( .A1(_05214_ ), .A2(_05218_ ), .ZN(_06820_ ) );
AOI21_X1 _14817_ ( .A(_06820_ ), .B1(_02764_ ), .B2(_05212_ ), .ZN(_06821_ ) );
INV_X1 _14818_ ( .A(_06821_ ), .ZN(_06822_ ) );
AND2_X1 _14819_ ( .A1(_05260_ ), .A2(_05256_ ), .ZN(_06823_ ) );
AOI221_X4 _14820_ ( .A(_05264_ ), .B1(_05256_ ), .B2(_06819_ ), .C1(_06822_ ), .C2(_06823_ ), .ZN(_06824_ ) );
AND2_X1 _14821_ ( .A1(_06817_ ), .A2(_06824_ ), .ZN(_06825_ ) );
INV_X1 _14822_ ( .A(_06825_ ), .ZN(_06826_ ) );
AND2_X1 _14823_ ( .A1(_05182_ ), .A2(_05176_ ), .ZN(_06827_ ) );
AND3_X1 _14824_ ( .A1(_06827_ ), .A2(_05171_ ), .A3(_05166_ ), .ZN(_06828_ ) );
INV_X1 _14825_ ( .A(_05208_ ), .ZN(_06829_ ) );
NOR3_X1 _14826_ ( .A1(_06829_ ), .A2(_05202_ ), .A3(_05203_ ), .ZN(_06830_ ) );
AND3_X1 _14827_ ( .A1(_06830_ ), .A2(_05190_ ), .A3(_05195_ ), .ZN(_06831_ ) );
NAND3_X1 _14828_ ( .A1(_06826_ ), .A2(_06828_ ), .A3(_06831_ ), .ZN(_06832_ ) );
NAND3_X1 _14829_ ( .A1(_06827_ ), .A2(_05171_ ), .A3(_05166_ ), .ZN(_06833_ ) );
INV_X1 _14830_ ( .A(_05203_ ), .ZN(_06834_ ) );
NOR2_X1 _14831_ ( .A1(_05207_ ), .A2(_05278_ ), .ZN(_06835_ ) );
AOI21_X1 _14832_ ( .A(_05202_ ), .B1(_06834_ ), .B2(_06835_ ), .ZN(_06836_ ) );
OR4_X1 _14833_ ( .A1(_05188_ ), .A2(_06836_ ), .A3(_05189_ ), .A4(_05196_ ), .ZN(_06837_ ) );
INV_X1 _14834_ ( .A(_03095_ ), .ZN(_06838_ ) );
NOR2_X1 _14835_ ( .A1(_05194_ ), .A2(_06838_ ), .ZN(_06839_ ) );
AOI21_X1 _14836_ ( .A(_05188_ ), .B1(_05190_ ), .B2(_06839_ ), .ZN(_06840_ ) );
AOI21_X1 _14837_ ( .A(_06833_ ), .B1(_06837_ ), .B2(_06840_ ), .ZN(_06841_ ) );
NOR2_X1 _14838_ ( .A1(_05170_ ), .A2(_05411_ ), .ZN(_06842_ ) );
NOR2_X1 _14839_ ( .A1(_05181_ ), .A2(_06574_ ), .ZN(_06843_ ) );
NOR2_X1 _14840_ ( .A1(_05175_ ), .A2(_05270_ ), .ZN(_06844_ ) );
AOI21_X1 _14841_ ( .A(_06843_ ), .B1(_05182_ ), .B2(_06844_ ), .ZN(_06845_ ) );
NOR3_X1 _14842_ ( .A1(_06845_ ), .A2(_05172_ ), .A3(_05167_ ), .ZN(_06846_ ) );
INV_X1 _14843_ ( .A(_03020_ ), .ZN(_06847_ ) );
NOR2_X1 _14844_ ( .A1(_05165_ ), .A2(_06847_ ), .ZN(_06848_ ) );
INV_X1 _14845_ ( .A(_06848_ ), .ZN(_06849_ ) );
AND2_X1 _14846_ ( .A1(_05170_ ), .A2(_05411_ ), .ZN(_06850_ ) );
NOR3_X1 _14847_ ( .A1(_06849_ ), .A2(_06842_ ), .A3(_06850_ ), .ZN(_06851_ ) );
NOR4_X1 _14848_ ( .A1(_06841_ ), .A2(_06842_ ), .A3(_06846_ ), .A4(_06851_ ), .ZN(_06852_ ) );
AND2_X1 _14849_ ( .A1(_06832_ ), .A2(_06852_ ), .ZN(_06853_ ) );
AND2_X1 _14850_ ( .A1(_05318_ ), .A2(_05323_ ), .ZN(_06854_ ) );
AND3_X1 _14851_ ( .A1(_06854_ ), .A2(_05289_ ), .A3(_05293_ ), .ZN(_06855_ ) );
INV_X1 _14852_ ( .A(_06855_ ), .ZN(_06856_ ) );
OR2_X1 _14853_ ( .A1(_06853_ ), .A2(_06856_ ), .ZN(_06857_ ) );
INV_X1 _14854_ ( .A(_05338_ ), .ZN(_06858_ ) );
INV_X1 _14855_ ( .A(_02709_ ), .ZN(_06859_ ) );
NOR2_X1 _14856_ ( .A1(_05292_ ), .A2(_06859_ ), .ZN(_06860_ ) );
AOI21_X1 _14857_ ( .A(_05339_ ), .B1(_06858_ ), .B2(_06860_ ), .ZN(_06861_ ) );
NOR3_X1 _14858_ ( .A1(_06861_ ), .A2(_05319_ ), .A3(_05324_ ), .ZN(_06862_ ) );
INV_X1 _14859_ ( .A(_04380_ ), .ZN(_06863_ ) );
NOR2_X1 _14860_ ( .A1(_05322_ ), .A2(_06863_ ), .ZN(_06864_ ) );
AND2_X1 _14861_ ( .A1(_05322_ ), .A2(_06863_ ), .ZN(_06865_ ) );
NOR4_X1 _14862_ ( .A1(_06865_ ), .A2(_06864_ ), .A3(_06538_ ), .A4(_05317_ ), .ZN(_06866_ ) );
NOR3_X1 _14863_ ( .A1(_06862_ ), .A2(_06864_ ), .A3(_06866_ ), .ZN(_06867_ ) );
AND2_X1 _14864_ ( .A1(_06857_ ), .A2(_06867_ ), .ZN(_06868_ ) );
INV_X1 _14865_ ( .A(_06868_ ), .ZN(_06869_ ) );
NAND2_X1 _14866_ ( .A1(_06869_ ), .A2(_05314_ ), .ZN(_06870_ ) );
NOR2_X1 _14867_ ( .A1(_05331_ ), .A2(_05313_ ), .ZN(_06871_ ) );
INV_X1 _14868_ ( .A(_06871_ ), .ZN(_06872_ ) );
AOI21_X1 _14869_ ( .A(_05303_ ), .B1(_06870_ ), .B2(_06872_ ), .ZN(_06873_ ) );
AOI211_X1 _14870_ ( .A(_05302_ ), .B(_06871_ ), .C1(_06869_ ), .C2(_05314_ ), .ZN(_06874_ ) );
BUF_X4 _14871_ ( .A(_05124_ ), .Z(_06875_ ) );
NOR2_X1 _14872_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06876_ ) );
INV_X1 _14873_ ( .A(_06876_ ), .ZN(_06877_ ) );
NOR2_X2 _14874_ ( .A1(_06875_ ), .A2(_06877_ ), .ZN(_06878_ ) );
INV_X1 _14875_ ( .A(_06878_ ), .ZN(_06879_ ) );
BUF_X2 _14876_ ( .A(_06879_ ), .Z(_06880_ ) );
OR3_X1 _14877_ ( .A1(_06873_ ), .A2(_06874_ ), .A3(_06880_ ), .ZN(_06881_ ) );
AND2_X2 _14878_ ( .A1(_05466_ ), .A2(\ID_EX_typ [2] ), .ZN(_06882_ ) );
BUF_X4 _14879_ ( .A(_06882_ ), .Z(_06883_ ) );
BUF_X4 _14880_ ( .A(_06883_ ), .Z(_06884_ ) );
OR2_X1 _14881_ ( .A1(_05259_ ), .A2(_05255_ ), .ZN(_06885_ ) );
AND2_X1 _14882_ ( .A1(_05237_ ), .A2(_05242_ ), .ZN(_06886_ ) );
AND2_X2 _14883_ ( .A1(_06886_ ), .A2(_05230_ ), .ZN(_06887_ ) );
AND2_X1 _14884_ ( .A1(_06887_ ), .A2(_05233_ ), .ZN(_06888_ ) );
AOI221_X4 _14885_ ( .A(_06885_ ), .B1(_05210_ ), .B2(_05211_ ), .C1(_06888_ ), .C2(_05217_ ), .ZN(_06889_ ) );
AND4_X1 _14886_ ( .A1(_05255_ ), .A2(_05212_ ), .A3(_05259_ ), .A4(_05217_ ), .ZN(_06890_ ) );
NAND4_X1 _14887_ ( .A1(_06890_ ), .A2(_05233_ ), .A3(_05230_ ), .A4(_06886_ ), .ZN(_06891_ ) );
NAND4_X1 _14888_ ( .A1(_05259_ ), .A2(_05255_ ), .A3(_05210_ ), .A4(_05211_ ), .ZN(_06892_ ) );
NAND2_X1 _14889_ ( .A1(_06891_ ), .A2(_06892_ ), .ZN(_06893_ ) );
OAI21_X1 _14890_ ( .A(_03243_ ), .B1(_06889_ ), .B2(_06893_ ), .ZN(_06894_ ) );
AND3_X1 _14891_ ( .A1(_05207_ ), .A2(_05199_ ), .A3(_05198_ ), .ZN(_06895_ ) );
AND2_X1 _14892_ ( .A1(_06893_ ), .A2(_06895_ ), .ZN(_06896_ ) );
INV_X1 _14893_ ( .A(_06896_ ), .ZN(_06897_ ) );
OR3_X1 _14894_ ( .A1(_06893_ ), .A2(_05200_ ), .A3(_05207_ ), .ZN(_06898_ ) );
AOI21_X1 _14895_ ( .A(_06894_ ), .B1(_06897_ ), .B2(_06898_ ), .ZN(_06899_ ) );
NAND3_X1 _14896_ ( .A1(_06893_ ), .A2(_05194_ ), .A3(_06895_ ), .ZN(_06900_ ) );
NOR2_X1 _14897_ ( .A1(_06900_ ), .A2(_05277_ ), .ZN(_06901_ ) );
AOI211_X1 _14898_ ( .A(_05186_ ), .B(_05194_ ), .C1(_06893_ ), .C2(_06895_ ), .ZN(_06902_ ) );
OAI21_X1 _14899_ ( .A(_06899_ ), .B1(_06901_ ), .B2(_06902_ ), .ZN(_06903_ ) );
NOR4_X1 _14900_ ( .A1(_05306_ ), .A2(_05301_ ), .A3(_05313_ ), .A4(_05296_ ), .ZN(_06904_ ) );
NOR4_X1 _14901_ ( .A1(_05170_ ), .A2(_05165_ ), .A3(_05181_ ), .A4(_05175_ ), .ZN(_06905_ ) );
OR2_X1 _14902_ ( .A1(_05322_ ), .A2(_05317_ ), .ZN(_06906_ ) );
NOR3_X1 _14903_ ( .A1(_06906_ ), .A2(_05288_ ), .A3(_05292_ ), .ZN(_06907_ ) );
AND3_X1 _14904_ ( .A1(_06904_ ), .A2(_06905_ ), .A3(_06907_ ), .ZN(_06908_ ) );
NOR4_X1 _14905_ ( .A1(_05350_ ), .A2(_05362_ ), .A3(_05357_ ), .A4(_05370_ ), .ZN(_06909_ ) );
AND4_X1 _14906_ ( .A1(_05153_ ), .A2(_05386_ ), .A3(_05159_ ), .A4(_05147_ ), .ZN(_06910_ ) );
NAND3_X1 _14907_ ( .A1(_06908_ ), .A2(_06909_ ), .A3(_06910_ ), .ZN(_06911_ ) );
NOR2_X1 _14908_ ( .A1(_06901_ ), .A2(_06911_ ), .ZN(_06912_ ) );
AND2_X1 _14909_ ( .A1(_05170_ ), .A2(_05165_ ), .ZN(_06913_ ) );
AND3_X1 _14910_ ( .A1(_06913_ ), .A2(_05181_ ), .A3(_05175_ ), .ZN(_06914_ ) );
AOI21_X1 _14911_ ( .A(_06912_ ), .B1(_06914_ ), .B2(_06901_ ), .ZN(_06915_ ) );
NOR2_X1 _14912_ ( .A1(_06903_ ), .A2(_06915_ ), .ZN(_06916_ ) );
NOR4_X1 _14913_ ( .A1(_05386_ ), .A2(_05159_ ), .A3(_05153_ ), .A4(_05147_ ), .ZN(_06917_ ) );
AOI22_X1 _14914_ ( .A1(_05348_ ), .A2(_05349_ ), .B1(_05355_ ), .B2(_05356_ ), .ZN(_06918_ ) );
AND4_X1 _14915_ ( .A1(_05362_ ), .A2(_06917_ ), .A3(_05370_ ), .A4(_06918_ ), .ZN(_06919_ ) );
AND4_X1 _14916_ ( .A1(_05321_ ), .A2(_05320_ ), .A3(_05315_ ), .A4(_05316_ ), .ZN(_06920_ ) );
AND3_X1 _14917_ ( .A1(_06920_ ), .A2(_05288_ ), .A3(_05292_ ), .ZN(_06921_ ) );
AND2_X1 _14918_ ( .A1(_05301_ ), .A2(_05313_ ), .ZN(_06922_ ) );
AND4_X1 _14919_ ( .A1(_05305_ ), .A2(_06922_ ), .A3(_05304_ ), .A4(_05296_ ), .ZN(_06923_ ) );
NAND3_X1 _14920_ ( .A1(_06919_ ), .A2(_06921_ ), .A3(_06923_ ), .ZN(_06924_ ) );
NAND3_X1 _14921_ ( .A1(_06924_ ), .A2(_06914_ ), .A3(_06901_ ), .ZN(_06925_ ) );
AND2_X2 _14922_ ( .A1(_06916_ ), .A2(_06925_ ), .ZN(_06926_ ) );
AND2_X1 _14923_ ( .A1(_06888_ ), .A2(_05217_ ), .ZN(_06927_ ) );
XNOR2_X1 _14924_ ( .A(_06927_ ), .B(_05212_ ), .ZN(_06928_ ) );
AND2_X2 _14925_ ( .A1(_06926_ ), .A2(_06928_ ), .ZN(_06929_ ) );
XNOR2_X1 _14926_ ( .A(_06888_ ), .B(_05217_ ), .ZN(_06930_ ) );
NOR2_X1 _14927_ ( .A1(_06930_ ), .A2(_05212_ ), .ZN(_06931_ ) );
NOR2_X1 _14928_ ( .A1(_06929_ ), .A2(_06931_ ), .ZN(_06932_ ) );
BUF_X2 _14929_ ( .A(_06926_ ), .Z(_06933_ ) );
XNOR2_X1 _14930_ ( .A(_06887_ ), .B(_05223_ ), .ZN(_06934_ ) );
INV_X1 _14931_ ( .A(_06934_ ), .ZN(_06935_ ) );
NAND2_X1 _14932_ ( .A1(_06933_ ), .A2(_06935_ ), .ZN(_06936_ ) );
BUF_X4 _14933_ ( .A(_05237_ ), .Z(_06937_ ) );
BUF_X4 _14934_ ( .A(_06937_ ), .Z(_06938_ ) );
BUF_X4 _14935_ ( .A(_06938_ ), .Z(_06939_ ) );
BUF_X4 _14936_ ( .A(_05242_ ), .Z(_06940_ ) );
BUF_X4 _14937_ ( .A(_06940_ ), .Z(_06941_ ) );
XNOR2_X1 _14938_ ( .A(_06939_ ), .B(_06941_ ), .ZN(_06942_ ) );
BUF_X4 _14939_ ( .A(_05231_ ), .Z(_06943_ ) );
BUF_X2 _14940_ ( .A(_06943_ ), .Z(_06944_ ) );
NOR2_X1 _14941_ ( .A1(_06942_ ), .A2(_06944_ ), .ZN(_06945_ ) );
NOR2_X1 _14942_ ( .A1(_06936_ ), .A2(_06945_ ), .ZN(_06946_ ) );
INV_X1 _14943_ ( .A(_06946_ ), .ZN(_06947_ ) );
INV_X1 _14944_ ( .A(_06930_ ), .ZN(_06948_ ) );
AOI21_X1 _14945_ ( .A(_06932_ ), .B1(_06947_ ), .B2(_06948_ ), .ZN(_06949_ ) );
BUF_X4 _14946_ ( .A(_05230_ ), .Z(_06950_ ) );
BUF_X4 _14947_ ( .A(_06950_ ), .Z(_06951_ ) );
AND3_X1 _14948_ ( .A1(_06940_ ), .A2(_03183_ ), .A3(_03163_ ), .ZN(_06952_ ) );
BUF_X2 _14949_ ( .A(_05242_ ), .Z(_06953_ ) );
BUF_X2 _14950_ ( .A(_06953_ ), .Z(_06954_ ) );
NOR2_X1 _14951_ ( .A1(_03207_ ), .A2(_06954_ ), .ZN(_06955_ ) );
OAI21_X1 _14952_ ( .A(_06938_ ), .B1(_06952_ ), .B2(_06955_ ), .ZN(_06956_ ) );
INV_X1 _14953_ ( .A(_05237_ ), .ZN(_06957_ ) );
BUF_X4 _14954_ ( .A(_06957_ ), .Z(_06958_ ) );
NOR2_X1 _14955_ ( .A1(_02448_ ), .A2(_06954_ ), .ZN(_06959_ ) );
BUF_X4 _14956_ ( .A(_05240_ ), .Z(_06960_ ) );
BUF_X4 _14957_ ( .A(_05241_ ), .Z(_06961_ ) );
AOI21_X1 _14958_ ( .A(_02487_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_06962_ ) );
OAI21_X1 _14959_ ( .A(_06958_ ), .B1(_06959_ ), .B2(_06962_ ), .ZN(_06963_ ) );
AOI21_X1 _14960_ ( .A(_06951_ ), .B1(_06956_ ), .B2(_06963_ ), .ZN(_06964_ ) );
BUF_X4 _14961_ ( .A(_05231_ ), .Z(_06965_ ) );
NOR2_X1 _14962_ ( .A1(_02535_ ), .A2(_06954_ ), .ZN(_06966_ ) );
AOI21_X1 _14963_ ( .A(_04505_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_06967_ ) );
OAI21_X1 _14964_ ( .A(_06938_ ), .B1(_06966_ ), .B2(_06967_ ), .ZN(_06968_ ) );
BUF_X4 _14965_ ( .A(_06957_ ), .Z(_06969_ ) );
NOR2_X1 _14966_ ( .A1(_02510_ ), .A2(_06954_ ), .ZN(_06970_ ) );
AOI21_X1 _14967_ ( .A(_02561_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_06971_ ) );
OAI21_X1 _14968_ ( .A(_06969_ ), .B1(_06970_ ), .B2(_06971_ ), .ZN(_06972_ ) );
AOI21_X1 _14969_ ( .A(_06965_ ), .B1(_06968_ ), .B2(_06972_ ), .ZN(_06973_ ) );
NOR2_X1 _14970_ ( .A1(_06964_ ), .A2(_06973_ ), .ZN(_06974_ ) );
INV_X2 _14971_ ( .A(_05242_ ), .ZN(_06975_ ) );
NAND3_X1 _14972_ ( .A1(_06975_ ), .A2(_02399_ ), .A3(_02400_ ), .ZN(_06976_ ) );
NAND3_X1 _14973_ ( .A1(_06953_ ), .A2(_02424_ ), .A3(_02423_ ), .ZN(_06977_ ) );
AND3_X1 _14974_ ( .A1(_06976_ ), .A2(_06937_ ), .A3(_06977_ ), .ZN(_06978_ ) );
AND2_X1 _14975_ ( .A1(_03243_ ), .A2(_06954_ ), .ZN(_06979_ ) );
AOI21_X1 _14976_ ( .A(_06978_ ), .B1(_06958_ ), .B2(_06979_ ), .ZN(_06980_ ) );
BUF_X2 _14977_ ( .A(_06965_ ), .Z(_06981_ ) );
NOR2_X1 _14978_ ( .A1(_06980_ ), .A2(_06981_ ), .ZN(_06982_ ) );
BUF_X4 _14979_ ( .A(_05223_ ), .Z(_06983_ ) );
BUF_X4 _14980_ ( .A(_06983_ ), .Z(_06984_ ) );
MUX2_X1 _14981_ ( .A(_06974_ ), .B(_06982_ ), .S(_06984_ ), .Z(_06985_ ) );
CLKBUF_X3 _14982_ ( .A(_05217_ ), .Z(_06986_ ) );
BUF_X2 _14983_ ( .A(_06986_ ), .Z(_06987_ ) );
BUF_X2 _14984_ ( .A(_06987_ ), .Z(_06988_ ) );
AND2_X1 _14985_ ( .A1(_06985_ ), .A2(_06988_ ), .ZN(_06989_ ) );
OAI21_X1 _14986_ ( .A(_06884_ ), .B1(_06949_ ), .B2(_06989_ ), .ZN(_06990_ ) );
AND2_X1 _14987_ ( .A1(_05126_ ), .A2(\ID_EX_typ [2] ), .ZN(_06991_ ) );
BUF_X4 _14988_ ( .A(_06991_ ), .Z(_06992_ ) );
BUF_X4 _14989_ ( .A(_06992_ ), .Z(_06993_ ) );
NAND3_X1 _14990_ ( .A1(_06985_ ), .A2(_06988_ ), .A3(_06993_ ), .ZN(_06994_ ) );
BUF_X2 _14991_ ( .A(_05217_ ), .Z(_06995_ ) );
BUF_X2 _14992_ ( .A(_06995_ ), .Z(_06996_ ) );
AOI21_X1 _14993_ ( .A(_03068_ ), .B1(_05240_ ), .B2(_05241_ ), .ZN(_06997_ ) );
NOR2_X1 _14994_ ( .A1(_06953_ ), .A2(_03045_ ), .ZN(_06998_ ) );
NOR3_X1 _14995_ ( .A1(_06969_ ), .A2(_06997_ ), .A3(_06998_ ), .ZN(_06999_ ) );
AOI21_X1 _14996_ ( .A(_02812_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_07000_ ) );
NOR2_X1 _14997_ ( .A1(_06953_ ), .A2(_02788_ ), .ZN(_07001_ ) );
NOR3_X1 _14998_ ( .A1(_07000_ ), .A2(_07001_ ), .A3(_06937_ ), .ZN(_07002_ ) );
NOR2_X1 _14999_ ( .A1(_06999_ ), .A2(_07002_ ), .ZN(_07003_ ) );
BUF_X4 _15000_ ( .A(_06950_ ), .Z(_07004_ ) );
BUF_X4 _15001_ ( .A(_07004_ ), .Z(_07005_ ) );
BUF_X2 _15002_ ( .A(_07005_ ), .Z(_07006_ ) );
NOR2_X1 _15003_ ( .A1(_07003_ ), .A2(_07006_ ), .ZN(_07007_ ) );
BUF_X4 _15004_ ( .A(_05233_ ), .Z(_07008_ ) );
BUF_X4 _15005_ ( .A(_07008_ ), .Z(_07009_ ) );
BUF_X4 _15006_ ( .A(_07009_ ), .Z(_07010_ ) );
BUF_X4 _15007_ ( .A(_06969_ ), .Z(_07011_ ) );
BUF_X4 _15008_ ( .A(_06960_ ), .Z(_07012_ ) );
BUF_X4 _15009_ ( .A(_06961_ ), .Z(_07013_ ) );
AOI21_X1 _15010_ ( .A(_04781_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07014_ ) );
BUF_X4 _15011_ ( .A(_06940_ ), .Z(_07015_ ) );
NOR2_X1 _15012_ ( .A1(_07015_ ), .A2(_02948_ ), .ZN(_07016_ ) );
OR3_X1 _15013_ ( .A1(_07011_ ), .A2(_07014_ ), .A3(_07016_ ), .ZN(_07017_ ) );
AOI21_X1 _15014_ ( .A(_04854_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07018_ ) );
NOR2_X1 _15015_ ( .A1(_07015_ ), .A2(_03095_ ), .ZN(_07019_ ) );
BUF_X2 _15016_ ( .A(_06937_ ), .Z(_07020_ ) );
OR3_X1 _15017_ ( .A1(_07018_ ), .A2(_07019_ ), .A3(_07020_ ), .ZN(_07021_ ) );
AOI21_X1 _15018_ ( .A(_06981_ ), .B1(_07017_ ), .B2(_07021_ ), .ZN(_07022_ ) );
NOR3_X1 _15019_ ( .A1(_07007_ ), .A2(_07010_ ), .A3(_07022_ ), .ZN(_07023_ ) );
BUF_X4 _15020_ ( .A(_06951_ ), .Z(_07024_ ) );
BUF_X2 _15021_ ( .A(_06969_ ), .Z(_07025_ ) );
AOI21_X1 _15022_ ( .A(_02684_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_07026_ ) );
NOR2_X1 _15023_ ( .A1(_07015_ ), .A2(_02709_ ), .ZN(_07027_ ) );
OR3_X1 _15024_ ( .A1(_07025_ ), .A2(_07026_ ), .A3(_07027_ ), .ZN(_07028_ ) );
AOI21_X1 _15025_ ( .A(_02996_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07029_ ) );
NOR2_X1 _15026_ ( .A1(_07015_ ), .A2(_03020_ ), .ZN(_07030_ ) );
OR3_X1 _15027_ ( .A1(_07029_ ), .A2(_07030_ ), .A3(_07020_ ), .ZN(_07031_ ) );
AOI21_X1 _15028_ ( .A(_07024_ ), .B1(_07028_ ), .B2(_07031_ ), .ZN(_07032_ ) );
BUF_X4 _15029_ ( .A(_06939_ ), .Z(_07033_ ) );
NOR2_X1 _15030_ ( .A1(_02610_ ), .A2(_06940_ ), .ZN(_07034_ ) );
OAI21_X1 _15031_ ( .A(_07033_ ), .B1(_07034_ ), .B2(_06967_ ), .ZN(_07035_ ) );
BUF_X4 _15032_ ( .A(_07011_ ), .Z(_07036_ ) );
NOR2_X1 _15033_ ( .A1(_02635_ ), .A2(_06940_ ), .ZN(_07037_ ) );
AOI21_X1 _15034_ ( .A(_04380_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_07038_ ) );
OAI21_X1 _15035_ ( .A(_07036_ ), .B1(_07037_ ), .B2(_07038_ ), .ZN(_07039_ ) );
BUF_X2 _15036_ ( .A(_07004_ ), .Z(_07040_ ) );
AND3_X1 _15037_ ( .A1(_07035_ ), .A2(_07039_ ), .A3(_07040_ ), .ZN(_07041_ ) );
BUF_X4 _15038_ ( .A(_06984_ ), .Z(_07042_ ) );
NOR3_X1 _15039_ ( .A1(_07032_ ), .A2(_07041_ ), .A3(_07042_ ), .ZN(_07043_ ) );
OAI21_X1 _15040_ ( .A(_06996_ ), .B1(_07023_ ), .B2(_07043_ ), .ZN(_07044_ ) );
INV_X1 _15041_ ( .A(_05464_ ), .ZN(_07045_ ) );
AND3_X1 _15042_ ( .A1(_06953_ ), .A2(_02908_ ), .A3(_02909_ ), .ZN(_07046_ ) );
NOR2_X1 _15043_ ( .A1(_06940_ ), .A2(_02886_ ), .ZN(_07047_ ) );
NOR3_X1 _15044_ ( .A1(_07046_ ), .A2(_06937_ ), .A3(_07047_ ), .ZN(_07048_ ) );
AOI21_X1 _15045_ ( .A(_02764_ ), .B1(_05240_ ), .B2(_05241_ ), .ZN(_07049_ ) );
NOR2_X1 _15046_ ( .A1(_06953_ ), .A2(_02735_ ), .ZN(_07050_ ) );
NOR3_X1 _15047_ ( .A1(_06969_ ), .A2(_07049_ ), .A3(_07050_ ), .ZN(_07051_ ) );
NOR2_X1 _15048_ ( .A1(_07048_ ), .A2(_07051_ ), .ZN(_07052_ ) );
NAND2_X1 _15049_ ( .A1(_07052_ ), .A2(_07006_ ), .ZN(_07053_ ) );
BUF_X2 _15050_ ( .A(_07008_ ), .Z(_07054_ ) );
BUF_X2 _15051_ ( .A(_07054_ ), .Z(_07055_ ) );
AND3_X1 _15052_ ( .A1(_06954_ ), .A2(_02834_ ), .A3(_02815_ ), .ZN(_07056_ ) );
NOR3_X1 _15053_ ( .A1(_07056_ ), .A2(_06958_ ), .A3(_05243_ ), .ZN(_07057_ ) );
OR2_X1 _15054_ ( .A1(_07057_ ), .A2(_07040_ ), .ZN(_07058_ ) );
NAND3_X1 _15055_ ( .A1(_07053_ ), .A2(_07055_ ), .A3(_07058_ ), .ZN(_07059_ ) );
BUF_X4 _15056_ ( .A(_05250_ ), .Z(_07060_ ) );
BUF_X4 _15057_ ( .A(_07060_ ), .Z(_07061_ ) );
AOI21_X1 _15058_ ( .A(_07045_ ), .B1(_07059_ ), .B2(_07061_ ), .ZN(_07062_ ) );
NAND2_X1 _15059_ ( .A1(_07044_ ), .A2(_07062_ ), .ZN(_07063_ ) );
INV_X1 _15060_ ( .A(_04505_ ), .ZN(_07064_ ) );
INV_X1 _15061_ ( .A(_06875_ ), .ZN(_07065_ ) );
OR3_X1 _15062_ ( .A1(_05301_ ), .A2(_07064_ ), .A3(_07065_ ), .ZN(_07066_ ) );
AOI21_X1 _15063_ ( .A(_05130_ ), .B1(_05301_ ), .B2(_07064_ ), .ZN(_07067_ ) );
BUF_X2 _15064_ ( .A(_05467_ ), .Z(_07068_ ) );
AOI21_X1 _15065_ ( .A(_07067_ ), .B1(_05302_ ), .B2(_07068_ ), .ZN(_07069_ ) );
AND4_X1 _15066_ ( .A1(_06994_ ), .A2(_07063_ ), .A3(_07066_ ), .A4(_07069_ ), .ZN(_07070_ ) );
NAND3_X1 _15067_ ( .A1(_06881_ ), .A2(_06990_ ), .A3(_07070_ ), .ZN(_07071_ ) );
OAI21_X1 _15068_ ( .A(_06785_ ), .B1(_06797_ ), .B2(_06784_ ), .ZN(_07072_ ) );
NOR2_X1 _15069_ ( .A1(_05481_ ), .A2(\ID_EX_typ [2] ), .ZN(_07073_ ) );
OAI211_X1 _15070_ ( .A(_07073_ ), .B(_05125_ ), .C1(_05144_ ), .C2(_04146_ ), .ZN(_07074_ ) );
AND2_X1 _15071_ ( .A1(_07072_ ), .A2(_07074_ ), .ZN(_07075_ ) );
NOR2_X1 _15072_ ( .A1(_07075_ ), .A2(_06802_ ), .ZN(_07076_ ) );
INV_X2 _15073_ ( .A(_07076_ ), .ZN(_07077_ ) );
BUF_X4 _15074_ ( .A(_07077_ ), .Z(_07078_ ) );
AOI21_X1 _15075_ ( .A(_06804_ ), .B1(_07071_ ), .B2(_07078_ ), .ZN(_07079_ ) );
BUF_X4 _15076_ ( .A(_06491_ ), .Z(_07080_ ) );
OAI21_X1 _15077_ ( .A(_07080_ ), .B1(_06198_ ), .B2(_05921_ ), .ZN(_07081_ ) );
OAI21_X1 _15078_ ( .A(_06783_ ), .B1(_07079_ ), .B2(_07081_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
NAND2_X1 _15079_ ( .A1(_05614_ ), .A2(_06494_ ), .ZN(_07082_ ) );
BUF_X4 _15080_ ( .A(_06786_ ), .Z(_07083_ ) );
BUF_X2 _15081_ ( .A(_07083_ ), .Z(_07084_ ) );
AND2_X1 _15082_ ( .A1(_06797_ ), .A2(_06785_ ), .ZN(_07085_ ) );
BUF_X4 _15083_ ( .A(_07085_ ), .Z(_07086_ ) );
BUF_X4 _15084_ ( .A(_07086_ ), .Z(_07087_ ) );
AOI22_X1 _15085_ ( .A1(_05617_ ), .A2(_07084_ ), .B1(\ID_EX_imm [20] ), .B2(_07087_ ), .ZN(_07088_ ) );
INV_X1 _15086_ ( .A(_06795_ ), .ZN(_07089_ ) );
AOI21_X1 _15087_ ( .A(_07089_ ), .B1(_06791_ ), .B2(_04504_ ), .ZN(_07090_ ) );
OAI21_X1 _15088_ ( .A(_07090_ ), .B1(_04504_ ), .B2(_06791_ ), .ZN(_07091_ ) );
AOI21_X1 _15089_ ( .A(_06803_ ), .B1(_07088_ ), .B2(_07091_ ), .ZN(_07092_ ) );
OR2_X1 _15090_ ( .A1(_07092_ ), .A2(_05838_ ), .ZN(_07093_ ) );
AOI21_X1 _15091_ ( .A(_06880_ ), .B1(_06869_ ), .B2(_05314_ ), .ZN(_07094_ ) );
OAI21_X1 _15092_ ( .A(_07094_ ), .B1(_05314_ ), .B2(_06869_ ), .ZN(_07095_ ) );
INV_X1 _15093_ ( .A(_06929_ ), .ZN(_07096_ ) );
INV_X1 _15094_ ( .A(_06931_ ), .ZN(_07097_ ) );
AOI21_X1 _15095_ ( .A(_06944_ ), .B1(_07033_ ), .B2(_06941_ ), .ZN(_07098_ ) );
INV_X1 _15096_ ( .A(_07098_ ), .ZN(_07099_ ) );
NAND3_X1 _15097_ ( .A1(_06933_ ), .A2(_06935_ ), .A3(_07099_ ), .ZN(_07100_ ) );
AOI22_X1 _15098_ ( .A1(_07096_ ), .A2(_07097_ ), .B1(_06948_ ), .B2(_07100_ ), .ZN(_07101_ ) );
AND3_X1 _15099_ ( .A1(_06953_ ), .A2(_02490_ ), .A3(_02509_ ), .ZN(_07102_ ) );
NOR2_X1 _15100_ ( .A1(_03184_ ), .A2(_06940_ ), .ZN(_07103_ ) );
NOR2_X1 _15101_ ( .A1(_07102_ ), .A2(_07103_ ), .ZN(_07104_ ) );
NOR2_X1 _15102_ ( .A1(_07104_ ), .A2(_06969_ ), .ZN(_07105_ ) );
AND3_X1 _15103_ ( .A1(_06953_ ), .A2(_03187_ ), .A3(_03206_ ), .ZN(_07106_ ) );
INV_X1 _15104_ ( .A(_07106_ ), .ZN(_07107_ ) );
NAND3_X1 _15105_ ( .A1(_05455_ ), .A2(_06960_ ), .A3(_06961_ ), .ZN(_07108_ ) );
AOI21_X1 _15106_ ( .A(_06937_ ), .B1(_07107_ ), .B2(_07108_ ), .ZN(_07109_ ) );
OR3_X1 _15107_ ( .A1(_07105_ ), .A2(_07109_ ), .A3(_05230_ ), .ZN(_07110_ ) );
AND3_X1 _15108_ ( .A1(_06940_ ), .A2(_02589_ ), .A3(_02609_ ), .ZN(_07111_ ) );
NOR2_X1 _15109_ ( .A1(_06954_ ), .A2(_04505_ ), .ZN(_07112_ ) );
OAI21_X1 _15110_ ( .A(_06938_ ), .B1(_07111_ ), .B2(_07112_ ), .ZN(_07113_ ) );
AND3_X1 _15111_ ( .A1(_06940_ ), .A2(_02514_ ), .A3(_02534_ ), .ZN(_07114_ ) );
NOR2_X1 _15112_ ( .A1(_06940_ ), .A2(_02561_ ), .ZN(_07115_ ) );
OAI21_X1 _15113_ ( .A(_06958_ ), .B1(_07114_ ), .B2(_07115_ ), .ZN(_07116_ ) );
NAND3_X1 _15114_ ( .A1(_07113_ ), .A2(_07116_ ), .A3(_06950_ ), .ZN(_07117_ ) );
NAND2_X1 _15115_ ( .A1(_07110_ ), .A2(_07117_ ), .ZN(_07118_ ) );
NAND3_X1 _15116_ ( .A1(_06975_ ), .A2(_02424_ ), .A3(_02423_ ), .ZN(_07119_ ) );
NAND3_X1 _15117_ ( .A1(_06953_ ), .A2(_02447_ ), .A3(_02428_ ), .ZN(_07120_ ) );
AND2_X1 _15118_ ( .A1(_07119_ ), .A2(_07120_ ), .ZN(_07121_ ) );
AND3_X1 _15119_ ( .A1(_02399_ ), .A2(_02400_ ), .A3(_06953_ ), .ZN(_07122_ ) );
AOI21_X1 _15120_ ( .A(_07122_ ), .B1(_05136_ ), .B2(_06975_ ), .ZN(_07123_ ) );
MUX2_X1 _15121_ ( .A(_07121_ ), .B(_07123_ ), .S(_06969_ ), .Z(_07124_ ) );
AND2_X1 _15122_ ( .A1(_07124_ ), .A2(_07004_ ), .ZN(_07125_ ) );
MUX2_X1 _15123_ ( .A(_07118_ ), .B(_07125_ ), .S(_06983_ ), .Z(_07126_ ) );
AND2_X1 _15124_ ( .A1(_07126_ ), .A2(_06988_ ), .ZN(_07127_ ) );
OAI21_X1 _15125_ ( .A(_06884_ ), .B1(_07101_ ), .B2(_07127_ ), .ZN(_07128_ ) );
BUF_X4 _15126_ ( .A(_05130_ ), .Z(_07129_ ) );
BUF_X4 _15127_ ( .A(_07129_ ), .Z(_07130_ ) );
AOI21_X1 _15128_ ( .A(_07130_ ), .B1(_05331_ ), .B2(_05313_ ), .ZN(_07131_ ) );
NOR2_X1 _15129_ ( .A1(_02910_ ), .A2(_06941_ ), .ZN(_07132_ ) );
AOI21_X1 _15130_ ( .A(_02735_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07133_ ) );
NOR3_X1 _15131_ ( .A1(_07132_ ), .A2(_07025_ ), .A3(_07133_ ), .ZN(_07134_ ) );
NOR2_X1 _15132_ ( .A1(_02835_ ), .A2(_07015_ ), .ZN(_07135_ ) );
AOI21_X1 _15133_ ( .A(_02886_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_07136_ ) );
BUF_X2 _15134_ ( .A(_06937_ ), .Z(_07137_ ) );
NOR3_X1 _15135_ ( .A1(_07135_ ), .A2(_07136_ ), .A3(_07137_ ), .ZN(_07138_ ) );
OAI21_X1 _15136_ ( .A(_07040_ ), .B1(_07134_ ), .B2(_07138_ ), .ZN(_07139_ ) );
BUF_X4 _15137_ ( .A(_06943_ ), .Z(_07140_ ) );
BUF_X4 _15138_ ( .A(_07020_ ), .Z(_07141_ ) );
BUF_X4 _15139_ ( .A(_07141_ ), .Z(_07142_ ) );
NAND4_X1 _15140_ ( .A1(_07140_ ), .A2(_05116_ ), .A3(_07142_ ), .A4(_06941_ ), .ZN(_07143_ ) );
AOI21_X1 _15141_ ( .A(_06984_ ), .B1(_07139_ ), .B2(_07143_ ), .ZN(_07144_ ) );
INV_X1 _15142_ ( .A(_07144_ ), .ZN(_07145_ ) );
BUF_X2 _15143_ ( .A(_07060_ ), .Z(_07146_ ) );
AOI21_X1 _15144_ ( .A(_07045_ ), .B1(_07145_ ), .B2(_07146_ ), .ZN(_07147_ ) );
AOI21_X1 _15145_ ( .A(_03045_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07148_ ) );
NOR2_X1 _15146_ ( .A1(_06954_ ), .A2(_02812_ ), .ZN(_07149_ ) );
NOR3_X1 _15147_ ( .A1(_07011_ ), .A2(_07148_ ), .A3(_07149_ ), .ZN(_07150_ ) );
AOI21_X1 _15148_ ( .A(_02788_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07151_ ) );
NOR2_X1 _15149_ ( .A1(_07015_ ), .A2(_02764_ ), .ZN(_07152_ ) );
NOR3_X1 _15150_ ( .A1(_07151_ ), .A2(_07152_ ), .A3(_07020_ ), .ZN(_07153_ ) );
NOR2_X1 _15151_ ( .A1(_07150_ ), .A2(_07153_ ), .ZN(_07154_ ) );
NOR2_X1 _15152_ ( .A1(_07154_ ), .A2(_07040_ ), .ZN(_07155_ ) );
AOI21_X1 _15153_ ( .A(_03095_ ), .B1(_06960_ ), .B2(_06961_ ), .ZN(_07156_ ) );
INV_X1 _15154_ ( .A(_07156_ ), .ZN(_07157_ ) );
NOR2_X1 _15155_ ( .A1(_07015_ ), .A2(_03068_ ), .ZN(_07158_ ) );
INV_X1 _15156_ ( .A(_07158_ ), .ZN(_07159_ ) );
NAND3_X1 _15157_ ( .A1(_07157_ ), .A2(_07036_ ), .A3(_07159_ ), .ZN(_07160_ ) );
AOI21_X1 _15158_ ( .A(_02948_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07161_ ) );
INV_X1 _15159_ ( .A(_07161_ ), .ZN(_07162_ ) );
NOR2_X1 _15160_ ( .A1(_07015_ ), .A2(_04854_ ), .ZN(_07163_ ) );
INV_X1 _15161_ ( .A(_07163_ ), .ZN(_07164_ ) );
NAND3_X1 _15162_ ( .A1(_07162_ ), .A2(_07033_ ), .A3(_07164_ ), .ZN(_07165_ ) );
AOI21_X1 _15163_ ( .A(_07140_ ), .B1(_07160_ ), .B2(_07165_ ), .ZN(_07166_ ) );
NOR3_X1 _15164_ ( .A1(_07155_ ), .A2(_07054_ ), .A3(_07166_ ), .ZN(_07167_ ) );
AOI21_X1 _15165_ ( .A(_03020_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07168_ ) );
INV_X1 _15166_ ( .A(_07168_ ), .ZN(_07169_ ) );
NOR2_X1 _15167_ ( .A1(_07015_ ), .A2(_04781_ ), .ZN(_07170_ ) );
INV_X1 _15168_ ( .A(_07170_ ), .ZN(_07171_ ) );
NAND3_X1 _15169_ ( .A1(_07169_ ), .A2(_07011_ ), .A3(_07171_ ), .ZN(_07172_ ) );
AOI21_X1 _15170_ ( .A(_02709_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07173_ ) );
INV_X1 _15171_ ( .A(_07173_ ), .ZN(_07174_ ) );
NOR2_X1 _15172_ ( .A1(_06941_ ), .A2(_02996_ ), .ZN(_07175_ ) );
INV_X1 _15173_ ( .A(_07175_ ), .ZN(_07176_ ) );
NAND3_X1 _15174_ ( .A1(_07174_ ), .A2(_06939_ ), .A3(_07176_ ), .ZN(_07177_ ) );
AND3_X1 _15175_ ( .A1(_07172_ ), .A2(_07177_ ), .A3(_06943_ ), .ZN(_07178_ ) );
NOR2_X1 _15176_ ( .A1(_06954_ ), .A2(_04380_ ), .ZN(_07179_ ) );
OAI21_X1 _15177_ ( .A(_07141_ ), .B1(_07111_ ), .B2(_07179_ ), .ZN(_07180_ ) );
BUF_X4 _15178_ ( .A(_06958_ ), .Z(_07181_ ) );
AND3_X1 _15179_ ( .A1(_06954_ ), .A2(_02614_ ), .A3(_02633_ ), .ZN(_07182_ ) );
NOR2_X1 _15180_ ( .A1(_07015_ ), .A2(_02684_ ), .ZN(_07183_ ) );
OAI21_X1 _15181_ ( .A(_07181_ ), .B1(_07182_ ), .B2(_07183_ ), .ZN(_07184_ ) );
AOI21_X1 _15182_ ( .A(_06965_ ), .B1(_07180_ ), .B2(_07184_ ), .ZN(_07185_ ) );
OR2_X1 _15183_ ( .A1(_07178_ ), .A2(_07185_ ), .ZN(_07186_ ) );
AOI21_X1 _15184_ ( .A(_07167_ ), .B1(_07010_ ), .B2(_07186_ ), .ZN(_07187_ ) );
OAI21_X1 _15185_ ( .A(_07147_ ), .B1(_07187_ ), .B2(_07061_ ), .ZN(_07188_ ) );
NAND3_X1 _15186_ ( .A1(_07126_ ), .A2(_06996_ ), .A3(_06992_ ), .ZN(_07189_ ) );
BUF_X4 _15187_ ( .A(_07065_ ), .Z(_07190_ ) );
OAI211_X1 _15188_ ( .A(_07188_ ), .B(_07189_ ), .C1(_06872_ ), .C2(_07190_ ), .ZN(_07191_ ) );
BUF_X2 _15189_ ( .A(_07068_ ), .Z(_07192_ ) );
AOI211_X1 _15190_ ( .A(_07131_ ), .B(_07191_ ), .C1(_05314_ ), .C2(_07192_ ), .ZN(_07193_ ) );
NAND3_X1 _15191_ ( .A1(_07095_ ), .A2(_07128_ ), .A3(_07193_ ), .ZN(_07194_ ) );
AOI21_X1 _15192_ ( .A(_07093_ ), .B1(_07194_ ), .B2(_07078_ ), .ZN(_07195_ ) );
OAI21_X1 _15193_ ( .A(_07080_ ), .B1(_05616_ ), .B2(_05921_ ), .ZN(_07196_ ) );
OAI21_X1 _15194_ ( .A(_07082_ ), .B1(_07195_ ), .B2(_07196_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OR2_X1 _15195_ ( .A1(_05658_ ), .A2(_06502_ ), .ZN(_07197_ ) );
INV_X1 _15196_ ( .A(_04353_ ), .ZN(_07198_ ) );
INV_X1 _15197_ ( .A(_04378_ ), .ZN(_07199_ ) );
AOI211_X1 _15198_ ( .A(_07198_ ), .B(_07199_ ), .C1(_05409_ ), .C2(_05424_ ), .ZN(_07200_ ) );
OR3_X1 _15199_ ( .A1(_07200_ ), .A2(_04376_ ), .A3(_05429_ ), .ZN(_07201_ ) );
NAND2_X1 _15200_ ( .A1(_07201_ ), .A2(_04431_ ), .ZN(_07202_ ) );
INV_X1 _15201_ ( .A(_04408_ ), .ZN(_07203_ ) );
NAND2_X1 _15202_ ( .A1(_02635_ ), .A2(_04429_ ), .ZN(_07204_ ) );
AND3_X1 _15203_ ( .A1(_07202_ ), .A2(_07203_ ), .A3(_07204_ ), .ZN(_07205_ ) );
AOI21_X1 _15204_ ( .A(_07203_ ), .B1(_07202_ ), .B2(_07204_ ), .ZN(_07206_ ) );
BUF_X4 _15205_ ( .A(_07089_ ), .Z(_07207_ ) );
NOR3_X1 _15206_ ( .A1(_07205_ ), .A2(_07206_ ), .A3(_07207_ ), .ZN(_07208_ ) );
AND2_X1 _15207_ ( .A1(_05631_ ), .A2(_07084_ ), .ZN(_07209_ ) );
AND3_X1 _15208_ ( .A1(_06797_ ), .A2(\ID_EX_imm [19] ), .A3(_06785_ ), .ZN(_07210_ ) );
NOR3_X1 _15209_ ( .A1(_07208_ ), .A2(_07209_ ), .A3(_07210_ ), .ZN(_07211_ ) );
OAI21_X1 _15210_ ( .A(_06141_ ), .B1(_07211_ ), .B2(_06803_ ), .ZN(_07212_ ) );
AND2_X1 _15211_ ( .A1(_06929_ ), .A2(_06930_ ), .ZN(_07213_ ) );
XNOR2_X1 _15212_ ( .A(_06886_ ), .B(_06950_ ), .ZN(_07214_ ) );
AND4_X1 _15213_ ( .A1(_06935_ ), .A2(_06926_ ), .A3(_07214_ ), .A4(_06928_ ), .ZN(_07215_ ) );
OAI21_X1 _15214_ ( .A(_06958_ ), .B1(_06952_ ), .B2(_06955_ ), .ZN(_07216_ ) );
OAI21_X1 _15215_ ( .A(_06938_ ), .B1(_06970_ ), .B2(_06971_ ), .ZN(_07217_ ) );
AOI21_X1 _15216_ ( .A(_06950_ ), .B1(_07216_ ), .B2(_07217_ ), .ZN(_07218_ ) );
OAI21_X1 _15217_ ( .A(_06938_ ), .B1(_07034_ ), .B2(_07038_ ), .ZN(_07219_ ) );
OAI21_X1 _15218_ ( .A(_06958_ ), .B1(_06966_ ), .B2(_06967_ ), .ZN(_07220_ ) );
AOI21_X1 _15219_ ( .A(_05231_ ), .B1(_07219_ ), .B2(_07220_ ), .ZN(_07221_ ) );
NOR2_X1 _15220_ ( .A1(_07218_ ), .A2(_07221_ ), .ZN(_07222_ ) );
INV_X1 _15221_ ( .A(_06959_ ), .ZN(_07223_ ) );
INV_X1 _15222_ ( .A(_06962_ ), .ZN(_07224_ ) );
NAND3_X1 _15223_ ( .A1(_07223_ ), .A2(_06938_ ), .A3(_07224_ ), .ZN(_07225_ ) );
NAND3_X1 _15224_ ( .A1(_06976_ ), .A2(_06969_ ), .A3(_06977_ ), .ZN(_07226_ ) );
AOI21_X1 _15225_ ( .A(_05231_ ), .B1(_07225_ ), .B2(_07226_ ), .ZN(_07227_ ) );
AND4_X1 _15226_ ( .A1(_03243_ ), .A2(_05231_ ), .A3(_06937_ ), .A4(_06941_ ), .ZN(_07228_ ) );
OR2_X1 _15227_ ( .A1(_07227_ ), .A2(_07228_ ), .ZN(_07229_ ) );
MUX2_X1 _15228_ ( .A(_07222_ ), .B(_07229_ ), .S(_06983_ ), .Z(_07230_ ) );
AND2_X1 _15229_ ( .A1(_07230_ ), .A2(_06986_ ), .ZN(_07231_ ) );
OR3_X1 _15230_ ( .A1(_07213_ ), .A2(_07215_ ), .A3(_07231_ ), .ZN(_07232_ ) );
AND2_X1 _15231_ ( .A1(_07232_ ), .A2(_06883_ ), .ZN(_07233_ ) );
BUF_X2 _15232_ ( .A(_06987_ ), .Z(_07234_ ) );
AND3_X1 _15233_ ( .A1(_07230_ ), .A2(_07234_ ), .A3(_06992_ ), .ZN(_07235_ ) );
NOR3_X1 _15234_ ( .A1(_05322_ ), .A2(_06863_ ), .A3(_07190_ ), .ZN(_07236_ ) );
OAI22_X1 _15235_ ( .A1(_05324_ ), .A2(_05468_ ), .B1(_06865_ ), .B2(_07129_ ), .ZN(_07237_ ) );
NOR4_X1 _15236_ ( .A1(_07233_ ), .A2(_07235_ ), .A3(_07236_ ), .A4(_07237_ ), .ZN(_07238_ ) );
INV_X1 _15237_ ( .A(_06853_ ), .ZN(_07239_ ) );
NAND3_X1 _15238_ ( .A1(_07239_ ), .A2(_05289_ ), .A3(_05293_ ), .ZN(_07240_ ) );
AOI21_X1 _15239_ ( .A(_05319_ ), .B1(_07240_ ), .B2(_06861_ ), .ZN(_07241_ ) );
INV_X1 _15240_ ( .A(_07241_ ), .ZN(_07242_ ) );
NOR2_X1 _15241_ ( .A1(_06538_ ), .A2(_05317_ ), .ZN(_07243_ ) );
INV_X1 _15242_ ( .A(_07243_ ), .ZN(_07244_ ) );
NAND3_X1 _15243_ ( .A1(_07242_ ), .A2(_05324_ ), .A3(_07244_ ), .ZN(_07245_ ) );
BUF_X4 _15244_ ( .A(_06878_ ), .Z(_07246_ ) );
OAI21_X1 _15245_ ( .A(_05323_ ), .B1(_07241_ ), .B2(_07243_ ), .ZN(_07247_ ) );
NAND3_X1 _15246_ ( .A1(_07245_ ), .A2(_07246_ ), .A3(_07247_ ), .ZN(_07248_ ) );
OAI21_X1 _15247_ ( .A(_07141_ ), .B1(_07037_ ), .B2(_07038_ ), .ZN(_07249_ ) );
OAI21_X1 _15248_ ( .A(_07181_ ), .B1(_07026_ ), .B2(_07027_ ), .ZN(_07250_ ) );
NAND2_X1 _15249_ ( .A1(_07249_ ), .A2(_07250_ ), .ZN(_07251_ ) );
NOR3_X1 _15250_ ( .A1(_07181_ ), .A2(_07029_ ), .A3(_07030_ ), .ZN(_07252_ ) );
NOR3_X1 _15251_ ( .A1(_07014_ ), .A2(_07016_ ), .A3(_06939_ ), .ZN(_07253_ ) );
NOR2_X1 _15252_ ( .A1(_07252_ ), .A2(_07253_ ), .ZN(_07254_ ) );
BUF_X4 _15253_ ( .A(_07140_ ), .Z(_07255_ ) );
MUX2_X1 _15254_ ( .A(_07251_ ), .B(_07254_ ), .S(_07255_ ), .Z(_07256_ ) );
BUF_X2 _15255_ ( .A(_07042_ ), .Z(_07257_ ) );
OR2_X1 _15256_ ( .A1(_07256_ ), .A2(_07257_ ), .ZN(_07258_ ) );
NOR3_X1 _15257_ ( .A1(_07025_ ), .A2(_07018_ ), .A3(_07019_ ), .ZN(_07259_ ) );
NOR3_X1 _15258_ ( .A1(_06997_ ), .A2(_06998_ ), .A3(_07020_ ), .ZN(_07260_ ) );
NOR2_X1 _15259_ ( .A1(_07259_ ), .A2(_07260_ ), .ZN(_07261_ ) );
NAND2_X1 _15260_ ( .A1(_07261_ ), .A2(_06951_ ), .ZN(_07262_ ) );
NOR3_X1 _15261_ ( .A1(_07025_ ), .A2(_07000_ ), .A3(_07001_ ), .ZN(_07263_ ) );
NOR3_X1 _15262_ ( .A1(_07049_ ), .A2(_07050_ ), .A3(_07020_ ), .ZN(_07264_ ) );
NOR2_X1 _15263_ ( .A1(_07263_ ), .A2(_07264_ ), .ZN(_07265_ ) );
NAND2_X1 _15264_ ( .A1(_07265_ ), .A2(_06965_ ), .ZN(_07266_ ) );
NAND3_X1 _15265_ ( .A1(_07262_ ), .A2(_07266_ ), .A3(_07257_ ), .ZN(_07267_ ) );
NAND3_X1 _15266_ ( .A1(_07258_ ), .A2(_06988_ ), .A3(_07267_ ), .ZN(_07268_ ) );
OAI21_X1 _15267_ ( .A(_07025_ ), .B1(_07056_ ), .B2(_05243_ ), .ZN(_07269_ ) );
NOR2_X1 _15268_ ( .A1(_07046_ ), .A2(_07047_ ), .ZN(_07270_ ) );
OAI21_X1 _15269_ ( .A(_07269_ ), .B1(_07270_ ), .B2(_07011_ ), .ZN(_07271_ ) );
INV_X1 _15270_ ( .A(_07271_ ), .ZN(_07272_ ) );
NAND3_X1 _15271_ ( .A1(_07272_ ), .A2(_07008_ ), .A3(_07040_ ), .ZN(_07273_ ) );
AOI21_X1 _15272_ ( .A(_07045_ ), .B1(_07273_ ), .B2(_07061_ ), .ZN(_07274_ ) );
NAND2_X1 _15273_ ( .A1(_07268_ ), .A2(_07274_ ), .ZN(_07275_ ) );
NAND3_X1 _15274_ ( .A1(_07238_ ), .A2(_07248_ ), .A3(_07275_ ), .ZN(_07276_ ) );
AOI21_X1 _15275_ ( .A(_07212_ ), .B1(_07276_ ), .B2(_07078_ ), .ZN(_07277_ ) );
NAND2_X1 _15276_ ( .A1(_05636_ ), .A2(_05553_ ), .ZN(_07278_ ) );
NAND2_X1 _15277_ ( .A1(_07278_ ), .A2(_06492_ ), .ZN(_07279_ ) );
OAI21_X1 _15278_ ( .A(_07197_ ), .B1(_07277_ ), .B2(_07279_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
NAND2_X1 _15279_ ( .A1(_05683_ ), .A2(_06494_ ), .ZN(_07280_ ) );
BUF_X4 _15280_ ( .A(_06802_ ), .Z(_07281_ ) );
AOI21_X1 _15281_ ( .A(_07207_ ), .B1(_07201_ ), .B2(_04431_ ), .ZN(_07282_ ) );
OAI21_X1 _15282_ ( .A(_07282_ ), .B1(_04431_ ), .B2(_07201_ ), .ZN(_07283_ ) );
AOI22_X1 _15283_ ( .A1(_05667_ ), .A2(_07084_ ), .B1(\ID_EX_imm [18] ), .B2(_07087_ ), .ZN(_07284_ ) );
AOI21_X1 _15284_ ( .A(_07281_ ), .B1(_07283_ ), .B2(_07284_ ), .ZN(_07285_ ) );
OR2_X1 _15285_ ( .A1(_07285_ ), .A2(_05838_ ), .ZN(_07286_ ) );
AND2_X1 _15286_ ( .A1(_06926_ ), .A2(_07214_ ), .ZN(_07287_ ) );
INV_X1 _15287_ ( .A(_07287_ ), .ZN(_07288_ ) );
AND2_X1 _15288_ ( .A1(_06975_ ), .A2(_07142_ ), .ZN(_07289_ ) );
OR3_X1 _15289_ ( .A1(_07288_ ), .A2(_07289_ ), .A3(_06934_ ), .ZN(_07290_ ) );
AOI21_X1 _15290_ ( .A(_06932_ ), .B1(_07290_ ), .B2(_06948_ ), .ZN(_07291_ ) );
NOR3_X1 _15291_ ( .A1(_07102_ ), .A2(_07103_ ), .A3(_06937_ ), .ZN(_07292_ ) );
NOR3_X1 _15292_ ( .A1(_07114_ ), .A2(_06969_ ), .A3(_07115_ ), .ZN(_07293_ ) );
OAI21_X1 _15293_ ( .A(_06965_ ), .B1(_07292_ ), .B2(_07293_ ), .ZN(_07294_ ) );
NOR3_X1 _15294_ ( .A1(_07182_ ), .A2(_07025_ ), .A3(_07179_ ), .ZN(_07295_ ) );
NOR3_X1 _15295_ ( .A1(_07111_ ), .A2(_07020_ ), .A3(_07112_ ), .ZN(_07296_ ) );
OAI21_X1 _15296_ ( .A(_07004_ ), .B1(_07295_ ), .B2(_07296_ ), .ZN(_07297_ ) );
NAND2_X1 _15297_ ( .A1(_07294_ ), .A2(_07297_ ), .ZN(_07298_ ) );
AOI21_X1 _15298_ ( .A(_06958_ ), .B1(_07107_ ), .B2(_07108_ ), .ZN(_07299_ ) );
AOI21_X1 _15299_ ( .A(_06938_ ), .B1(_07119_ ), .B2(_07120_ ), .ZN(_07300_ ) );
OAI21_X1 _15300_ ( .A(_06950_ ), .B1(_07299_ ), .B2(_07300_ ), .ZN(_07301_ ) );
AND2_X1 _15301_ ( .A1(_07123_ ), .A2(_07137_ ), .ZN(_07302_ ) );
OAI21_X1 _15302_ ( .A(_07301_ ), .B1(_07302_ ), .B2(_07004_ ), .ZN(_07303_ ) );
INV_X1 _15303_ ( .A(_07303_ ), .ZN(_07304_ ) );
MUX2_X1 _15304_ ( .A(_07298_ ), .B(_07304_ ), .S(_06984_ ), .Z(_07305_ ) );
AND2_X1 _15305_ ( .A1(_07305_ ), .A2(_06988_ ), .ZN(_07306_ ) );
OAI21_X1 _15306_ ( .A(_06884_ ), .B1(_07291_ ), .B2(_07306_ ), .ZN(_07307_ ) );
NAND3_X1 _15307_ ( .A1(_07240_ ), .A2(_05319_ ), .A3(_06861_ ), .ZN(_07308_ ) );
NAND3_X1 _15308_ ( .A1(_07242_ ), .A2(_07246_ ), .A3(_07308_ ), .ZN(_07309_ ) );
AND3_X1 _15309_ ( .A1(_07305_ ), .A2(_07234_ ), .A3(_06992_ ), .ZN(_07310_ ) );
OAI211_X1 _15310_ ( .A(_05235_ ), .B(_05236_ ), .C1(_06975_ ), .C2(_06805_ ), .ZN(_07311_ ) );
NOR2_X1 _15311_ ( .A1(_07135_ ), .A2(_07136_ ), .ZN(_07312_ ) );
OAI21_X1 _15312_ ( .A(_07311_ ), .B1(_07312_ ), .B2(_07011_ ), .ZN(_07313_ ) );
NOR2_X1 _15313_ ( .A1(_07313_ ), .A2(_07255_ ), .ZN(_07314_ ) );
BUF_X2 _15314_ ( .A(_07008_ ), .Z(_07315_ ) );
AND2_X1 _15315_ ( .A1(_07314_ ), .A2(_07315_ ), .ZN(_07316_ ) );
OAI21_X1 _15316_ ( .A(_05464_ ), .B1(_07316_ ), .B2(_06996_ ), .ZN(_07317_ ) );
INV_X1 _15317_ ( .A(_07183_ ), .ZN(_07318_ ) );
OAI211_X1 _15318_ ( .A(_07318_ ), .B(_06939_ ), .C1(_02635_ ), .C2(_06975_ ), .ZN(_07319_ ) );
NAND3_X1 _15319_ ( .A1(_07174_ ), .A2(_07011_ ), .A3(_07176_ ), .ZN(_07320_ ) );
NAND3_X1 _15320_ ( .A1(_07319_ ), .A2(_07320_ ), .A3(_07024_ ), .ZN(_07321_ ) );
NAND3_X1 _15321_ ( .A1(_07162_ ), .A2(_07025_ ), .A3(_07164_ ), .ZN(_07322_ ) );
NAND3_X1 _15322_ ( .A1(_07169_ ), .A2(_07137_ ), .A3(_07171_ ), .ZN(_07323_ ) );
NAND3_X1 _15323_ ( .A1(_07322_ ), .A2(_07323_ ), .A3(_06981_ ), .ZN(_07324_ ) );
NAND2_X1 _15324_ ( .A1(_07321_ ), .A2(_07324_ ), .ZN(_07325_ ) );
NOR3_X1 _15325_ ( .A1(_06958_ ), .A2(_07156_ ), .A3(_07158_ ), .ZN(_07326_ ) );
NOR3_X1 _15326_ ( .A1(_07148_ ), .A2(_07149_ ), .A3(_06938_ ), .ZN(_07327_ ) );
NOR2_X1 _15327_ ( .A1(_07326_ ), .A2(_07327_ ), .ZN(_07328_ ) );
NAND2_X1 _15328_ ( .A1(_07328_ ), .A2(_07006_ ), .ZN(_07329_ ) );
OAI21_X1 _15329_ ( .A(_07025_ ), .B1(_07132_ ), .B2(_07133_ ), .ZN(_07330_ ) );
OAI21_X1 _15330_ ( .A(_07137_ ), .B1(_07151_ ), .B2(_07152_ ), .ZN(_07331_ ) );
NAND2_X1 _15331_ ( .A1(_07330_ ), .A2(_07331_ ), .ZN(_07332_ ) );
NAND2_X1 _15332_ ( .A1(_07332_ ), .A2(_06981_ ), .ZN(_07333_ ) );
NAND2_X1 _15333_ ( .A1(_07329_ ), .A2(_07333_ ), .ZN(_07334_ ) );
MUX2_X1 _15334_ ( .A(_07325_ ), .B(_07334_ ), .S(_07042_ ), .Z(_07335_ ) );
AOI21_X1 _15335_ ( .A(_07317_ ), .B1(_06988_ ), .B2(_07335_ ), .ZN(_07336_ ) );
AOI21_X1 _15336_ ( .A(_07129_ ), .B1(_06538_ ), .B2(_05317_ ), .ZN(_07337_ ) );
OAI22_X1 _15337_ ( .A1(_05319_ ), .A2(_05468_ ), .B1(_07244_ ), .B2(_07190_ ), .ZN(_07338_ ) );
NOR4_X1 _15338_ ( .A1(_07310_ ), .A2(_07336_ ), .A3(_07337_ ), .A4(_07338_ ), .ZN(_07339_ ) );
NAND3_X1 _15339_ ( .A1(_07307_ ), .A2(_07309_ ), .A3(_07339_ ), .ZN(_07340_ ) );
AOI21_X1 _15340_ ( .A(_07286_ ), .B1(_07340_ ), .B2(_07078_ ), .ZN(_07341_ ) );
OAI21_X1 _15341_ ( .A(_07080_ ), .B1(_05665_ ), .B2(_05921_ ), .ZN(_07342_ ) );
OAI21_X1 _15342_ ( .A(_07280_ ), .B1(_07341_ ), .B2(_07342_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
OR2_X1 _15343_ ( .A1(_05707_ ), .A2(_06502_ ), .ZN(_07343_ ) );
NOR2_X1 _15344_ ( .A1(_05425_ ), .A2(_07198_ ), .ZN(_07344_ ) );
INV_X1 _15345_ ( .A(_07344_ ), .ZN(_07345_ ) );
AND3_X1 _15346_ ( .A1(_07345_ ), .A2(_05428_ ), .A3(_07199_ ), .ZN(_07346_ ) );
AOI21_X1 _15347_ ( .A(_07199_ ), .B1(_07345_ ), .B2(_05428_ ), .ZN(_07347_ ) );
OR3_X1 _15348_ ( .A1(_07346_ ), .A2(_07347_ ), .A3(_07089_ ), .ZN(_07348_ ) );
AOI22_X1 _15349_ ( .A1(_05690_ ), .A2(_07084_ ), .B1(\ID_EX_imm [17] ), .B2(_07087_ ), .ZN(_07349_ ) );
AOI21_X1 _15350_ ( .A(_07281_ ), .B1(_07348_ ), .B2(_07349_ ), .ZN(_07350_ ) );
OR2_X1 _15351_ ( .A1(_07350_ ), .A2(_05838_ ), .ZN(_07351_ ) );
NAND2_X1 _15352_ ( .A1(_07239_ ), .A2(_05293_ ), .ZN(_07352_ ) );
INV_X1 _15353_ ( .A(_06860_ ), .ZN(_07353_ ) );
NAND2_X1 _15354_ ( .A1(_07352_ ), .A2(_07353_ ), .ZN(_07354_ ) );
AOI21_X1 _15355_ ( .A(_06879_ ), .B1(_07354_ ), .B2(_05289_ ), .ZN(_07355_ ) );
OAI21_X1 _15356_ ( .A(_07355_ ), .B1(_05289_ ), .B2(_07354_ ), .ZN(_07356_ ) );
OR3_X1 _15357_ ( .A1(_07037_ ), .A2(_06969_ ), .A3(_07026_ ), .ZN(_07357_ ) );
OR3_X1 _15358_ ( .A1(_07034_ ), .A2(_07038_ ), .A3(_06937_ ), .ZN(_07358_ ) );
AOI21_X1 _15359_ ( .A(_06943_ ), .B1(_07357_ ), .B2(_07358_ ), .ZN(_07359_ ) );
AND3_X1 _15360_ ( .A1(_06968_ ), .A2(_06972_ ), .A3(_05231_ ), .ZN(_07360_ ) );
NOR2_X1 _15361_ ( .A1(_07359_ ), .A2(_07360_ ), .ZN(_07361_ ) );
NAND2_X1 _15362_ ( .A1(_06980_ ), .A2(_06943_ ), .ZN(_07362_ ) );
NAND2_X1 _15363_ ( .A1(_06956_ ), .A2(_06963_ ), .ZN(_07363_ ) );
NAND2_X1 _15364_ ( .A1(_07363_ ), .A2(_06950_ ), .ZN(_07364_ ) );
NAND2_X1 _15365_ ( .A1(_07362_ ), .A2(_07364_ ), .ZN(_07365_ ) );
MUX2_X1 _15366_ ( .A(_07361_ ), .B(_07365_ ), .S(_06983_ ), .Z(_07366_ ) );
NOR2_X1 _15367_ ( .A1(_07366_ ), .A2(_07061_ ), .ZN(_07367_ ) );
BUF_X2 _15368_ ( .A(_06875_ ), .Z(_07368_ ) );
AOI22_X1 _15369_ ( .A1(_07367_ ), .A2(_06993_ ), .B1(_05339_ ), .B2(_07368_ ), .ZN(_07369_ ) );
AND2_X1 _15370_ ( .A1(_07356_ ), .A2(_07369_ ), .ZN(_07370_ ) );
AND3_X1 _15371_ ( .A1(_06933_ ), .A2(_06935_ ), .A3(_07214_ ), .ZN(_07371_ ) );
NAND2_X1 _15372_ ( .A1(_07371_ ), .A2(_06942_ ), .ZN(_07372_ ) );
AOI22_X1 _15373_ ( .A1(_07372_ ), .A2(_06948_ ), .B1(_07096_ ), .B2(_07097_ ), .ZN(_07373_ ) );
OAI21_X1 _15374_ ( .A(_06884_ ), .B1(_07373_ ), .B2(_07367_ ), .ZN(_07374_ ) );
AND3_X1 _15375_ ( .A1(_07057_ ), .A2(_07008_ ), .A3(_07040_ ), .ZN(_07375_ ) );
OAI21_X1 _15376_ ( .A(_05464_ ), .B1(_07375_ ), .B2(_06995_ ), .ZN(_07376_ ) );
NAND2_X1 _15377_ ( .A1(_07052_ ), .A2(_05231_ ), .ZN(_07377_ ) );
NAND2_X1 _15378_ ( .A1(_07003_ ), .A2(_06950_ ), .ZN(_07378_ ) );
NAND2_X1 _15379_ ( .A1(_07377_ ), .A2(_07378_ ), .ZN(_07379_ ) );
AOI21_X1 _15380_ ( .A(_06951_ ), .B1(_07017_ ), .B2(_07021_ ), .ZN(_07380_ ) );
AOI21_X1 _15381_ ( .A(_06944_ ), .B1(_07028_ ), .B2(_07031_ ), .ZN(_07381_ ) );
NOR2_X1 _15382_ ( .A1(_07380_ ), .A2(_07381_ ), .ZN(_07382_ ) );
MUX2_X1 _15383_ ( .A(_07379_ ), .B(_07382_ ), .S(_07054_ ), .Z(_07383_ ) );
AOI21_X1 _15384_ ( .A(_07376_ ), .B1(_07383_ ), .B2(_06987_ ), .ZN(_07384_ ) );
AOI221_X4 _15385_ ( .A(_07384_ ), .B1(_06858_ ), .B2(_05129_ ), .C1(_05289_ ), .C2(_07068_ ), .ZN(_07385_ ) );
NAND3_X1 _15386_ ( .A1(_07370_ ), .A2(_07374_ ), .A3(_07385_ ), .ZN(_07386_ ) );
AOI21_X1 _15387_ ( .A(_07351_ ), .B1(_07386_ ), .B2(_07078_ ), .ZN(_07387_ ) );
NAND2_X1 _15388_ ( .A1(_05695_ ), .A2(_05553_ ), .ZN(_07388_ ) );
NAND2_X1 _15389_ ( .A1(_07388_ ), .A2(_06563_ ), .ZN(_07389_ ) );
OAI21_X1 _15390_ ( .A(_07343_ ), .B1(_07387_ ), .B2(_07389_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
OR2_X1 _15391_ ( .A1(_05725_ ), .A2(_06502_ ), .ZN(_07390_ ) );
INV_X1 _15392_ ( .A(_05425_ ), .ZN(_07391_ ) );
AOI21_X1 _15393_ ( .A(_07089_ ), .B1(_07391_ ), .B2(_04353_ ), .ZN(_07392_ ) );
OAI21_X1 _15394_ ( .A(_07392_ ), .B1(_04353_ ), .B2(_07391_ ), .ZN(_07393_ ) );
AOI22_X1 _15395_ ( .A1(_05727_ ), .A2(_07084_ ), .B1(\ID_EX_imm [16] ), .B2(_07087_ ), .ZN(_07394_ ) );
AOI21_X1 _15396_ ( .A(_07281_ ), .B1(_07393_ ), .B2(_07394_ ), .ZN(_07395_ ) );
OR2_X1 _15397_ ( .A1(_07395_ ), .A2(_05838_ ), .ZN(_07396_ ) );
INV_X1 _15398_ ( .A(_06928_ ), .ZN(_07397_ ) );
INV_X1 _15399_ ( .A(_06926_ ), .ZN(_07398_ ) );
INV_X1 _15400_ ( .A(_06888_ ), .ZN(_07399_ ) );
AOI211_X1 _15401_ ( .A(_07397_ ), .B(_07398_ ), .C1(_07234_ ), .C2(_07399_ ), .ZN(_07400_ ) );
OR3_X1 _15402_ ( .A1(_07182_ ), .A2(_06938_ ), .A3(_07179_ ), .ZN(_07401_ ) );
NAND3_X1 _15403_ ( .A1(_07174_ ), .A2(_07137_ ), .A3(_07318_ ), .ZN(_07402_ ) );
AOI21_X1 _15404_ ( .A(_06943_ ), .B1(_07401_ ), .B2(_07402_ ), .ZN(_07403_ ) );
AND3_X1 _15405_ ( .A1(_07113_ ), .A2(_07116_ ), .A3(_05231_ ), .ZN(_07404_ ) );
NOR3_X1 _15406_ ( .A1(_07403_ ), .A2(_07404_ ), .A3(_06983_ ), .ZN(_07405_ ) );
OAI21_X1 _15407_ ( .A(_06951_ ), .B1(_07105_ ), .B2(_07109_ ), .ZN(_07406_ ) );
OAI21_X1 _15408_ ( .A(_07406_ ), .B1(_07124_ ), .B2(_07005_ ), .ZN(_07407_ ) );
AOI21_X1 _15409_ ( .A(_07405_ ), .B1(_07407_ ), .B2(_07042_ ), .ZN(_07408_ ) );
AND2_X1 _15410_ ( .A1(_07408_ ), .A2(_06996_ ), .ZN(_07409_ ) );
OAI21_X1 _15411_ ( .A(_06883_ ), .B1(_07400_ ), .B2(_07409_ ), .ZN(_07410_ ) );
OAI21_X1 _15412_ ( .A(_06965_ ), .B1(_07134_ ), .B2(_07138_ ), .ZN(_07411_ ) );
OAI21_X1 _15413_ ( .A(_06951_ ), .B1(_07150_ ), .B2(_07153_ ), .ZN(_07412_ ) );
NAND2_X1 _15414_ ( .A1(_07411_ ), .A2(_07412_ ), .ZN(_07413_ ) );
BUF_X2 _15415_ ( .A(_06983_ ), .Z(_07414_ ) );
BUF_X2 _15416_ ( .A(_07414_ ), .Z(_07415_ ) );
NAND2_X1 _15417_ ( .A1(_07413_ ), .A2(_07415_ ), .ZN(_07416_ ) );
NAND3_X1 _15418_ ( .A1(_07172_ ), .A2(_07177_ ), .A3(_07024_ ), .ZN(_07417_ ) );
NAND3_X1 _15419_ ( .A1(_07160_ ), .A2(_07165_ ), .A3(_06981_ ), .ZN(_07418_ ) );
NAND3_X1 _15420_ ( .A1(_07417_ ), .A2(_07418_ ), .A3(_07055_ ), .ZN(_07419_ ) );
AOI21_X1 _15421_ ( .A(_07061_ ), .B1(_07416_ ), .B2(_07419_ ), .ZN(_07420_ ) );
AND4_X1 _15422_ ( .A1(_05116_ ), .A2(_06887_ ), .A3(_07146_ ), .A4(_07055_ ), .ZN(_07421_ ) );
OAI21_X1 _15423_ ( .A(_05464_ ), .B1(_07420_ ), .B2(_07421_ ), .ZN(_07422_ ) );
NAND3_X1 _15424_ ( .A1(_07408_ ), .A2(_06988_ ), .A3(_06993_ ), .ZN(_07423_ ) );
AND3_X1 _15425_ ( .A1(_07410_ ), .A2(_07422_ ), .A3(_07423_ ), .ZN(_07424_ ) );
AOI21_X1 _15426_ ( .A(_06880_ ), .B1(_07239_ ), .B2(_05293_ ), .ZN(_07425_ ) );
OAI21_X1 _15427_ ( .A(_07425_ ), .B1(_05293_ ), .B2(_07239_ ), .ZN(_07426_ ) );
AND2_X1 _15428_ ( .A1(_05293_ ), .A2(_07192_ ), .ZN(_07427_ ) );
NOR3_X1 _15429_ ( .A1(_05292_ ), .A2(_06859_ ), .A3(_07190_ ), .ZN(_07428_ ) );
AOI21_X1 _15430_ ( .A(_07130_ ), .B1(_05292_ ), .B2(_06859_ ), .ZN(_07429_ ) );
NOR3_X1 _15431_ ( .A1(_07427_ ), .A2(_07428_ ), .A3(_07429_ ), .ZN(_07430_ ) );
NAND3_X1 _15432_ ( .A1(_07424_ ), .A2(_07426_ ), .A3(_07430_ ), .ZN(_07431_ ) );
AOI21_X1 _15433_ ( .A(_07396_ ), .B1(_07431_ ), .B2(_07078_ ), .ZN(_07432_ ) );
NAND2_X1 _15434_ ( .A1(_05729_ ), .A2(_05553_ ), .ZN(_07433_ ) );
NAND2_X1 _15435_ ( .A1(_07433_ ), .A2(_06563_ ), .ZN(_07434_ ) );
OAI21_X1 _15436_ ( .A(_07390_ ), .B1(_07432_ ), .B2(_07434_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OR2_X1 _15437_ ( .A1(_05752_ ), .A2(_06502_ ), .ZN(_07435_ ) );
INV_X1 _15438_ ( .A(_04806_ ), .ZN(_07436_ ) );
INV_X1 _15439_ ( .A(_04828_ ), .ZN(_07437_ ) );
INV_X1 _15440_ ( .A(_05408_ ), .ZN(_07438_ ) );
NAND2_X1 _15441_ ( .A1(_07438_ ), .A2(_04928_ ), .ZN(_07439_ ) );
AOI211_X1 _15442_ ( .A(_07436_ ), .B(_07437_ ), .C1(_07439_ ), .C2(_05418_ ), .ZN(_07440_ ) );
OAI21_X1 _15443_ ( .A(_04753_ ), .B1(_07440_ ), .B2(_05423_ ), .ZN(_07441_ ) );
NAND2_X1 _15444_ ( .A1(_03020_ ), .A2(_04752_ ), .ZN(_07442_ ) );
AND2_X1 _15445_ ( .A1(_07441_ ), .A2(_07442_ ), .ZN(_07443_ ) );
XNOR2_X1 _15446_ ( .A(_07443_ ), .B(_04779_ ), .ZN(_07444_ ) );
BUF_X4 _15447_ ( .A(_06795_ ), .Z(_07445_ ) );
NAND2_X1 _15448_ ( .A1(_07444_ ), .A2(_07445_ ), .ZN(_07446_ ) );
AOI22_X1 _15449_ ( .A1(_05739_ ), .A2(_07083_ ), .B1(\ID_EX_imm [15] ), .B2(_07087_ ), .ZN(_07447_ ) );
AOI21_X1 _15450_ ( .A(_07281_ ), .B1(_07446_ ), .B2(_07447_ ), .ZN(_07448_ ) );
OR2_X1 _15451_ ( .A1(_07448_ ), .A2(_05838_ ), .ZN(_07449_ ) );
NAND2_X1 _15452_ ( .A1(_06826_ ), .A2(_06831_ ), .ZN(_07450_ ) );
AND2_X1 _15453_ ( .A1(_06837_ ), .A2(_06840_ ), .ZN(_07451_ ) );
AND2_X1 _15454_ ( .A1(_07450_ ), .A2(_07451_ ), .ZN(_07452_ ) );
INV_X1 _15455_ ( .A(_07452_ ), .ZN(_07453_ ) );
NAND2_X1 _15456_ ( .A1(_07453_ ), .A2(_06827_ ), .ZN(_07454_ ) );
AOI21_X1 _15457_ ( .A(_05167_ ), .B1(_07454_ ), .B2(_06845_ ), .ZN(_07455_ ) );
INV_X1 _15458_ ( .A(_07455_ ), .ZN(_07456_ ) );
NAND3_X1 _15459_ ( .A1(_07456_ ), .A2(_05172_ ), .A3(_06849_ ), .ZN(_07457_ ) );
OAI21_X1 _15460_ ( .A(_05171_ ), .B1(_07455_ ), .B2(_06848_ ), .ZN(_07458_ ) );
NAND3_X1 _15461_ ( .A1(_07457_ ), .A2(_07246_ ), .A3(_07458_ ), .ZN(_07459_ ) );
NAND4_X1 _15462_ ( .A1(_06933_ ), .A2(_06884_ ), .A3(_06930_ ), .A4(_06928_ ), .ZN(_07460_ ) );
NAND2_X1 _15463_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_07461_ ) );
NOR3_X1 _15464_ ( .A1(_07037_ ), .A2(_07026_ ), .A3(_06939_ ), .ZN(_07462_ ) );
NOR3_X1 _15465_ ( .A1(_07181_ ), .A2(_07029_ ), .A3(_07027_ ), .ZN(_07463_ ) );
OAI21_X1 _15466_ ( .A(_07005_ ), .B1(_07462_ ), .B2(_07463_ ), .ZN(_07464_ ) );
NAND3_X1 _15467_ ( .A1(_07219_ ), .A2(_07220_ ), .A3(_06944_ ), .ZN(_07465_ ) );
AND2_X1 _15468_ ( .A1(_07464_ ), .A2(_07465_ ), .ZN(_07466_ ) );
OR2_X1 _15469_ ( .A1(_07466_ ), .A2(_07414_ ), .ZN(_07467_ ) );
AND3_X1 _15470_ ( .A1(_07225_ ), .A2(_06944_ ), .A3(_07226_ ), .ZN(_07468_ ) );
AOI21_X1 _15471_ ( .A(_06944_ ), .B1(_07216_ ), .B2(_07217_ ), .ZN(_07469_ ) );
OR3_X1 _15472_ ( .A1(_07468_ ), .A2(_07009_ ), .A3(_07469_ ), .ZN(_07470_ ) );
AND3_X1 _15473_ ( .A1(_07467_ ), .A2(_06987_ ), .A3(_07470_ ), .ZN(_07471_ ) );
NAND3_X1 _15474_ ( .A1(_06887_ ), .A2(_03243_ ), .A3(_05233_ ), .ZN(_07472_ ) );
AOI211_X1 _15475_ ( .A(_07461_ ), .B(_07471_ ), .C1(_07061_ ), .C2(_07472_ ), .ZN(_07473_ ) );
MUX2_X1 _15476_ ( .A(_07271_ ), .B(_07265_ ), .S(_07004_ ), .Z(_07474_ ) );
NAND2_X1 _15477_ ( .A1(_07474_ ), .A2(_07414_ ), .ZN(_07475_ ) );
OAI21_X1 _15478_ ( .A(_07140_ ), .B1(_07259_ ), .B2(_07260_ ), .ZN(_07476_ ) );
OAI21_X1 _15479_ ( .A(_07005_ ), .B1(_07252_ ), .B2(_07253_ ), .ZN(_07477_ ) );
NAND3_X1 _15480_ ( .A1(_07476_ ), .A2(_07477_ ), .A3(_07009_ ), .ZN(_07478_ ) );
AND2_X1 _15481_ ( .A1(_05217_ ), .A2(_05464_ ), .ZN(_07479_ ) );
BUF_X2 _15482_ ( .A(_07479_ ), .Z(_07480_ ) );
AND3_X1 _15483_ ( .A1(_07475_ ), .A2(_07478_ ), .A3(_07480_ ), .ZN(_07481_ ) );
NOR3_X1 _15484_ ( .A1(_06850_ ), .A2(_06842_ ), .A3(_05468_ ), .ZN(_07482_ ) );
NAND2_X1 _15485_ ( .A1(_06842_ ), .A2(_06875_ ), .ZN(_07483_ ) );
OAI21_X1 _15486_ ( .A(_07483_ ), .B1(_06850_ ), .B2(_07129_ ), .ZN(_07484_ ) );
NOR4_X1 _15487_ ( .A1(_07473_ ), .A2(_07481_ ), .A3(_07482_ ), .A4(_07484_ ), .ZN(_07485_ ) );
NAND3_X1 _15488_ ( .A1(_07459_ ), .A2(_07460_ ), .A3(_07485_ ), .ZN(_07486_ ) );
AOI21_X1 _15489_ ( .A(_07449_ ), .B1(_07486_ ), .B2(_07078_ ), .ZN(_07487_ ) );
NAND2_X1 _15490_ ( .A1(_05742_ ), .A2(_05553_ ), .ZN(_07488_ ) );
NAND2_X1 _15491_ ( .A1(_07488_ ), .A2(_06563_ ), .ZN(_07489_ ) );
OAI21_X1 _15492_ ( .A(_07435_ ), .B1(_07487_ ), .B2(_07489_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
OR2_X1 _15493_ ( .A1(_05767_ ), .A2(_06502_ ), .ZN(_07490_ ) );
OR3_X1 _15494_ ( .A1(_07440_ ), .A2(_04753_ ), .A3(_05423_ ), .ZN(_07491_ ) );
NAND3_X1 _15495_ ( .A1(_07491_ ), .A2(_07445_ ), .A3(_07441_ ), .ZN(_07492_ ) );
AOI22_X1 _15496_ ( .A1(_05772_ ), .A2(_07083_ ), .B1(\ID_EX_imm [14] ), .B2(_07086_ ), .ZN(_07493_ ) );
AOI21_X1 _15497_ ( .A(_07281_ ), .B1(_07492_ ), .B2(_07493_ ), .ZN(_07494_ ) );
OR2_X1 _15498_ ( .A1(_07494_ ), .A2(_05552_ ), .ZN(_07495_ ) );
NAND3_X1 _15499_ ( .A1(_07454_ ), .A2(_05167_ ), .A3(_06845_ ), .ZN(_07496_ ) );
NAND3_X1 _15500_ ( .A1(_07456_ ), .A2(_07246_ ), .A3(_07496_ ), .ZN(_07497_ ) );
AND2_X1 _15501_ ( .A1(_06928_ ), .A2(_06930_ ), .ZN(_07498_ ) );
INV_X1 _15502_ ( .A(_07498_ ), .ZN(_07499_ ) );
NOR2_X1 _15503_ ( .A1(_06936_ ), .A2(_07499_ ), .ZN(_07500_ ) );
BUF_X2 _15504_ ( .A(_07498_ ), .Z(_07501_ ) );
NAND3_X1 _15505_ ( .A1(_06975_ ), .A2(_07033_ ), .A3(_06951_ ), .ZN(_07502_ ) );
NAND4_X1 _15506_ ( .A1(_06916_ ), .A2(_06925_ ), .A3(_07501_ ), .A4(_07502_ ), .ZN(_07503_ ) );
OR3_X1 _15507_ ( .A1(_07292_ ), .A2(_07293_ ), .A3(_05231_ ), .ZN(_07504_ ) );
OAI21_X1 _15508_ ( .A(_06943_ ), .B1(_07299_ ), .B2(_07300_ ), .ZN(_07505_ ) );
NAND3_X1 _15509_ ( .A1(_07504_ ), .A2(_07042_ ), .A3(_07505_ ), .ZN(_07506_ ) );
OAI21_X1 _15510_ ( .A(_06981_ ), .B1(_07295_ ), .B2(_07296_ ), .ZN(_07507_ ) );
OAI21_X1 _15511_ ( .A(_07033_ ), .B1(_07168_ ), .B2(_07175_ ), .ZN(_07508_ ) );
OAI21_X1 _15512_ ( .A(_07036_ ), .B1(_07173_ ), .B2(_07183_ ), .ZN(_07509_ ) );
NAND3_X1 _15513_ ( .A1(_07508_ ), .A2(_07509_ ), .A3(_07024_ ), .ZN(_07510_ ) );
AND2_X1 _15514_ ( .A1(_07507_ ), .A2(_07510_ ), .ZN(_07511_ ) );
OAI211_X1 _15515_ ( .A(_07506_ ), .B(_06996_ ), .C1(_07511_ ), .C2(_07415_ ), .ZN(_07512_ ) );
AND3_X1 _15516_ ( .A1(_07123_ ), .A2(_06950_ ), .A3(_07137_ ), .ZN(_07513_ ) );
INV_X1 _15517_ ( .A(_07513_ ), .ZN(_07514_ ) );
OAI21_X1 _15518_ ( .A(_07061_ ), .B1(_07514_ ), .B2(_07415_ ), .ZN(_07515_ ) );
NAND2_X1 _15519_ ( .A1(_07512_ ), .A2(_07515_ ), .ZN(_07516_ ) );
NAND2_X1 _15520_ ( .A1(_07503_ ), .A2(_07516_ ), .ZN(_07517_ ) );
OAI21_X1 _15521_ ( .A(_06884_ ), .B1(_07500_ ), .B2(_07517_ ), .ZN(_07518_ ) );
NAND3_X1 _15522_ ( .A1(_07512_ ), .A2(_06993_ ), .A3(_07515_ ), .ZN(_07519_ ) );
NOR2_X1 _15523_ ( .A1(_07328_ ), .A2(_07004_ ), .ZN(_07520_ ) );
AOI21_X1 _15524_ ( .A(_06943_ ), .B1(_07322_ ), .B2(_07323_ ), .ZN(_07521_ ) );
OR2_X1 _15525_ ( .A1(_07520_ ), .A2(_07521_ ), .ZN(_07522_ ) );
AND2_X1 _15526_ ( .A1(_07522_ ), .A2(_07009_ ), .ZN(_07523_ ) );
MUX2_X1 _15527_ ( .A(_07332_ ), .B(_07313_ ), .S(_06965_ ), .Z(_07524_ ) );
NOR2_X1 _15528_ ( .A1(_07524_ ), .A2(_07009_ ), .ZN(_07525_ ) );
OAI21_X1 _15529_ ( .A(_07480_ ), .B1(_07523_ ), .B2(_07525_ ), .ZN(_07526_ ) );
NAND2_X1 _15530_ ( .A1(_06848_ ), .A2(_07368_ ), .ZN(_07527_ ) );
AOI21_X1 _15531_ ( .A(_05130_ ), .B1(_05165_ ), .B2(_06847_ ), .ZN(_07528_ ) );
AOI21_X1 _15532_ ( .A(_07528_ ), .B1(_05166_ ), .B2(_07068_ ), .ZN(_07529_ ) );
AND4_X1 _15533_ ( .A1(_07519_ ), .A2(_07526_ ), .A3(_07527_ ), .A4(_07529_ ), .ZN(_07530_ ) );
NAND3_X1 _15534_ ( .A1(_07497_ ), .A2(_07518_ ), .A3(_07530_ ), .ZN(_07531_ ) );
AOI21_X1 _15535_ ( .A(_07495_ ), .B1(_07531_ ), .B2(_07078_ ), .ZN(_07532_ ) );
OAI21_X1 _15536_ ( .A(_07080_ ), .B1(_05770_ ), .B2(_05921_ ), .ZN(_07533_ ) );
OAI21_X1 _15537_ ( .A(_07490_ ), .B1(_07532_ ), .B2(_07533_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
NAND2_X1 _15538_ ( .A1(_05786_ ), .A2(_06494_ ), .ZN(_07534_ ) );
AND2_X1 _15539_ ( .A1(_07439_ ), .A2(_05418_ ), .ZN(_07535_ ) );
OR2_X1 _15540_ ( .A1(_07535_ ), .A2(_07437_ ), .ZN(_07536_ ) );
INV_X1 _15541_ ( .A(_05420_ ), .ZN(_07537_ ) );
AND3_X1 _15542_ ( .A1(_07536_ ), .A2(_07436_ ), .A3(_07537_ ), .ZN(_07538_ ) );
AOI21_X1 _15543_ ( .A(_07436_ ), .B1(_07536_ ), .B2(_07537_ ), .ZN(_07539_ ) );
OR3_X1 _15544_ ( .A1(_07538_ ), .A2(_07539_ ), .A3(_07089_ ), .ZN(_07540_ ) );
AOI22_X1 _15545_ ( .A1(_05790_ ), .A2(_07083_ ), .B1(\ID_EX_imm [13] ), .B2(_07086_ ), .ZN(_07541_ ) );
AOI21_X1 _15546_ ( .A(_07281_ ), .B1(_07540_ ), .B2(_07541_ ), .ZN(_07542_ ) );
OR2_X1 _15547_ ( .A1(_07542_ ), .A2(_05552_ ), .ZN(_07543_ ) );
INV_X1 _15548_ ( .A(_06882_ ), .ZN(_07544_ ) );
AND2_X1 _15549_ ( .A1(_06934_ ), .A2(_06945_ ), .ZN(_07545_ ) );
OR4_X1 _15550_ ( .A1(_06948_ ), .A2(_07398_ ), .A3(_07397_ ), .A4(_07545_ ), .ZN(_07546_ ) );
NAND3_X1 _15551_ ( .A1(_07357_ ), .A2(_07358_ ), .A3(_07140_ ), .ZN(_07547_ ) );
OR3_X1 _15552_ ( .A1(_07025_ ), .A2(_07014_ ), .A3(_07030_ ), .ZN(_07548_ ) );
OR3_X1 _15553_ ( .A1(_07029_ ), .A2(_07027_ ), .A3(_07020_ ), .ZN(_07549_ ) );
NAND3_X1 _15554_ ( .A1(_07548_ ), .A2(_07040_ ), .A3(_07549_ ), .ZN(_07550_ ) );
AOI21_X1 _15555_ ( .A(_07414_ ), .B1(_07547_ ), .B2(_07550_ ), .ZN(_07551_ ) );
NOR2_X1 _15556_ ( .A1(_06974_ ), .A2(_07315_ ), .ZN(_07552_ ) );
AOI211_X1 _15557_ ( .A(_07551_ ), .B(_07552_ ), .C1(_05215_ ), .C2(_05216_ ), .ZN(_07553_ ) );
NOR4_X1 _15558_ ( .A1(_06980_ ), .A2(_06995_ ), .A3(_07042_ ), .A4(_07255_ ), .ZN(_07554_ ) );
NOR2_X1 _15559_ ( .A1(_07553_ ), .A2(_07554_ ), .ZN(_07555_ ) );
AOI21_X1 _15560_ ( .A(_07544_ ), .B1(_07546_ ), .B2(_07555_ ), .ZN(_07556_ ) );
INV_X1 _15561_ ( .A(_06991_ ), .ZN(_07557_ ) );
NOR2_X1 _15562_ ( .A1(_07555_ ), .A2(_07557_ ), .ZN(_07558_ ) );
INV_X1 _15563_ ( .A(_07479_ ), .ZN(_07559_ ) );
OAI21_X1 _15564_ ( .A(_07010_ ), .B1(_07007_ ), .B2(_07022_ ), .ZN(_07560_ ) );
NAND3_X1 _15565_ ( .A1(_07053_ ), .A2(_07042_ ), .A3(_07058_ ), .ZN(_07561_ ) );
AOI21_X1 _15566_ ( .A(_07559_ ), .B1(_07560_ ), .B2(_07561_ ), .ZN(_07562_ ) );
NAND2_X1 _15567_ ( .A1(_05182_ ), .A2(_07068_ ), .ZN(_07563_ ) );
NAND2_X1 _15568_ ( .A1(_06843_ ), .A2(_07368_ ), .ZN(_07564_ ) );
NAND2_X1 _15569_ ( .A1(_07563_ ), .A2(_07564_ ), .ZN(_07565_ ) );
NOR4_X1 _15570_ ( .A1(_07556_ ), .A2(_07558_ ), .A3(_07562_ ), .A4(_07565_ ), .ZN(_07566_ ) );
AOI21_X1 _15571_ ( .A(_05177_ ), .B1(_07450_ ), .B2(_07451_ ), .ZN(_07567_ ) );
OR2_X1 _15572_ ( .A1(_07567_ ), .A2(_06844_ ), .ZN(_07568_ ) );
AOI21_X1 _15573_ ( .A(_06880_ ), .B1(_07568_ ), .B2(_05182_ ), .ZN(_07569_ ) );
OAI21_X1 _15574_ ( .A(_07569_ ), .B1(_05182_ ), .B2(_07568_ ), .ZN(_07570_ ) );
AND2_X1 _15575_ ( .A1(_05181_ ), .A2(_06574_ ), .ZN(_07571_ ) );
OR2_X1 _15576_ ( .A1(_07571_ ), .A2(_07130_ ), .ZN(_07572_ ) );
NAND3_X1 _15577_ ( .A1(_07566_ ), .A2(_07570_ ), .A3(_07572_ ), .ZN(_07573_ ) );
AOI21_X1 _15578_ ( .A(_07543_ ), .B1(_07573_ ), .B2(_07078_ ), .ZN(_07574_ ) );
OAI21_X1 _15579_ ( .A(_07080_ ), .B1(_05787_ ), .B2(_05921_ ), .ZN(_07575_ ) );
OAI21_X1 _15580_ ( .A(_07534_ ), .B1(_07574_ ), .B2(_07575_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
OR2_X1 _15581_ ( .A1(_05810_ ), .A2(_06491_ ), .ZN(_07576_ ) );
NAND3_X1 _15582_ ( .A1(_07439_ ), .A2(_07437_ ), .A3(_05418_ ), .ZN(_07577_ ) );
NAND3_X1 _15583_ ( .A1(_07536_ ), .A2(_07445_ ), .A3(_07577_ ), .ZN(_07578_ ) );
AOI22_X1 _15584_ ( .A1(_05796_ ), .A2(_07083_ ), .B1(\ID_EX_imm [12] ), .B2(_07086_ ), .ZN(_07579_ ) );
AOI21_X1 _15585_ ( .A(_07281_ ), .B1(_07578_ ), .B2(_07579_ ), .ZN(_07580_ ) );
OR2_X1 _15586_ ( .A1(_07580_ ), .A2(_05552_ ), .ZN(_07581_ ) );
NAND3_X1 _15587_ ( .A1(_07401_ ), .A2(_06965_ ), .A3(_07402_ ), .ZN(_07582_ ) );
OAI21_X1 _15588_ ( .A(_07137_ ), .B1(_07161_ ), .B2(_07170_ ), .ZN(_07583_ ) );
OAI21_X1 _15589_ ( .A(_06958_ ), .B1(_07168_ ), .B2(_07175_ ), .ZN(_07584_ ) );
AND2_X1 _15590_ ( .A1(_07583_ ), .A2(_07584_ ), .ZN(_07585_ ) );
OAI21_X1 _15591_ ( .A(_07582_ ), .B1(_06944_ ), .B2(_07585_ ), .ZN(_07586_ ) );
NAND2_X1 _15592_ ( .A1(_07586_ ), .A2(_07054_ ), .ZN(_07587_ ) );
OAI211_X1 _15593_ ( .A(_07587_ ), .B(_06995_ ), .C1(_07118_ ), .C2(_07315_ ), .ZN(_07588_ ) );
NAND4_X1 _15594_ ( .A1(_07124_ ), .A2(_07060_ ), .A3(_07315_ ), .A4(_07006_ ), .ZN(_07589_ ) );
AND2_X1 _15595_ ( .A1(_07588_ ), .A2(_07589_ ), .ZN(_07590_ ) );
OAI21_X1 _15596_ ( .A(_07590_ ), .B1(_06936_ ), .B2(_07499_ ), .ZN(_07591_ ) );
AND4_X1 _15597_ ( .A1(_06934_ ), .A2(_06933_ ), .A3(_07099_ ), .A4(_07501_ ), .ZN(_07592_ ) );
OAI21_X1 _15598_ ( .A(_06884_ ), .B1(_07591_ ), .B2(_07592_ ), .ZN(_07593_ ) );
NOR2_X1 _15599_ ( .A1(_07567_ ), .A2(_06880_ ), .ZN(_07594_ ) );
OAI21_X1 _15600_ ( .A(_07594_ ), .B1(_05176_ ), .B2(_07453_ ), .ZN(_07595_ ) );
OR2_X1 _15601_ ( .A1(_07590_ ), .A2(_07557_ ), .ZN(_07596_ ) );
OAI21_X1 _15602_ ( .A(_07010_ ), .B1(_07155_ ), .B2(_07166_ ), .ZN(_07597_ ) );
AND2_X1 _15603_ ( .A1(_07139_ ), .A2(_07143_ ), .ZN(_07598_ ) );
OAI21_X1 _15604_ ( .A(_07597_ ), .B1(_07598_ ), .B2(_07055_ ), .ZN(_07599_ ) );
NAND2_X1 _15605_ ( .A1(_07599_ ), .A2(_07480_ ), .ZN(_07600_ ) );
NAND3_X1 _15606_ ( .A1(_05271_ ), .A2(_02948_ ), .A3(_07368_ ), .ZN(_07601_ ) );
AOI21_X1 _15607_ ( .A(_05130_ ), .B1(_05175_ ), .B2(_05270_ ), .ZN(_07602_ ) );
AOI21_X1 _15608_ ( .A(_07602_ ), .B1(_05176_ ), .B2(_07068_ ), .ZN(_07603_ ) );
AND4_X1 _15609_ ( .A1(_07596_ ), .A2(_07600_ ), .A3(_07601_ ), .A4(_07603_ ), .ZN(_07604_ ) );
NAND3_X1 _15610_ ( .A1(_07593_ ), .A2(_07595_ ), .A3(_07604_ ), .ZN(_07605_ ) );
AOI21_X1 _15611_ ( .A(_07581_ ), .B1(_07605_ ), .B2(_07078_ ), .ZN(_07606_ ) );
OAI21_X1 _15612_ ( .A(_07080_ ), .B1(_05798_ ), .B2(_05921_ ), .ZN(_07607_ ) );
OAI21_X1 _15613_ ( .A(_07576_ ), .B1(_07606_ ), .B2(_07607_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
OR2_X1 _15614_ ( .A1(_05549_ ), .A2(_06491_ ), .ZN(_07608_ ) );
OR2_X1 _15615_ ( .A1(_04179_ ), .A2(_05479_ ), .ZN(_07609_ ) );
AOI22_X1 _15616_ ( .A1(_04290_ ), .A2(_07084_ ), .B1(\ID_EX_imm [30] ), .B2(_07087_ ), .ZN(_07610_ ) );
NAND2_X1 _15617_ ( .A1(_07391_ ), .A2(_04531_ ), .ZN(_07611_ ) );
NAND2_X1 _15618_ ( .A1(_07611_ ), .A2(_05442_ ), .ZN(_07612_ ) );
NAND2_X1 _15619_ ( .A1(_07612_ ), .A2(_04678_ ), .ZN(_07613_ ) );
NAND2_X1 _15620_ ( .A1(_07613_ ), .A2(_05459_ ), .ZN(_07614_ ) );
AOI21_X1 _15621_ ( .A(_05456_ ), .B1(_07614_ ), .B2(_04724_ ), .ZN(_07615_ ) );
INV_X1 _15622_ ( .A(_04560_ ), .ZN(_07616_ ) );
NOR4_X1 _15623_ ( .A1(_07615_ ), .A2(_04583_ ), .A3(_04582_ ), .A4(_07616_ ), .ZN(_07617_ ) );
OR2_X1 _15624_ ( .A1(_07617_ ), .A2(_05447_ ), .ZN(_07618_ ) );
AOI21_X1 _15625_ ( .A(_07207_ ), .B1(_07618_ ), .B2(_04607_ ), .ZN(_07619_ ) );
OAI21_X1 _15626_ ( .A(_07619_ ), .B1(_04607_ ), .B2(_07618_ ), .ZN(_07620_ ) );
AOI21_X1 _15627_ ( .A(_06803_ ), .B1(_07610_ ), .B2(_07620_ ), .ZN(_07621_ ) );
OR2_X1 _15628_ ( .A1(_07621_ ), .A2(_05838_ ), .ZN(_07622_ ) );
AND4_X1 _15629_ ( .A1(_05358_ ), .A2(_05354_ ), .A3(_05366_ ), .A4(_05371_ ), .ZN(_07623_ ) );
NOR3_X1 _15630_ ( .A1(_05298_ ), .A2(_05308_ ), .A3(_05309_ ), .ZN(_07624_ ) );
NAND3_X1 _15631_ ( .A1(_07624_ ), .A2(_05302_ ), .A3(_05314_ ), .ZN(_07625_ ) );
AOI211_X1 _15632_ ( .A(_06856_ ), .B(_07625_ ), .C1(_06832_ ), .C2(_06852_ ), .ZN(_07626_ ) );
OR2_X1 _15633_ ( .A1(_06867_ ), .A2(_07625_ ), .ZN(_07627_ ) );
INV_X1 _15634_ ( .A(_05308_ ), .ZN(_07628_ ) );
NAND2_X1 _15635_ ( .A1(_05302_ ), .A2(_06871_ ), .ZN(_07629_ ) );
OAI21_X1 _15636_ ( .A(_07629_ ), .B1(_07064_ ), .B2(_05301_ ), .ZN(_07630_ ) );
NAND3_X1 _15637_ ( .A1(_07630_ ), .A2(_05328_ ), .A3(_05297_ ), .ZN(_07631_ ) );
INV_X1 _15638_ ( .A(_05309_ ), .ZN(_07632_ ) );
INV_X1 _15639_ ( .A(_02535_ ), .ZN(_07633_ ) );
NOR2_X1 _15640_ ( .A1(_07633_ ), .A2(_05296_ ), .ZN(_07634_ ) );
NAND3_X1 _15641_ ( .A1(_07628_ ), .A2(_07632_ ), .A3(_07634_ ), .ZN(_07635_ ) );
NAND4_X1 _15642_ ( .A1(_07627_ ), .A2(_07628_ ), .A3(_07631_ ), .A4(_07635_ ), .ZN(_07636_ ) );
OAI21_X1 _15643_ ( .A(_07623_ ), .B1(_07626_ ), .B2(_07636_ ), .ZN(_07637_ ) );
NOR2_X1 _15644_ ( .A1(_05455_ ), .A2(_05357_ ), .ZN(_07638_ ) );
INV_X1 _15645_ ( .A(_05370_ ), .ZN(_07639_ ) );
AND2_X1 _15646_ ( .A1(_07639_ ), .A2(_03184_ ), .ZN(_07640_ ) );
AOI21_X1 _15647_ ( .A(_07640_ ), .B1(_05364_ ), .B2(_05371_ ), .ZN(_07641_ ) );
NOR4_X1 _15648_ ( .A1(_07641_ ), .A2(_05378_ ), .A3(_05353_ ), .A4(_05352_ ), .ZN(_07642_ ) );
AOI211_X1 _15649_ ( .A(_07638_ ), .B(_07642_ ), .C1(_05358_ ), .C2(_05352_ ), .ZN(_07643_ ) );
AND2_X1 _15650_ ( .A1(_07637_ ), .A2(_07643_ ), .ZN(_07644_ ) );
INV_X1 _15651_ ( .A(_05161_ ), .ZN(_07645_ ) );
OR4_X1 _15652_ ( .A1(_05154_ ), .A2(_07644_ ), .A3(_05155_ ), .A4(_07645_ ), .ZN(_07646_ ) );
INV_X1 _15653_ ( .A(_05148_ ), .ZN(_07647_ ) );
AND2_X1 _15654_ ( .A1(_05159_ ), .A2(_02448_ ), .ZN(_07648_ ) );
AOI21_X1 _15655_ ( .A(_05154_ ), .B1(_07648_ ), .B2(_05156_ ), .ZN(_07649_ ) );
AND3_X1 _15656_ ( .A1(_07646_ ), .A2(_07647_ ), .A3(_07649_ ), .ZN(_07650_ ) );
AOI21_X1 _15657_ ( .A(_07647_ ), .B1(_07646_ ), .B2(_07649_ ), .ZN(_07651_ ) );
OR3_X1 _15658_ ( .A1(_07650_ ), .A2(_07651_ ), .A3(_06880_ ), .ZN(_07652_ ) );
AND4_X1 _15659_ ( .A1(_06935_ ), .A2(_06916_ ), .A3(_06925_ ), .A4(_06931_ ), .ZN(_07653_ ) );
NOR2_X1 _15660_ ( .A1(_07213_ ), .A2(_07653_ ), .ZN(_07654_ ) );
INV_X1 _15661_ ( .A(_07654_ ), .ZN(_07655_ ) );
OAI211_X1 _15662_ ( .A(_06926_ ), .B(_07502_ ), .C1(_06928_ ), .C2(_06931_ ), .ZN(_07656_ ) );
INV_X1 _15663_ ( .A(_07656_ ), .ZN(_07657_ ) );
AND2_X1 _15664_ ( .A1(_07513_ ), .A2(_07008_ ), .ZN(_07658_ ) );
AND2_X1 _15665_ ( .A1(_07658_ ), .A2(_06986_ ), .ZN(_07659_ ) );
OR2_X1 _15666_ ( .A1(_07657_ ), .A2(_07659_ ), .ZN(_07660_ ) );
OAI21_X1 _15667_ ( .A(_06882_ ), .B1(_07655_ ), .B2(_07660_ ), .ZN(_07661_ ) );
OR3_X1 _15668_ ( .A1(_07523_ ), .A2(_06995_ ), .A3(_07525_ ), .ZN(_07662_ ) );
AND2_X1 _15669_ ( .A1(_07108_ ), .A2(_07120_ ), .ZN(_07663_ ) );
AOI21_X1 _15670_ ( .A(_07122_ ), .B1(_05389_ ), .B2(_06975_ ), .ZN(_07664_ ) );
MUX2_X1 _15671_ ( .A(_07663_ ), .B(_07664_ ), .S(_07033_ ), .Z(_07665_ ) );
OR2_X1 _15672_ ( .A1(_07665_ ), .A2(_06981_ ), .ZN(_07666_ ) );
NOR2_X1 _15673_ ( .A1(_07106_ ), .A2(_07103_ ), .ZN(_07667_ ) );
NAND2_X1 _15674_ ( .A1(_07667_ ), .A2(_07142_ ), .ZN(_07668_ ) );
OR3_X1 _15675_ ( .A1(_07102_ ), .A2(_07033_ ), .A3(_07115_ ), .ZN(_07669_ ) );
NAND3_X1 _15676_ ( .A1(_07668_ ), .A2(_07669_ ), .A3(_07255_ ), .ZN(_07670_ ) );
NAND3_X1 _15677_ ( .A1(_07666_ ), .A2(_07010_ ), .A3(_07670_ ), .ZN(_07671_ ) );
OAI21_X1 _15678_ ( .A(_06939_ ), .B1(_07114_ ), .B2(_07112_ ), .ZN(_07672_ ) );
OAI21_X1 _15679_ ( .A(_07011_ ), .B1(_07111_ ), .B2(_07179_ ), .ZN(_07673_ ) );
AND3_X1 _15680_ ( .A1(_07672_ ), .A2(_07673_ ), .A3(_07004_ ), .ZN(_07674_ ) );
AOI21_X1 _15681_ ( .A(_07004_ ), .B1(_07319_ ), .B2(_07320_ ), .ZN(_07675_ ) );
OAI21_X1 _15682_ ( .A(_07042_ ), .B1(_07674_ ), .B2(_07675_ ), .ZN(_07676_ ) );
NAND3_X1 _15683_ ( .A1(_07671_ ), .A2(_06996_ ), .A3(_07676_ ), .ZN(_07677_ ) );
NAND3_X1 _15684_ ( .A1(_07662_ ), .A2(_07677_ ), .A3(_05464_ ), .ZN(_07678_ ) );
NAND3_X1 _15685_ ( .A1(_07658_ ), .A2(_07234_ ), .A3(_06992_ ), .ZN(_07679_ ) );
NAND3_X1 _15686_ ( .A1(_07661_ ), .A2(_07678_ ), .A3(_07679_ ), .ZN(_07680_ ) );
AND2_X1 _15687_ ( .A1(_05148_ ), .A2(_07068_ ), .ZN(_07681_ ) );
INV_X1 _15688_ ( .A(_05147_ ), .ZN(_07682_ ) );
NOR3_X1 _15689_ ( .A1(_02401_ ), .A2(_07682_ ), .A3(_07065_ ), .ZN(_07683_ ) );
AOI21_X1 _15690_ ( .A(_07129_ ), .B1(_02401_ ), .B2(_07682_ ), .ZN(_07684_ ) );
NOR4_X1 _15691_ ( .A1(_07680_ ), .A2(_07681_ ), .A3(_07683_ ), .A4(_07684_ ), .ZN(_07685_ ) );
AOI21_X1 _15692_ ( .A(_07076_ ), .B1(_07652_ ), .B2(_07685_ ), .ZN(_07686_ ) );
OAI21_X1 _15693_ ( .A(_07609_ ), .B1(_07622_ ), .B2(_07686_ ), .ZN(_07687_ ) );
OAI21_X1 _15694_ ( .A(_07608_ ), .B1(_07687_ ), .B2(_06628_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
NAND2_X1 _15695_ ( .A1(_05829_ ), .A2(_06494_ ), .ZN(_07688_ ) );
NAND2_X1 _15696_ ( .A1(_07438_ ), .A2(_04902_ ), .ZN(_07689_ ) );
AND2_X1 _15697_ ( .A1(_07689_ ), .A2(_05416_ ), .ZN(_07690_ ) );
OAI21_X1 _15698_ ( .A(_05415_ ), .B1(_07690_ ), .B2(_04926_ ), .ZN(_07691_ ) );
NAND2_X1 _15699_ ( .A1(_07691_ ), .A2(_04878_ ), .ZN(_07692_ ) );
OAI21_X1 _15700_ ( .A(_07692_ ), .B1(_06838_ ), .B2(_04877_ ), .ZN(_07693_ ) );
XOR2_X1 _15701_ ( .A(_07693_ ), .B(_04855_ ), .Z(_07694_ ) );
NAND2_X1 _15702_ ( .A1(_07694_ ), .A2(_07445_ ), .ZN(_07695_ ) );
NOR2_X1 _15703_ ( .A1(_05819_ ), .A2(_06788_ ), .ZN(_07696_ ) );
AOI21_X1 _15704_ ( .A(_07696_ ), .B1(\ID_EX_imm [11] ), .B2(_07087_ ), .ZN(_07697_ ) );
AOI21_X1 _15705_ ( .A(_06803_ ), .B1(_07695_ ), .B2(_07697_ ), .ZN(_07698_ ) );
NAND2_X1 _15706_ ( .A1(_06826_ ), .A2(_06830_ ), .ZN(_07699_ ) );
AOI21_X1 _15707_ ( .A(_05196_ ), .B1(_07699_ ), .B2(_06836_ ), .ZN(_07700_ ) );
OR3_X1 _15708_ ( .A1(_07700_ ), .A2(_05190_ ), .A3(_06839_ ), .ZN(_07701_ ) );
OAI21_X1 _15709_ ( .A(_05190_ ), .B1(_07700_ ), .B2(_06839_ ), .ZN(_07702_ ) );
NAND3_X1 _15710_ ( .A1(_07701_ ), .A2(_06878_ ), .A3(_07702_ ), .ZN(_07703_ ) );
AND2_X1 _15711_ ( .A1(_07229_ ), .A2(_07009_ ), .ZN(_07704_ ) );
OR2_X1 _15712_ ( .A1(_07704_ ), .A2(_06987_ ), .ZN(_07705_ ) );
NOR2_X1 _15713_ ( .A1(_07222_ ), .A2(_07315_ ), .ZN(_07706_ ) );
OAI21_X1 _15714_ ( .A(_07140_ ), .B1(_07462_ ), .B2(_07463_ ), .ZN(_07707_ ) );
NOR3_X1 _15715_ ( .A1(_07181_ ), .A2(_07018_ ), .A3(_07016_ ), .ZN(_07708_ ) );
NOR3_X1 _15716_ ( .A1(_07014_ ), .A2(_07030_ ), .A3(_07141_ ), .ZN(_07709_ ) );
OAI21_X1 _15717_ ( .A(_07005_ ), .B1(_07708_ ), .B2(_07709_ ), .ZN(_07710_ ) );
AND3_X1 _15718_ ( .A1(_07707_ ), .A2(_07054_ ), .A3(_07710_ ), .ZN(_07711_ ) );
OAI21_X1 _15719_ ( .A(_06987_ ), .B1(_07706_ ), .B2(_07711_ ), .ZN(_07712_ ) );
NAND3_X1 _15720_ ( .A1(_07705_ ), .A2(_06992_ ), .A3(_07712_ ), .ZN(_07713_ ) );
OR2_X1 _15721_ ( .A1(_05189_ ), .A2(_07129_ ), .ZN(_07714_ ) );
NAND3_X1 _15722_ ( .A1(_07262_ ), .A2(_07266_ ), .A3(_07008_ ), .ZN(_07715_ ) );
NAND3_X1 _15723_ ( .A1(_07272_ ), .A2(_06983_ ), .A3(_07005_ ), .ZN(_07716_ ) );
AOI21_X1 _15724_ ( .A(_07559_ ), .B1(_07715_ ), .B2(_07716_ ), .ZN(_07717_ ) );
AOI221_X4 _15725_ ( .A(_07717_ ), .B1(_05188_ ), .B2(_06875_ ), .C1(_05190_ ), .C2(_05467_ ), .ZN(_07718_ ) );
AND4_X1 _15726_ ( .A1(_07703_ ), .A2(_07713_ ), .A3(_07714_ ), .A4(_07718_ ), .ZN(_07719_ ) );
NAND4_X1 _15727_ ( .A1(_06916_ ), .A2(_06925_ ), .A3(_07214_ ), .A4(_07501_ ), .ZN(_07720_ ) );
NAND2_X1 _15728_ ( .A1(_07705_ ), .A2(_07712_ ), .ZN(_07721_ ) );
OAI211_X1 _15729_ ( .A(_07720_ ), .B(_07721_ ), .C1(_06936_ ), .C2(_07499_ ), .ZN(_07722_ ) );
NAND2_X1 _15730_ ( .A1(_07722_ ), .A2(_06883_ ), .ZN(_07723_ ) );
AOI21_X1 _15731_ ( .A(_07076_ ), .B1(_07719_ ), .B2(_07723_ ), .ZN(_07724_ ) );
NOR3_X1 _15732_ ( .A1(_07698_ ), .A2(_05553_ ), .A3(_07724_ ), .ZN(_07725_ ) );
NAND2_X1 _15733_ ( .A1(_05814_ ), .A2(_05553_ ), .ZN(_07726_ ) );
NAND2_X1 _15734_ ( .A1(_07726_ ), .A2(_06563_ ), .ZN(_07727_ ) );
OAI21_X1 _15735_ ( .A(_07688_ ), .B1(_07725_ ), .B2(_07727_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OR2_X1 _15736_ ( .A1(_05888_ ), .A2(_06491_ ), .ZN(_07728_ ) );
AOI21_X1 _15737_ ( .A(_07089_ ), .B1(_07691_ ), .B2(_04878_ ), .ZN(_07729_ ) );
OAI21_X1 _15738_ ( .A(_07729_ ), .B1(_04878_ ), .B2(_07691_ ), .ZN(_07730_ ) );
AOI22_X1 _15739_ ( .A1(_05893_ ), .A2(_07083_ ), .B1(\ID_EX_imm [10] ), .B2(_07086_ ), .ZN(_07731_ ) );
AOI21_X1 _15740_ ( .A(_07281_ ), .B1(_07730_ ), .B2(_07731_ ), .ZN(_07732_ ) );
OR2_X1 _15741_ ( .A1(_07732_ ), .A2(_05552_ ), .ZN(_07733_ ) );
NAND3_X1 _15742_ ( .A1(_07304_ ), .A2(_07061_ ), .A3(_07055_ ), .ZN(_07734_ ) );
OAI21_X1 _15743_ ( .A(_07033_ ), .B1(_07156_ ), .B2(_07163_ ), .ZN(_07735_ ) );
OAI21_X1 _15744_ ( .A(_07036_ ), .B1(_07161_ ), .B2(_07170_ ), .ZN(_07736_ ) );
AOI21_X1 _15745_ ( .A(_07140_ ), .B1(_07735_ ), .B2(_07736_ ), .ZN(_07737_ ) );
AOI21_X1 _15746_ ( .A(_07005_ ), .B1(_07508_ ), .B2(_07509_ ), .ZN(_07738_ ) );
OAI21_X1 _15747_ ( .A(_07010_ ), .B1(_07737_ ), .B2(_07738_ ), .ZN(_07739_ ) );
OAI211_X1 _15748_ ( .A(_06996_ ), .B(_07739_ ), .C1(_07298_ ), .C2(_07055_ ), .ZN(_07740_ ) );
AOI21_X1 _15749_ ( .A(_07557_ ), .B1(_07734_ ), .B2(_07740_ ), .ZN(_07741_ ) );
NAND2_X1 _15750_ ( .A1(_07334_ ), .A2(_07055_ ), .ZN(_07742_ ) );
OAI21_X1 _15751_ ( .A(_07415_ ), .B1(_07313_ ), .B2(_07255_ ), .ZN(_07743_ ) );
AND3_X1 _15752_ ( .A1(_07742_ ), .A2(_07743_ ), .A3(_07480_ ), .ZN(_07744_ ) );
OAI211_X1 _15753_ ( .A(_07287_ ), .B(_07501_ ), .C1(_07036_ ), .C2(_06941_ ), .ZN(_07745_ ) );
INV_X1 _15754_ ( .A(_07500_ ), .ZN(_07746_ ) );
NAND4_X1 _15755_ ( .A1(_07745_ ), .A2(_07746_ ), .A3(_07740_ ), .A4(_07734_ ), .ZN(_07747_ ) );
AOI211_X1 _15756_ ( .A(_07741_ ), .B(_07744_ ), .C1(_07747_ ), .C2(_06883_ ), .ZN(_07748_ ) );
AND3_X1 _15757_ ( .A1(_07699_ ), .A2(_05196_ ), .A3(_06836_ ), .ZN(_07749_ ) );
OR3_X1 _15758_ ( .A1(_07749_ ), .A2(_07700_ ), .A3(_06880_ ), .ZN(_07750_ ) );
AND2_X1 _15759_ ( .A1(_05195_ ), .A2(_07192_ ), .ZN(_07751_ ) );
AOI21_X1 _15760_ ( .A(_07130_ ), .B1(_05194_ ), .B2(_06838_ ), .ZN(_07752_ ) );
NOR3_X1 _15761_ ( .A1(_05194_ ), .A2(_06838_ ), .A3(_07190_ ), .ZN(_07753_ ) );
NOR3_X1 _15762_ ( .A1(_07751_ ), .A2(_07752_ ), .A3(_07753_ ), .ZN(_07754_ ) );
NAND3_X1 _15763_ ( .A1(_07748_ ), .A2(_07750_ ), .A3(_07754_ ), .ZN(_07755_ ) );
BUF_X4 _15764_ ( .A(_07077_ ), .Z(_07756_ ) );
AOI21_X1 _15765_ ( .A(_07733_ ), .B1(_07755_ ), .B2(_07756_ ), .ZN(_07757_ ) );
OAI21_X1 _15766_ ( .A(_07080_ ), .B1(_05891_ ), .B2(_05921_ ), .ZN(_07758_ ) );
OAI21_X1 _15767_ ( .A(_07728_ ), .B1(_07757_ ), .B2(_07758_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
NAND2_X1 _15768_ ( .A1(_05914_ ), .A2(_06494_ ), .ZN(_07759_ ) );
AND4_X1 _15769_ ( .A1(_06942_ ), .A2(_07287_ ), .A3(_06934_ ), .A4(_07501_ ), .ZN(_07760_ ) );
OAI21_X1 _15770_ ( .A(_07060_ ), .B1(_07365_ ), .B2(_07414_ ), .ZN(_07761_ ) );
NAND3_X1 _15771_ ( .A1(_07548_ ), .A2(_06944_ ), .A3(_07549_ ), .ZN(_07762_ ) );
OR3_X1 _15772_ ( .A1(_07018_ ), .A2(_07016_ ), .A3(_07020_ ), .ZN(_07763_ ) );
NOR2_X1 _15773_ ( .A1(_06997_ ), .A2(_07019_ ), .ZN(_07764_ ) );
NAND2_X1 _15774_ ( .A1(_07764_ ), .A2(_07141_ ), .ZN(_07765_ ) );
NAND3_X1 _15775_ ( .A1(_07763_ ), .A2(_07765_ ), .A3(_06951_ ), .ZN(_07766_ ) );
NAND3_X1 _15776_ ( .A1(_07762_ ), .A2(_07766_ ), .A3(_07008_ ), .ZN(_07767_ ) );
OAI211_X1 _15777_ ( .A(_06986_ ), .B(_07767_ ), .C1(_07361_ ), .C2(_07009_ ), .ZN(_07768_ ) );
NAND2_X1 _15778_ ( .A1(_07761_ ), .A2(_07768_ ), .ZN(_07769_ ) );
OAI21_X1 _15779_ ( .A(_07769_ ), .B1(_06936_ ), .B2(_07499_ ), .ZN(_07770_ ) );
OAI21_X1 _15780_ ( .A(_06884_ ), .B1(_07760_ ), .B2(_07770_ ), .ZN(_07771_ ) );
NAND3_X1 _15781_ ( .A1(_07377_ ), .A2(_07378_ ), .A3(_05233_ ), .ZN(_07772_ ) );
NAND3_X1 _15782_ ( .A1(_07057_ ), .A2(_05223_ ), .A3(_06950_ ), .ZN(_07773_ ) );
AOI21_X1 _15783_ ( .A(_07559_ ), .B1(_07772_ ), .B2(_07773_ ), .ZN(_07774_ ) );
AOI221_X4 _15784_ ( .A(_07774_ ), .B1(_05202_ ), .B2(_06875_ ), .C1(_05204_ ), .C2(_05467_ ), .ZN(_07775_ ) );
OAI21_X1 _15785_ ( .A(_07775_ ), .B1(_07557_ ), .B2(_07769_ ), .ZN(_07776_ ) );
AOI21_X1 _15786_ ( .A(_06829_ ), .B1(_06817_ ), .B2(_06824_ ), .ZN(_07777_ ) );
NOR3_X1 _15787_ ( .A1(_07777_ ), .A2(_05204_ ), .A3(_06835_ ), .ZN(_07778_ ) );
NOR2_X1 _15788_ ( .A1(_07778_ ), .A2(_06879_ ), .ZN(_07779_ ) );
OAI21_X1 _15789_ ( .A(_05204_ ), .B1(_07777_ ), .B2(_06835_ ), .ZN(_07780_ ) );
AOI221_X4 _15790_ ( .A(_07776_ ), .B1(_06834_ ), .B2(_05129_ ), .C1(_07779_ ), .C2(_07780_ ), .ZN(_07781_ ) );
AOI21_X1 _15791_ ( .A(_07076_ ), .B1(_07771_ ), .B2(_07781_ ), .ZN(_07782_ ) );
XNOR2_X1 _15792_ ( .A(_07690_ ), .B(_04927_ ), .ZN(_07783_ ) );
NAND2_X1 _15793_ ( .A1(_07783_ ), .A2(_07445_ ), .ZN(_07784_ ) );
AOI22_X1 _15794_ ( .A1(_05903_ ), .A2(_07084_ ), .B1(\ID_EX_imm [9] ), .B2(_07087_ ), .ZN(_07785_ ) );
AOI21_X1 _15795_ ( .A(_06803_ ), .B1(_07784_ ), .B2(_07785_ ), .ZN(_07786_ ) );
NOR3_X1 _15796_ ( .A1(_07782_ ), .A2(_05553_ ), .A3(_07786_ ), .ZN(_07787_ ) );
BUF_X4 _15797_ ( .A(_05479_ ), .Z(_07788_ ) );
OAI21_X1 _15798_ ( .A(_07080_ ), .B1(_05900_ ), .B2(_07788_ ), .ZN(_07789_ ) );
OAI21_X1 _15799_ ( .A(_07759_ ), .B1(_07787_ ), .B2(_07789_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
NAND2_X1 _15800_ ( .A1(_05929_ ), .A2(_06494_ ), .ZN(_07790_ ) );
OAI211_X1 _15801_ ( .A(_06929_ ), .B(_06930_ ), .C1(_07257_ ), .C2(_06887_ ), .ZN(_07791_ ) );
OAI211_X1 _15802_ ( .A(_07159_ ), .B(_07137_ ), .C1(_03045_ ), .C2(_06975_ ), .ZN(_07792_ ) );
NAND3_X1 _15803_ ( .A1(_07157_ ), .A2(_07011_ ), .A3(_07164_ ), .ZN(_07793_ ) );
AOI21_X1 _15804_ ( .A(_06943_ ), .B1(_07792_ ), .B2(_07793_ ), .ZN(_07794_ ) );
AOI211_X1 _15805_ ( .A(_07042_ ), .B(_07794_ ), .C1(_07255_ ), .C2(_07585_ ), .ZN(_07795_ ) );
NOR3_X1 _15806_ ( .A1(_07403_ ), .A2(_07404_ ), .A3(_07010_ ), .ZN(_07796_ ) );
OAI21_X1 _15807_ ( .A(_06996_ ), .B1(_07795_ ), .B2(_07796_ ), .ZN(_07797_ ) );
OAI21_X1 _15808_ ( .A(_07061_ ), .B1(_07407_ ), .B2(_07415_ ), .ZN(_07798_ ) );
NAND2_X1 _15809_ ( .A1(_07797_ ), .A2(_07798_ ), .ZN(_07799_ ) );
AOI21_X1 _15810_ ( .A(_07544_ ), .B1(_07791_ ), .B2(_07799_ ), .ZN(_07800_ ) );
NOR2_X1 _15811_ ( .A1(_07777_ ), .A2(_06879_ ), .ZN(_07801_ ) );
OAI21_X1 _15812_ ( .A(_07801_ ), .B1(_05208_ ), .B2(_06826_ ), .ZN(_07802_ ) );
NAND3_X1 _15813_ ( .A1(_07797_ ), .A2(_06993_ ), .A3(_07798_ ), .ZN(_07803_ ) );
OAI21_X1 _15814_ ( .A(_05129_ ), .B1(_05279_ ), .B2(_03045_ ), .ZN(_07804_ ) );
NAND2_X1 _15815_ ( .A1(_07413_ ), .A2(_07009_ ), .ZN(_07805_ ) );
AND2_X1 _15816_ ( .A1(_06941_ ), .A2(_05116_ ), .ZN(_07806_ ) );
NAND4_X1 _15817_ ( .A1(_07806_ ), .A2(_06983_ ), .A3(_07005_ ), .A4(_07142_ ), .ZN(_07807_ ) );
AOI21_X1 _15818_ ( .A(_07559_ ), .B1(_07805_ ), .B2(_07807_ ), .ZN(_07808_ ) );
AOI221_X4 _15819_ ( .A(_07808_ ), .B1(_06835_ ), .B2(_06875_ ), .C1(_05208_ ), .C2(_07068_ ), .ZN(_07809_ ) );
NAND4_X1 _15820_ ( .A1(_07802_ ), .A2(_07803_ ), .A3(_07804_ ), .A4(_07809_ ), .ZN(_07810_ ) );
OAI21_X1 _15821_ ( .A(_07077_ ), .B1(_07800_ ), .B2(_07810_ ), .ZN(_07811_ ) );
AOI21_X1 _15822_ ( .A(_07207_ ), .B1(_07438_ ), .B2(_04902_ ), .ZN(_07812_ ) );
OAI21_X1 _15823_ ( .A(_07812_ ), .B1(_04902_ ), .B2(_07438_ ), .ZN(_07813_ ) );
AOI22_X1 _15824_ ( .A1(_05930_ ), .A2(_07084_ ), .B1(\ID_EX_imm [8] ), .B2(_07087_ ), .ZN(_07814_ ) );
NAND2_X1 _15825_ ( .A1(_07813_ ), .A2(_07814_ ), .ZN(_07815_ ) );
BUF_X4 _15826_ ( .A(_06801_ ), .Z(_07816_ ) );
NAND2_X1 _15827_ ( .A1(_07815_ ), .A2(_07816_ ), .ZN(_07817_ ) );
AND3_X1 _15828_ ( .A1(_07811_ ), .A2(_05601_ ), .A3(_07817_ ), .ZN(_07818_ ) );
NAND2_X1 _15829_ ( .A1(_05932_ ), .A2(_05838_ ), .ZN(_07819_ ) );
NAND2_X1 _15830_ ( .A1(_07819_ ), .A2(_06563_ ), .ZN(_07820_ ) );
OAI21_X1 _15831_ ( .A(_07790_ ), .B1(_07818_ ), .B2(_07820_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
NAND2_X1 _15832_ ( .A1(_05943_ ), .A2(_06494_ ), .ZN(_07821_ ) );
AND3_X1 _15833_ ( .A1(_05399_ ), .A2(_05400_ ), .A3(_05401_ ), .ZN(_07822_ ) );
NOR2_X1 _15834_ ( .A1(_07822_ ), .A2(_05406_ ), .ZN(_07823_ ) );
OR2_X1 _15835_ ( .A1(_07823_ ), .A2(_05070_ ), .ZN(_07824_ ) );
NAND2_X1 _15836_ ( .A1(_02788_ ), .A2(_05069_ ), .ZN(_07825_ ) );
AND3_X1 _15837_ ( .A1(_07824_ ), .A2(_05048_ ), .A3(_07825_ ), .ZN(_07826_ ) );
AOI21_X1 _15838_ ( .A(_05048_ ), .B1(_07824_ ), .B2(_07825_ ), .ZN(_07827_ ) );
OR3_X1 _15839_ ( .A1(_07826_ ), .A2(_07827_ ), .A3(_07089_ ), .ZN(_07828_ ) );
AOI22_X1 _15840_ ( .A1(_05948_ ), .A2(_07083_ ), .B1(\ID_EX_imm [7] ), .B2(_07086_ ), .ZN(_07829_ ) );
AOI21_X1 _15841_ ( .A(_07281_ ), .B1(_07828_ ), .B2(_07829_ ), .ZN(_07830_ ) );
OR2_X1 _15842_ ( .A1(_07830_ ), .A2(_05552_ ), .ZN(_07831_ ) );
AND4_X1 _15843_ ( .A1(_05214_ ), .A2(_06814_ ), .A3(_06815_ ), .A4(_05220_ ), .ZN(_07832_ ) );
OR2_X1 _15844_ ( .A1(_07832_ ), .A2(_06822_ ), .ZN(_07833_ ) );
AND2_X1 _15845_ ( .A1(_07833_ ), .A2(_05260_ ), .ZN(_07834_ ) );
OR3_X1 _15846_ ( .A1(_07834_ ), .A2(_05256_ ), .A3(_06819_ ), .ZN(_07835_ ) );
OAI21_X1 _15847_ ( .A(_05256_ ), .B1(_07834_ ), .B2(_06819_ ), .ZN(_07836_ ) );
NAND3_X1 _15848_ ( .A1(_07835_ ), .A2(_07246_ ), .A3(_07836_ ), .ZN(_07837_ ) );
NAND4_X1 _15849_ ( .A1(_06933_ ), .A2(_06884_ ), .A3(_06935_ ), .A4(_07501_ ), .ZN(_07838_ ) );
OR3_X1 _15850_ ( .A1(_07468_ ), .A2(_06984_ ), .A3(_07469_ ), .ZN(_07839_ ) );
NAND4_X1 _15851_ ( .A1(_06979_ ), .A2(_07414_ ), .A3(_07006_ ), .A4(_07142_ ), .ZN(_07840_ ) );
AND3_X1 _15852_ ( .A1(_07839_ ), .A2(_07146_ ), .A3(_07840_ ), .ZN(_07841_ ) );
NOR2_X1 _15853_ ( .A1(_07708_ ), .A2(_07709_ ), .ZN(_07842_ ) );
NOR3_X1 _15854_ ( .A1(_07181_ ), .A2(_07000_ ), .A3(_06998_ ), .ZN(_07843_ ) );
NOR3_X1 _15855_ ( .A1(_06997_ ), .A2(_07019_ ), .A3(_07141_ ), .ZN(_07844_ ) );
NOR2_X1 _15856_ ( .A1(_07843_ ), .A2(_07844_ ), .ZN(_07845_ ) );
MUX2_X1 _15857_ ( .A(_07842_ ), .B(_07845_ ), .S(_07024_ ), .Z(_07846_ ) );
MUX2_X1 _15858_ ( .A(_07466_ ), .B(_07846_ ), .S(_07010_ ), .Z(_07847_ ) );
AOI211_X1 _15859_ ( .A(_07461_ ), .B(_07841_ ), .C1(_06988_ ), .C2(_07847_ ), .ZN(_07848_ ) );
NOR3_X1 _15860_ ( .A1(_07474_ ), .A2(_07257_ ), .A3(_07559_ ), .ZN(_07849_ ) );
NOR3_X1 _15861_ ( .A1(_05263_ ), .A2(_05264_ ), .A3(_05468_ ), .ZN(_07850_ ) );
NAND3_X1 _15862_ ( .A1(_05266_ ), .A2(_02812_ ), .A3(_06875_ ), .ZN(_07851_ ) );
OAI21_X1 _15863_ ( .A(_07851_ ), .B1(_05263_ ), .B2(_07129_ ), .ZN(_07852_ ) );
NOR4_X1 _15864_ ( .A1(_07848_ ), .A2(_07849_ ), .A3(_07850_ ), .A4(_07852_ ), .ZN(_07853_ ) );
NAND3_X1 _15865_ ( .A1(_07837_ ), .A2(_07838_ ), .A3(_07853_ ), .ZN(_07854_ ) );
AOI21_X1 _15866_ ( .A(_07831_ ), .B1(_07854_ ), .B2(_07756_ ), .ZN(_07855_ ) );
OAI21_X1 _15867_ ( .A(_07080_ ), .B1(_05945_ ), .B2(_07788_ ), .ZN(_07856_ ) );
OAI21_X1 _15868_ ( .A(_07821_ ), .B1(_07855_ ), .B2(_07856_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
OR2_X1 _15869_ ( .A1(_05972_ ), .A2(_06491_ ), .ZN(_07857_ ) );
NAND2_X1 _15870_ ( .A1(_07823_ ), .A2(_05070_ ), .ZN(_07858_ ) );
NAND3_X1 _15871_ ( .A1(_07824_ ), .A2(_07445_ ), .A3(_07858_ ), .ZN(_07859_ ) );
AOI22_X1 _15872_ ( .A1(_05960_ ), .A2(_07083_ ), .B1(\ID_EX_imm [6] ), .B2(_07086_ ), .ZN(_07860_ ) );
AOI21_X1 _15873_ ( .A(_07281_ ), .B1(_07859_ ), .B2(_07860_ ), .ZN(_07861_ ) );
OR2_X1 _15874_ ( .A1(_07861_ ), .A2(_05552_ ), .ZN(_07862_ ) );
NAND3_X1 _15875_ ( .A1(_06916_ ), .A2(_06925_ ), .A3(_07502_ ), .ZN(_07863_ ) );
NOR3_X1 _15876_ ( .A1(_07863_ ), .A2(_06934_ ), .A3(_07499_ ), .ZN(_07864_ ) );
NAND3_X1 _15877_ ( .A1(_07504_ ), .A2(_05233_ ), .A3(_07505_ ), .ZN(_07865_ ) );
OAI21_X1 _15878_ ( .A(_07865_ ), .B1(_07008_ ), .B2(_07514_ ), .ZN(_07866_ ) );
AND2_X1 _15879_ ( .A1(_07866_ ), .A2(_07146_ ), .ZN(_07867_ ) );
OAI21_X1 _15880_ ( .A(_07033_ ), .B1(_07151_ ), .B2(_07149_ ), .ZN(_07868_ ) );
OAI21_X1 _15881_ ( .A(_07036_ ), .B1(_07148_ ), .B2(_07158_ ), .ZN(_07869_ ) );
NAND3_X1 _15882_ ( .A1(_07868_ ), .A2(_07869_ ), .A3(_07024_ ), .ZN(_07870_ ) );
NAND3_X1 _15883_ ( .A1(_07735_ ), .A2(_07736_ ), .A3(_06981_ ), .ZN(_07871_ ) );
AND3_X1 _15884_ ( .A1(_07870_ ), .A2(_07871_ ), .A3(_07054_ ), .ZN(_07872_ ) );
AOI211_X1 _15885_ ( .A(_07146_ ), .B(_07872_ ), .C1(_07511_ ), .C2(_07415_ ), .ZN(_07873_ ) );
OR2_X1 _15886_ ( .A1(_07867_ ), .A2(_07873_ ), .ZN(_07874_ ) );
OAI21_X1 _15887_ ( .A(_06884_ ), .B1(_07864_ ), .B2(_07874_ ), .ZN(_07875_ ) );
AOI21_X1 _15888_ ( .A(_06880_ ), .B1(_07833_ ), .B2(_05260_ ), .ZN(_07876_ ) );
OAI21_X1 _15889_ ( .A(_07876_ ), .B1(_05260_ ), .B2(_07833_ ), .ZN(_07877_ ) );
AOI21_X1 _15890_ ( .A(_07130_ ), .B1(_05259_ ), .B2(_06818_ ), .ZN(_07878_ ) );
OR3_X1 _15891_ ( .A1(_07524_ ), .A2(_07415_ ), .A3(_07559_ ), .ZN(_07879_ ) );
NAND2_X1 _15892_ ( .A1(_05260_ ), .A2(_07068_ ), .ZN(_07880_ ) );
NAND2_X1 _15893_ ( .A1(_06819_ ), .A2(_07368_ ), .ZN(_07881_ ) );
NAND3_X1 _15894_ ( .A1(_07879_ ), .A2(_07880_ ), .A3(_07881_ ), .ZN(_07882_ ) );
AOI211_X1 _15895_ ( .A(_07878_ ), .B(_07882_ ), .C1(_07874_ ), .C2(_06993_ ), .ZN(_07883_ ) );
NAND3_X1 _15896_ ( .A1(_07875_ ), .A2(_07877_ ), .A3(_07883_ ), .ZN(_07884_ ) );
AOI21_X1 _15897_ ( .A(_07862_ ), .B1(_07884_ ), .B2(_07756_ ), .ZN(_07885_ ) );
OAI21_X1 _15898_ ( .A(_07080_ ), .B1(_05959_ ), .B2(_07788_ ), .ZN(_07886_ ) );
OAI21_X1 _15899_ ( .A(_07857_ ), .B1(_07885_ ), .B2(_07886_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
OR2_X1 _15900_ ( .A1(_05987_ ), .A2(_06491_ ), .ZN(_07887_ ) );
AND3_X1 _15901_ ( .A1(_05399_ ), .A2(_05400_ ), .A3(_04999_ ), .ZN(_07888_ ) );
OR3_X1 _15902_ ( .A1(_07888_ ), .A2(_05092_ ), .A3(_05404_ ), .ZN(_07889_ ) );
OAI21_X1 _15903_ ( .A(_05092_ ), .B1(_07888_ ), .B2(_05404_ ), .ZN(_07890_ ) );
NAND3_X1 _15904_ ( .A1(_07889_ ), .A2(_07445_ ), .A3(_07890_ ), .ZN(_07891_ ) );
AOI22_X1 _15905_ ( .A1(_05990_ ), .A2(_07083_ ), .B1(\ID_EX_imm [5] ), .B2(_07086_ ), .ZN(_07892_ ) );
AOI21_X1 _15906_ ( .A(_06802_ ), .B1(_07891_ ), .B2(_07892_ ), .ZN(_07893_ ) );
OR2_X1 _15907_ ( .A1(_07893_ ), .A2(_05552_ ), .ZN(_07894_ ) );
NOR3_X1 _15908_ ( .A1(_06936_ ), .A2(_06945_ ), .A3(_07499_ ), .ZN(_07895_ ) );
NAND2_X1 _15909_ ( .A1(_06985_ ), .A2(_07146_ ), .ZN(_07896_ ) );
AOI21_X1 _15910_ ( .A(_07054_ ), .B1(_07547_ ), .B2(_07550_ ), .ZN(_07897_ ) );
NAND3_X1 _15911_ ( .A1(_07763_ ), .A2(_07765_ ), .A3(_07140_ ), .ZN(_07898_ ) );
OAI21_X1 _15912_ ( .A(_07141_ ), .B1(_07049_ ), .B2(_07001_ ), .ZN(_07899_ ) );
OAI21_X1 _15913_ ( .A(_07181_ ), .B1(_07000_ ), .B2(_06998_ ), .ZN(_07900_ ) );
NAND2_X1 _15914_ ( .A1(_07899_ ), .A2(_07900_ ), .ZN(_07901_ ) );
NAND2_X1 _15915_ ( .A1(_07901_ ), .A2(_07040_ ), .ZN(_07902_ ) );
AOI21_X1 _15916_ ( .A(_06984_ ), .B1(_07898_ ), .B2(_07902_ ), .ZN(_07903_ ) );
OR3_X1 _15917_ ( .A1(_07897_ ), .A2(_07903_ ), .A3(_07060_ ), .ZN(_07904_ ) );
NAND2_X1 _15918_ ( .A1(_07896_ ), .A2(_07904_ ), .ZN(_07905_ ) );
OAI21_X1 _15919_ ( .A(_06883_ ), .B1(_07895_ ), .B2(_07905_ ), .ZN(_07906_ ) );
NAND2_X1 _15920_ ( .A1(_07905_ ), .A2(_06993_ ), .ZN(_07907_ ) );
OR2_X1 _15921_ ( .A1(_07059_ ), .A2(_07559_ ), .ZN(_07908_ ) );
AND3_X1 _15922_ ( .A1(_07906_ ), .A2(_07907_ ), .A3(_07908_ ), .ZN(_07909_ ) );
NAND2_X1 _15923_ ( .A1(_06814_ ), .A2(_06815_ ), .ZN(_07910_ ) );
INV_X1 _15924_ ( .A(_05220_ ), .ZN(_07911_ ) );
NOR2_X1 _15925_ ( .A1(_07910_ ), .A2(_07911_ ), .ZN(_07912_ ) );
NOR2_X1 _15926_ ( .A1(_07912_ ), .A2(_05218_ ), .ZN(_07913_ ) );
XNOR2_X1 _15927_ ( .A(_07913_ ), .B(_05214_ ), .ZN(_07914_ ) );
NAND2_X1 _15928_ ( .A1(_07914_ ), .A2(_07246_ ), .ZN(_07915_ ) );
NAND2_X1 _15929_ ( .A1(_05214_ ), .A2(_07192_ ), .ZN(_07916_ ) );
NAND3_X1 _15930_ ( .A1(_05212_ ), .A2(_02764_ ), .A3(_07368_ ), .ZN(_07917_ ) );
OAI21_X1 _15931_ ( .A(_05129_ ), .B1(_05212_ ), .B2(_02764_ ), .ZN(_07918_ ) );
AND3_X1 _15932_ ( .A1(_07916_ ), .A2(_07917_ ), .A3(_07918_ ), .ZN(_07919_ ) );
NAND3_X1 _15933_ ( .A1(_07909_ ), .A2(_07915_ ), .A3(_07919_ ), .ZN(_07920_ ) );
AOI21_X1 _15934_ ( .A(_07894_ ), .B1(_07920_ ), .B2(_07756_ ), .ZN(_07921_ ) );
NAND2_X1 _15935_ ( .A1(_05992_ ), .A2(_05838_ ), .ZN(_07922_ ) );
NAND2_X1 _15936_ ( .A1(_07922_ ), .A2(_06563_ ), .ZN(_07923_ ) );
OAI21_X1 _15937_ ( .A(_07887_ ), .B1(_07921_ ), .B2(_07923_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
AND2_X1 _15938_ ( .A1(_05999_ ), .A2(_05552_ ), .ZN(_07924_ ) );
NAND4_X1 _15939_ ( .A1(_06933_ ), .A2(_06935_ ), .A3(_07099_ ), .A4(_07501_ ), .ZN(_07925_ ) );
NAND2_X1 _15940_ ( .A1(_07126_ ), .A2(_07060_ ), .ZN(_07926_ ) );
NAND2_X1 _15941_ ( .A1(_07586_ ), .A2(_06984_ ), .ZN(_07927_ ) );
AND3_X1 _15942_ ( .A1(_07792_ ), .A2(_06943_ ), .A3(_07793_ ), .ZN(_07928_ ) );
NOR3_X1 _15943_ ( .A1(_07011_ ), .A2(_07133_ ), .A3(_07152_ ), .ZN(_07929_ ) );
NOR3_X1 _15944_ ( .A1(_07151_ ), .A2(_07149_ ), .A3(_07020_ ), .ZN(_07930_ ) );
NOR2_X1 _15945_ ( .A1(_07929_ ), .A2(_07930_ ), .ZN(_07931_ ) );
AOI21_X1 _15946_ ( .A(_07928_ ), .B1(_07040_ ), .B2(_07931_ ), .ZN(_07932_ ) );
OAI211_X1 _15947_ ( .A(_07927_ ), .B(_06986_ ), .C1(_07414_ ), .C2(_07932_ ), .ZN(_07933_ ) );
AND2_X1 _15948_ ( .A1(_07926_ ), .A2(_07933_ ), .ZN(_07934_ ) );
AOI21_X1 _15949_ ( .A(_07544_ ), .B1(_07925_ ), .B2(_07934_ ), .ZN(_07935_ ) );
NAND3_X1 _15950_ ( .A1(_07146_ ), .A2(_02735_ ), .A3(_06875_ ), .ZN(_07936_ ) );
OAI221_X1 _15951_ ( .A(_07936_ ), .B1(_07911_ ), .B2(_05468_ ), .C1(_07145_ ), .C2(_07559_ ), .ZN(_07937_ ) );
OR2_X1 _15952_ ( .A1(_07935_ ), .A2(_07937_ ), .ZN(_07938_ ) );
AOI21_X1 _15953_ ( .A(_06879_ ), .B1(_07910_ ), .B2(_07911_ ), .ZN(_07939_ ) );
OAI21_X1 _15954_ ( .A(_07939_ ), .B1(_07911_ ), .B2(_07910_ ), .ZN(_07940_ ) );
OAI221_X1 _15955_ ( .A(_07940_ ), .B1(_05219_ ), .B2(_07129_ ), .C1(_07934_ ), .C2(_07557_ ), .ZN(_07941_ ) );
OAI21_X1 _15956_ ( .A(_07077_ ), .B1(_07938_ ), .B2(_07941_ ), .ZN(_07942_ ) );
AOI21_X1 _15957_ ( .A(_04999_ ), .B1(_05399_ ), .B2(_05400_ ), .ZN(_07943_ ) );
NOR3_X1 _15958_ ( .A1(_07888_ ), .A2(_07943_ ), .A3(_07207_ ), .ZN(_07944_ ) );
INV_X1 _15959_ ( .A(_07086_ ), .ZN(_07945_ ) );
OAI22_X1 _15960_ ( .A1(_06002_ ), .A2(_06787_ ), .B1(_02736_ ), .B2(_07945_ ), .ZN(_07946_ ) );
OAI21_X1 _15961_ ( .A(_07816_ ), .B1(_07944_ ), .B2(_07946_ ), .ZN(_07947_ ) );
AND2_X1 _15962_ ( .A1(_07947_ ), .A2(_05600_ ), .ZN(_07948_ ) );
AOI21_X1 _15963_ ( .A(_07924_ ), .B1(_07942_ ), .B2(_07948_ ), .ZN(_07949_ ) );
MUX2_X1 _15964_ ( .A(_06014_ ), .B(_07949_ ), .S(_06502_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
AND3_X1 _15965_ ( .A1(_06033_ ), .A2(\ID_EX_typ [7] ), .A3(_06800_ ), .ZN(_07950_ ) );
NAND4_X1 _15966_ ( .A1(_06933_ ), .A2(_06935_ ), .A3(_07214_ ), .A4(_07501_ ), .ZN(_07951_ ) );
OR2_X1 _15967_ ( .A1(_07230_ ), .A2(_06987_ ), .ZN(_07952_ ) );
NOR3_X1 _15968_ ( .A1(_07049_ ), .A2(_07001_ ), .A3(_07141_ ), .ZN(_07953_ ) );
NOR2_X1 _15969_ ( .A1(_07046_ ), .A2(_07050_ ), .ZN(_07954_ ) );
AOI211_X1 _15970_ ( .A(_06944_ ), .B(_07953_ ), .C1(_07142_ ), .C2(_07954_ ), .ZN(_07955_ ) );
NOR3_X1 _15971_ ( .A1(_07843_ ), .A2(_07844_ ), .A3(_07005_ ), .ZN(_07956_ ) );
NOR3_X1 _15972_ ( .A1(_07955_ ), .A2(_07414_ ), .A3(_07956_ ), .ZN(_07957_ ) );
AOI21_X1 _15973_ ( .A(_07009_ ), .B1(_07707_ ), .B2(_07710_ ), .ZN(_07958_ ) );
OR3_X1 _15974_ ( .A1(_07957_ ), .A2(_07060_ ), .A3(_07958_ ), .ZN(_07959_ ) );
NAND2_X1 _15975_ ( .A1(_07952_ ), .A2(_07959_ ), .ZN(_07960_ ) );
AOI21_X1 _15976_ ( .A(_07544_ ), .B1(_07951_ ), .B2(_07960_ ), .ZN(_07961_ ) );
NAND3_X1 _15977_ ( .A1(_07952_ ), .A2(_06992_ ), .A3(_07959_ ), .ZN(_07962_ ) );
OR3_X1 _15978_ ( .A1(_06812_ ), .A2(_05226_ ), .A3(_06813_ ), .ZN(_07963_ ) );
OAI21_X1 _15979_ ( .A(_05226_ ), .B1(_06812_ ), .B2(_06813_ ), .ZN(_07964_ ) );
NAND3_X1 _15980_ ( .A1(_07963_ ), .A2(_06878_ ), .A3(_07964_ ), .ZN(_07965_ ) );
OAI21_X1 _15981_ ( .A(_05129_ ), .B1(_02910_ ), .B2(_07257_ ), .ZN(_07966_ ) );
NOR2_X1 _15982_ ( .A1(_07273_ ), .A2(_07559_ ), .ZN(_07967_ ) );
AOI221_X4 _15983_ ( .A(_07967_ ), .B1(_05224_ ), .B2(_06875_ ), .C1(_05226_ ), .C2(_05467_ ), .ZN(_07968_ ) );
NAND4_X1 _15984_ ( .A1(_07962_ ), .A2(_07965_ ), .A3(_07966_ ), .A4(_07968_ ), .ZN(_07969_ ) );
OAI21_X1 _15985_ ( .A(_07077_ ), .B1(_07961_ ), .B2(_07969_ ), .ZN(_07970_ ) );
OR2_X1 _15986_ ( .A1(_05397_ ), .A2(_05398_ ), .ZN(_07971_ ) );
AND3_X1 _15987_ ( .A1(_07971_ ), .A2(_04953_ ), .A3(_05395_ ), .ZN(_07972_ ) );
AOI21_X1 _15988_ ( .A(_04953_ ), .B1(_07971_ ), .B2(_05395_ ), .ZN(_07973_ ) );
NOR3_X1 _15989_ ( .A1(_07972_ ), .A2(_07973_ ), .A3(_07207_ ), .ZN(_07974_ ) );
OAI22_X1 _15990_ ( .A1(_06031_ ), .A2(_06787_ ), .B1(_02911_ ), .B2(_07945_ ), .ZN(_07975_ ) );
OAI21_X1 _15991_ ( .A(_07816_ ), .B1(_07974_ ), .B2(_07975_ ), .ZN(_07976_ ) );
AND2_X1 _15992_ ( .A1(_07976_ ), .A2(_05600_ ), .ZN(_07977_ ) );
AOI21_X1 _15993_ ( .A(_07950_ ), .B1(_07970_ ), .B2(_07977_ ), .ZN(_07978_ ) );
MUX2_X1 _15994_ ( .A(_06027_ ), .B(_07978_ ), .S(_06502_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
NAND2_X1 _15995_ ( .A1(_06045_ ), .A2(_06494_ ), .ZN(_07979_ ) );
NAND2_X1 _15996_ ( .A1(_05397_ ), .A2(_05398_ ), .ZN(_07980_ ) );
NAND3_X1 _15997_ ( .A1(_07971_ ), .A2(_07445_ ), .A3(_07980_ ), .ZN(_07981_ ) );
AOI22_X1 _15998_ ( .A1(_06047_ ), .A2(_07083_ ), .B1(\ID_EX_imm [2] ), .B2(_07086_ ), .ZN(_07982_ ) );
AOI21_X1 _15999_ ( .A(_06802_ ), .B1(_07981_ ), .B2(_07982_ ), .ZN(_07983_ ) );
OR2_X1 _16000_ ( .A1(_07983_ ), .A2(_05552_ ), .ZN(_07984_ ) );
NAND2_X1 _16001_ ( .A1(_07305_ ), .A2(_07060_ ), .ZN(_07985_ ) );
OAI21_X1 _16002_ ( .A(_07414_ ), .B1(_07737_ ), .B2(_07738_ ), .ZN(_07986_ ) );
OAI21_X1 _16003_ ( .A(_07036_ ), .B1(_07133_ ), .B2(_07152_ ), .ZN(_07987_ ) );
NOR2_X1 _16004_ ( .A1(_07132_ ), .A2(_07136_ ), .ZN(_07988_ ) );
OAI211_X1 _16005_ ( .A(_07040_ ), .B(_07987_ ), .C1(_07988_ ), .C2(_07036_ ), .ZN(_07989_ ) );
NAND3_X1 _16006_ ( .A1(_07868_ ), .A2(_07869_ ), .A3(_07140_ ), .ZN(_07990_ ) );
NAND3_X1 _16007_ ( .A1(_07989_ ), .A2(_07054_ ), .A3(_07990_ ), .ZN(_07991_ ) );
NAND3_X1 _16008_ ( .A1(_07986_ ), .A2(_06995_ ), .A3(_07991_ ), .ZN(_07992_ ) );
AOI21_X1 _16009_ ( .A(_07557_ ), .B1(_07985_ ), .B2(_07992_ ), .ZN(_07993_ ) );
NOR2_X1 _16010_ ( .A1(_07288_ ), .A2(_07289_ ), .ZN(_07994_ ) );
NAND3_X1 _16011_ ( .A1(_07994_ ), .A2(_06935_ ), .A3(_07501_ ), .ZN(_07995_ ) );
NAND3_X1 _16012_ ( .A1(_07995_ ), .A2(_07992_ ), .A3(_07985_ ), .ZN(_07996_ ) );
AOI221_X4 _16013_ ( .A(_07993_ ), .B1(_07316_ ), .B2(_07480_ ), .C1(_07996_ ), .C2(_06883_ ), .ZN(_07997_ ) );
AOI21_X1 _16014_ ( .A(_06880_ ), .B1(_06811_ ), .B2(_05246_ ), .ZN(_07998_ ) );
OAI21_X1 _16015_ ( .A(_07998_ ), .B1(_05246_ ), .B2(_06811_ ), .ZN(_07999_ ) );
NAND2_X1 _16016_ ( .A1(_05245_ ), .A2(_07192_ ), .ZN(_08000_ ) );
NAND3_X1 _16017_ ( .A1(_07255_ ), .A2(_02886_ ), .A3(_07368_ ), .ZN(_08001_ ) );
OAI21_X1 _16018_ ( .A(_05129_ ), .B1(_07255_ ), .B2(_02886_ ), .ZN(_08002_ ) );
AND3_X1 _16019_ ( .A1(_08000_ ), .A2(_08001_ ), .A3(_08002_ ), .ZN(_08003_ ) );
NAND3_X1 _16020_ ( .A1(_07997_ ), .A2(_07999_ ), .A3(_08003_ ), .ZN(_08004_ ) );
AOI21_X1 _16021_ ( .A(_07984_ ), .B1(_08004_ ), .B2(_07756_ ), .ZN(_08005_ ) );
BUF_X4 _16022_ ( .A(_06491_ ), .Z(_08006_ ) );
OAI21_X1 _16023_ ( .A(_08006_ ), .B1(_05620_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08007_ ) );
OAI21_X1 _16024_ ( .A(_07979_ ), .B1(_08005_ ), .B2(_08007_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
BUF_X4 _16025_ ( .A(_06489_ ), .Z(_08008_ ) );
NAND2_X1 _16026_ ( .A1(_05597_ ), .A2(_08008_ ), .ZN(_08009_ ) );
OAI22_X1 _16027_ ( .A1(_05577_ ), .A2(_06788_ ), .B1(_02426_ ), .B2(_07945_ ), .ZN(_08010_ ) );
NOR2_X1 _16028_ ( .A1(_07615_ ), .A2(_07616_ ), .ZN(_08011_ ) );
AND2_X1 _16029_ ( .A1(_02448_ ), .A2(_05445_ ), .ZN(_08012_ ) );
OR3_X1 _16030_ ( .A1(_08011_ ), .A2(_04584_ ), .A3(_08012_ ), .ZN(_08013_ ) );
OAI21_X1 _16031_ ( .A(_04584_ ), .B1(_08011_ ), .B2(_08012_ ), .ZN(_08014_ ) );
AND3_X1 _16032_ ( .A1(_08013_ ), .A2(_06795_ ), .A3(_08014_ ), .ZN(_08015_ ) );
OAI21_X1 _16033_ ( .A(_07816_ ), .B1(_08010_ ), .B2(_08015_ ), .ZN(_08016_ ) );
NAND2_X1 _16034_ ( .A1(_08016_ ), .A2(_05601_ ), .ZN(_08017_ ) );
NAND3_X1 _16035_ ( .A1(_07560_ ), .A2(_07146_ ), .A3(_07561_ ), .ZN(_08018_ ) );
OAI211_X1 _16036_ ( .A(_07224_ ), .B(_07036_ ), .C1(_03207_ ), .C2(_06941_ ), .ZN(_08019_ ) );
NAND2_X1 _16037_ ( .A1(_07223_ ), .A2(_06977_ ), .ZN(_08020_ ) );
OAI211_X1 _16038_ ( .A(_08019_ ), .B(_07024_ ), .C1(_07036_ ), .C2(_08020_ ), .ZN(_08021_ ) );
NOR2_X1 _16039_ ( .A1(_06966_ ), .A2(_06971_ ), .ZN(_08022_ ) );
NOR2_X1 _16040_ ( .A1(_06952_ ), .A2(_06970_ ), .ZN(_08023_ ) );
MUX2_X1 _16041_ ( .A(_08022_ ), .B(_08023_ ), .S(_07142_ ), .Z(_08024_ ) );
OAI211_X1 _16042_ ( .A(_07010_ ), .B(_08021_ ), .C1(_08024_ ), .C2(_07006_ ), .ZN(_08025_ ) );
OAI21_X1 _16043_ ( .A(_07042_ ), .B1(_07032_ ), .B2(_07041_ ), .ZN(_08026_ ) );
NAND3_X1 _16044_ ( .A1(_08025_ ), .A2(_06987_ ), .A3(_08026_ ), .ZN(_08027_ ) );
AND3_X1 _16045_ ( .A1(_08018_ ), .A2(_05464_ ), .A3(_08027_ ), .ZN(_08028_ ) );
NOR3_X1 _16046_ ( .A1(_06980_ ), .A2(_07414_ ), .A3(_06981_ ), .ZN(_08029_ ) );
AND2_X1 _16047_ ( .A1(_08029_ ), .A2(_06995_ ), .ZN(_08030_ ) );
AOI21_X1 _16048_ ( .A(_08030_ ), .B1(_06929_ ), .B2(_06930_ ), .ZN(_08031_ ) );
OR3_X1 _16049_ ( .A1(_07398_ ), .A2(_07397_ ), .A3(_07545_ ), .ZN(_08032_ ) );
AOI21_X1 _16050_ ( .A(_07544_ ), .B1(_08031_ ), .B2(_08032_ ), .ZN(_08033_ ) );
AOI211_X1 _16051_ ( .A(_08028_ ), .B(_08033_ ), .C1(_06993_ ), .C2(_08030_ ), .ZN(_08034_ ) );
AOI21_X1 _16052_ ( .A(_07645_ ), .B1(_07637_ ), .B2(_07643_ ), .ZN(_08035_ ) );
OR3_X1 _16053_ ( .A1(_08035_ ), .A2(_05156_ ), .A3(_07648_ ), .ZN(_08036_ ) );
OAI21_X1 _16054_ ( .A(_05156_ ), .B1(_08035_ ), .B2(_07648_ ), .ZN(_08037_ ) );
NAND3_X1 _16055_ ( .A1(_08036_ ), .A2(_07246_ ), .A3(_08037_ ), .ZN(_08038_ ) );
NOR3_X1 _16056_ ( .A1(_05154_ ), .A2(_05155_ ), .A3(_05468_ ), .ZN(_08039_ ) );
NOR2_X1 _16057_ ( .A1(_05155_ ), .A2(_07130_ ), .ZN(_08040_ ) );
AND3_X1 _16058_ ( .A1(_05153_ ), .A2(_02425_ ), .A3(_07368_ ), .ZN(_08041_ ) );
NOR3_X1 _16059_ ( .A1(_08039_ ), .A2(_08040_ ), .A3(_08041_ ), .ZN(_08042_ ) );
NAND3_X1 _16060_ ( .A1(_08034_ ), .A2(_08038_ ), .A3(_08042_ ), .ZN(_08043_ ) );
AOI21_X1 _16061_ ( .A(_08017_ ), .B1(_08043_ ), .B2(_07756_ ), .ZN(_08044_ ) );
OAI21_X1 _16062_ ( .A(_08006_ ), .B1(_05571_ ), .B2(_07788_ ), .ZN(_08045_ ) );
OAI21_X1 _16063_ ( .A(_08009_ ), .B1(_08044_ ), .B2(_08045_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
NAND2_X1 _16064_ ( .A1(_06066_ ), .A2(_08008_ ), .ZN(_08046_ ) );
NOR2_X1 _16065_ ( .A1(_05115_ ), .A2(_05118_ ), .ZN(_08047_ ) );
NOR3_X1 _16066_ ( .A1(_05119_ ), .A2(_08047_ ), .A3(_07207_ ), .ZN(_08048_ ) );
AND2_X1 _16067_ ( .A1(_06053_ ), .A2(_07084_ ), .ZN(_08049_ ) );
AND3_X1 _16068_ ( .A1(_06797_ ), .A2(\ID_EX_imm [1] ), .A3(_06785_ ), .ZN(_08050_ ) );
NOR3_X1 _16069_ ( .A1(_08048_ ), .A2(_08049_ ), .A3(_08050_ ), .ZN(_08051_ ) );
OAI21_X1 _16070_ ( .A(_06141_ ), .B1(_08051_ ), .B2(_06803_ ), .ZN(_08052_ ) );
OR2_X1 _16071_ ( .A1(_07366_ ), .A2(_06986_ ), .ZN(_08053_ ) );
OAI21_X1 _16072_ ( .A(_07033_ ), .B1(_07056_ ), .B2(_07047_ ), .ZN(_08054_ ) );
OAI211_X1 _16073_ ( .A(_08054_ ), .B(_07005_ ), .C1(_07954_ ), .C2(_07142_ ), .ZN(_08055_ ) );
OAI211_X1 _16074_ ( .A(_08055_ ), .B(_07009_ ), .C1(_07024_ ), .C2(_07901_ ), .ZN(_08056_ ) );
AND2_X1 _16075_ ( .A1(_07766_ ), .A2(_07762_ ), .ZN(_08057_ ) );
OAI211_X1 _16076_ ( .A(_06995_ ), .B(_08056_ ), .C1(_08057_ ), .C2(_07315_ ), .ZN(_08058_ ) );
AOI21_X1 _16077_ ( .A(_07557_ ), .B1(_08053_ ), .B2(_08058_ ), .ZN(_08059_ ) );
NAND4_X1 _16078_ ( .A1(_07287_ ), .A2(_06942_ ), .A3(_06935_ ), .A4(_07501_ ), .ZN(_08060_ ) );
NAND3_X1 _16079_ ( .A1(_08060_ ), .A2(_08058_ ), .A3(_08053_ ), .ZN(_08061_ ) );
AOI221_X4 _16080_ ( .A(_08059_ ), .B1(_07375_ ), .B2(_07480_ ), .C1(_08061_ ), .C2(_06882_ ), .ZN(_08062_ ) );
OAI21_X1 _16081_ ( .A(_06878_ ), .B1(_05239_ ), .B2(_06806_ ), .ZN(_08063_ ) );
OR2_X1 _16082_ ( .A1(_08063_ ), .A2(_06810_ ), .ZN(_08064_ ) );
NOR3_X1 _16083_ ( .A1(_06808_ ), .A2(_06809_ ), .A3(_05468_ ), .ZN(_08065_ ) );
NOR3_X1 _16084_ ( .A1(_02862_ ), .A2(_07142_ ), .A3(_07190_ ), .ZN(_08066_ ) );
AOI21_X1 _16085_ ( .A(_07130_ ), .B1(_02862_ ), .B2(_07142_ ), .ZN(_08067_ ) );
NOR3_X1 _16086_ ( .A1(_08065_ ), .A2(_08066_ ), .A3(_08067_ ), .ZN(_08068_ ) );
NAND3_X1 _16087_ ( .A1(_08062_ ), .A2(_08064_ ), .A3(_08068_ ), .ZN(_08069_ ) );
AOI21_X1 _16088_ ( .A(_08052_ ), .B1(_08069_ ), .B2(_07756_ ), .ZN(_08070_ ) );
OAI21_X1 _16089_ ( .A(_08006_ ), .B1(_05620_ ), .B2(\ID_EX_pc [1] ), .ZN(_08071_ ) );
OAI21_X1 _16090_ ( .A(_08046_ ), .B1(_08070_ ), .B2(_08071_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
OR2_X1 _16091_ ( .A1(_06097_ ), .A2(_06491_ ), .ZN(_08072_ ) );
AND2_X1 _16092_ ( .A1(_04291_ ), .A2(\ID_EX_typ [2] ), .ZN(_08073_ ) );
OAI21_X1 _16093_ ( .A(_08073_ ), .B1(_05386_ ), .B2(_05136_ ), .ZN(_08074_ ) );
AOI211_X1 _16094_ ( .A(_08074_ ), .B(_05385_ ), .C1(_05149_ ), .C2(_05390_ ), .ZN(_08075_ ) );
AND2_X1 _16095_ ( .A1(_05383_ ), .A2(_08075_ ), .ZN(_08076_ ) );
NAND4_X1 _16096_ ( .A1(_06933_ ), .A2(_05212_ ), .A3(_06882_ ), .A4(_06927_ ), .ZN(_00340_ ) );
AOI211_X1 _16097_ ( .A(_06986_ ), .B(_07405_ ), .C1(_07407_ ), .C2(_06984_ ), .ZN(_00341_ ) );
AOI211_X1 _16098_ ( .A(_07008_ ), .B(_07794_ ), .C1(_07140_ ), .C2(_07585_ ), .ZN(_00342_ ) );
NOR2_X1 _16099_ ( .A1(_07931_ ), .A2(_06951_ ), .ZN(_00343_ ) );
OAI21_X1 _16100_ ( .A(_07025_ ), .B1(_07132_ ), .B2(_07136_ ), .ZN(_00344_ ) );
AOI21_X1 _16101_ ( .A(_05116_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_00345_ ) );
OAI21_X1 _16102_ ( .A(_07137_ ), .B1(_07135_ ), .B2(_00345_ ), .ZN(_00346_ ) );
AND3_X1 _16103_ ( .A1(_00344_ ), .A2(_00346_ ), .A3(_07004_ ), .ZN(_00347_ ) );
NOR3_X1 _16104_ ( .A1(_00343_ ), .A2(_06983_ ), .A3(_00347_ ), .ZN(_00348_ ) );
NOR3_X1 _16105_ ( .A1(_00342_ ), .A2(_00348_ ), .A3(_07060_ ), .ZN(_00349_ ) );
NOR2_X1 _16106_ ( .A1(_00341_ ), .A2(_00349_ ), .ZN(_00350_ ) );
AOI21_X1 _16107_ ( .A(_07461_ ), .B1(_00340_ ), .B2(_00350_ ), .ZN(_00351_ ) );
AND3_X1 _16108_ ( .A1(_06888_ ), .A2(_05116_ ), .A3(_07479_ ), .ZN(_00352_ ) );
OR3_X1 _16109_ ( .A1(_08076_ ), .A2(_00351_ ), .A3(_00352_ ), .ZN(_00353_ ) );
NOR3_X1 _16110_ ( .A1(_06806_ ), .A2(_00345_ ), .A3(_06879_ ), .ZN(_00354_ ) );
OAI21_X1 _16111_ ( .A(_07068_ ), .B1(_07806_ ), .B2(_05243_ ), .ZN(_00355_ ) );
OAI221_X1 _16112_ ( .A(_00355_ ), .B1(_07129_ ), .B2(_00345_ ), .C1(_07190_ ), .C2(_06807_ ), .ZN(_00356_ ) );
NOR3_X1 _16113_ ( .A1(_00353_ ), .A2(_00354_ ), .A3(_00356_ ), .ZN(_00357_ ) );
OAI21_X1 _16114_ ( .A(_06141_ ), .B1(_00357_ ), .B2(_07076_ ), .ZN(_00358_ ) );
AND3_X1 _16115_ ( .A1(_05123_ ), .A2(_07073_ ), .A3(_05144_ ), .ZN(_00359_ ) );
AND4_X1 _16116_ ( .A1(\ID_EX_typ [4] ), .A2(_04291_ ), .A3(\ID_EX_typ [3] ), .A4(_05127_ ), .ZN(_00360_ ) );
OAI21_X1 _16117_ ( .A(_05392_ ), .B1(_00359_ ), .B2(_00360_ ), .ZN(_00361_ ) );
AND3_X1 _16118_ ( .A1(_06797_ ), .A2(\ID_EX_imm [0] ), .A3(_06785_ ), .ZN(_00362_ ) );
AOI21_X1 _16119_ ( .A(_00362_ ), .B1(_06099_ ), .B2(_07084_ ), .ZN(_00363_ ) );
OAI21_X1 _16120_ ( .A(_07445_ ), .B1(_04977_ ), .B2(_05117_ ), .ZN(_00364_ ) );
NAND3_X1 _16121_ ( .A1(_00361_ ), .A2(_00363_ ), .A3(_00364_ ), .ZN(_00365_ ) );
AOI21_X1 _16122_ ( .A(_00358_ ), .B1(_07816_ ), .B2(_00365_ ), .ZN(_00366_ ) );
OAI21_X1 _16123_ ( .A(_08006_ ), .B1(_05480_ ), .B2(\ID_EX_pc [0] ), .ZN(_00367_ ) );
OAI21_X1 _16124_ ( .A(_08072_ ), .B1(_00366_ ), .B2(_00367_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
NAND2_X1 _16125_ ( .A1(_05874_ ), .A2(_08008_ ), .ZN(_00368_ ) );
NOR2_X1 _16126_ ( .A1(_05868_ ), .A2(_06788_ ), .ZN(_00369_ ) );
OAI21_X1 _16127_ ( .A(_06795_ ), .B1(_07615_ ), .B2(_07616_ ), .ZN(_00370_ ) );
AOI21_X1 _16128_ ( .A(_00370_ ), .B1(_07616_ ), .B2(_07615_ ), .ZN(_00371_ ) );
AND3_X1 _16129_ ( .A1(_06797_ ), .A2(\ID_EX_imm [28] ), .A3(_06785_ ), .ZN(_00372_ ) );
NOR3_X1 _16130_ ( .A1(_00369_ ), .A2(_00371_ ), .A3(_00372_ ), .ZN(_00373_ ) );
OAI21_X1 _16131_ ( .A(_06141_ ), .B1(_00373_ ), .B2(_06803_ ), .ZN(_00374_ ) );
AND3_X1 _16132_ ( .A1(_06926_ ), .A2(_06934_ ), .A3(_07099_ ), .ZN(_00375_ ) );
OAI21_X1 _16133_ ( .A(_00375_ ), .B1(_06929_ ), .B2(_06931_ ), .ZN(_00376_ ) );
NAND3_X1 _16134_ ( .A1(_07124_ ), .A2(_07010_ ), .A3(_07006_ ), .ZN(_00377_ ) );
OAI211_X1 _16135_ ( .A(_07654_ ), .B(_00376_ ), .C1(_07061_ ), .C2(_00377_ ), .ZN(_00378_ ) );
NAND2_X1 _16136_ ( .A1(_00378_ ), .A2(_06883_ ), .ZN(_00379_ ) );
MUX2_X1 _16137_ ( .A(_07667_ ), .B(_07663_ ), .S(_07137_ ), .Z(_00380_ ) );
OR2_X1 _16138_ ( .A1(_00380_ ), .A2(_06944_ ), .ZN(_00381_ ) );
OAI21_X1 _16139_ ( .A(_07141_ ), .B1(_07102_ ), .B2(_07115_ ), .ZN(_00382_ ) );
OAI21_X1 _16140_ ( .A(_07181_ ), .B1(_07114_ ), .B2(_07112_ ), .ZN(_00383_ ) );
AND2_X1 _16141_ ( .A1(_00382_ ), .A2(_00383_ ), .ZN(_00384_ ) );
OAI21_X1 _16142_ ( .A(_00381_ ), .B1(_00384_ ), .B2(_07024_ ), .ZN(_00385_ ) );
MUX2_X1 _16143_ ( .A(_07186_ ), .B(_00385_ ), .S(_07315_ ), .Z(_00386_ ) );
AOI21_X1 _16144_ ( .A(_07045_ ), .B1(_00386_ ), .B2(_06996_ ), .ZN(_00387_ ) );
OAI21_X1 _16145_ ( .A(_00387_ ), .B1(_07234_ ), .B2(_07599_ ), .ZN(_00388_ ) );
OR3_X1 _16146_ ( .A1(_00377_ ), .A2(_07146_ ), .A3(_07557_ ), .ZN(_00389_ ) );
NAND3_X1 _16147_ ( .A1(_00379_ ), .A2(_00388_ ), .A3(_00389_ ), .ZN(_00390_ ) );
OAI21_X1 _16148_ ( .A(_06878_ ), .B1(_07644_ ), .B2(_07645_ ), .ZN(_00391_ ) );
AOI21_X1 _16149_ ( .A(_00391_ ), .B1(_07645_ ), .B2(_07644_ ), .ZN(_00392_ ) );
NAND2_X1 _16150_ ( .A1(_05161_ ), .A2(_07192_ ), .ZN(_00393_ ) );
NAND3_X1 _16151_ ( .A1(_05159_ ), .A2(_02448_ ), .A3(_07368_ ), .ZN(_00394_ ) );
OAI21_X1 _16152_ ( .A(_05129_ ), .B1(_05159_ ), .B2(_02448_ ), .ZN(_00395_ ) );
NAND3_X1 _16153_ ( .A1(_00393_ ), .A2(_00394_ ), .A3(_00395_ ), .ZN(_00396_ ) );
OR3_X1 _16154_ ( .A1(_00390_ ), .A2(_00392_ ), .A3(_00396_ ), .ZN(_00397_ ) );
AOI21_X1 _16155_ ( .A(_00374_ ), .B1(_00397_ ), .B2(_07756_ ), .ZN(_00398_ ) );
OAI21_X1 _16156_ ( .A(_08006_ ), .B1(_05840_ ), .B2(_07788_ ), .ZN(_00399_ ) );
OAI21_X1 _16157_ ( .A(_00368_ ), .B1(_00398_ ), .B2(_00399_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _16158_ ( .A1(_06085_ ), .A2(_08008_ ), .ZN(_00400_ ) );
OAI22_X1 _16159_ ( .A1(_06076_ ), .A2(_06788_ ), .B1(_02488_ ), .B2(_07945_ ), .ZN(_00401_ ) );
AND2_X1 _16160_ ( .A1(_07614_ ), .A2(_04701_ ), .ZN(_00402_ ) );
OR3_X1 _16161_ ( .A1(_00402_ ), .A2(_04723_ ), .A3(_05453_ ), .ZN(_00403_ ) );
OAI21_X1 _16162_ ( .A(_04723_ ), .B1(_00402_ ), .B2(_05453_ ), .ZN(_00404_ ) );
AND3_X1 _16163_ ( .A1(_00403_ ), .A2(_06795_ ), .A3(_00404_ ), .ZN(_00405_ ) );
OAI21_X1 _16164_ ( .A(_07816_ ), .B1(_00401_ ), .B2(_00405_ ), .ZN(_00406_ ) );
NAND2_X1 _16165_ ( .A1(_00406_ ), .A2(_05601_ ), .ZN(_00407_ ) );
NAND2_X1 _16166_ ( .A1(_08023_ ), .A2(_07181_ ), .ZN(_00408_ ) );
OAI211_X1 _16167_ ( .A(_07224_ ), .B(_06939_ ), .C1(_03207_ ), .C2(_06941_ ), .ZN(_00409_ ) );
NAND2_X1 _16168_ ( .A1(_00408_ ), .A2(_00409_ ), .ZN(_00410_ ) );
NOR3_X1 _16169_ ( .A1(_06966_ ), .A2(_07181_ ), .A3(_06971_ ), .ZN(_00411_ ) );
NOR3_X1 _16170_ ( .A1(_07034_ ), .A2(_06967_ ), .A3(_06939_ ), .ZN(_00412_ ) );
OR2_X1 _16171_ ( .A1(_00411_ ), .A2(_00412_ ), .ZN(_00413_ ) );
MUX2_X1 _16172_ ( .A(_00410_ ), .B(_00413_ ), .S(_07255_ ), .Z(_00414_ ) );
OAI21_X1 _16173_ ( .A(_07480_ ), .B1(_00414_ ), .B2(_07257_ ), .ZN(_00415_ ) );
AND2_X1 _16174_ ( .A1(_07256_ ), .A2(_07257_ ), .ZN(_00416_ ) );
NOR2_X1 _16175_ ( .A1(_00415_ ), .A2(_00416_ ), .ZN(_00417_ ) );
INV_X1 _16176_ ( .A(_07213_ ), .ZN(_00418_ ) );
INV_X1 _16177_ ( .A(_07653_ ), .ZN(_00419_ ) );
OAI211_X1 _16178_ ( .A(_06933_ ), .B(_07214_ ), .C1(_06928_ ), .C2(_06931_ ), .ZN(_00420_ ) );
NAND2_X1 _16179_ ( .A1(_07704_ ), .A2(_06995_ ), .ZN(_00421_ ) );
NAND4_X1 _16180_ ( .A1(_00418_ ), .A2(_00419_ ), .A3(_00420_ ), .A4(_00421_ ), .ZN(_00422_ ) );
NAND2_X1 _16181_ ( .A1(_00422_ ), .A2(_06882_ ), .ZN(_00423_ ) );
OAI21_X1 _16182_ ( .A(_00423_ ), .B1(_07557_ ), .B2(_00421_ ), .ZN(_00424_ ) );
NAND2_X1 _16183_ ( .A1(_07715_ ), .A2(_07716_ ), .ZN(_00425_ ) );
NOR2_X1 _16184_ ( .A1(_05217_ ), .A2(_07045_ ), .ZN(_00426_ ) );
AOI211_X1 _16185_ ( .A(_00417_ ), .B(_00424_ ), .C1(_00425_ ), .C2(_00426_ ), .ZN(_00427_ ) );
INV_X1 _16186_ ( .A(_05354_ ), .ZN(_00428_ ) );
OAI211_X1 _16187_ ( .A(_05366_ ), .B(_05371_ ), .C1(_07626_ ), .C2(_07636_ ), .ZN(_00429_ ) );
AOI21_X1 _16188_ ( .A(_00428_ ), .B1(_00429_ ), .B2(_07641_ ), .ZN(_00430_ ) );
OR3_X1 _16189_ ( .A1(_00430_ ), .A2(_05358_ ), .A3(_05352_ ), .ZN(_00431_ ) );
OAI21_X1 _16190_ ( .A(_05358_ ), .B1(_00430_ ), .B2(_05352_ ), .ZN(_00432_ ) );
NAND3_X1 _16191_ ( .A1(_00431_ ), .A2(_07246_ ), .A3(_00432_ ), .ZN(_00433_ ) );
AND2_X1 _16192_ ( .A1(_05358_ ), .A2(_07192_ ), .ZN(_00434_ ) );
NOR3_X1 _16193_ ( .A1(_05455_ ), .A2(_05357_ ), .A3(_07190_ ), .ZN(_00435_ ) );
AOI21_X1 _16194_ ( .A(_07130_ ), .B1(_05455_ ), .B2(_05357_ ), .ZN(_00436_ ) );
NOR3_X1 _16195_ ( .A1(_00434_ ), .A2(_00435_ ), .A3(_00436_ ), .ZN(_00437_ ) );
NAND3_X1 _16196_ ( .A1(_00427_ ), .A2(_00433_ ), .A3(_00437_ ), .ZN(_00438_ ) );
AOI21_X1 _16197_ ( .A(_00407_ ), .B1(_00438_ ), .B2(_07756_ ), .ZN(_00439_ ) );
OAI21_X1 _16198_ ( .A(_08006_ ), .B1(_06071_ ), .B2(_07788_ ), .ZN(_00440_ ) );
OAI21_X1 _16199_ ( .A(_00400_ ), .B1(_00439_ ), .B2(_00440_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
NAND2_X1 _16200_ ( .A1(_06114_ ), .A2(_08008_ ), .ZN(_00441_ ) );
OAI22_X1 _16201_ ( .A1(_06106_ ), .A2(_06788_ ), .B1(_03208_ ), .B2(_07945_ ), .ZN(_00442_ ) );
NOR2_X1 _16202_ ( .A1(_07614_ ), .A2(_04701_ ), .ZN(_00443_ ) );
NOR3_X1 _16203_ ( .A1(_00402_ ), .A2(_00443_ ), .A3(_07207_ ), .ZN(_00444_ ) );
OAI21_X1 _16204_ ( .A(_07816_ ), .B1(_00442_ ), .B2(_00444_ ), .ZN(_00445_ ) );
NAND2_X1 _16205_ ( .A1(_00445_ ), .A2(_05601_ ), .ZN(_00446_ ) );
NOR2_X1 _16206_ ( .A1(_07303_ ), .A2(_06984_ ), .ZN(_00447_ ) );
AND2_X1 _16207_ ( .A1(_00447_ ), .A2(_06986_ ), .ZN(_00448_ ) );
OR3_X1 _16208_ ( .A1(_07213_ ), .A2(_07653_ ), .A3(_00448_ ), .ZN(_00449_ ) );
NOR3_X1 _16209_ ( .A1(_06932_ ), .A2(_07288_ ), .A3(_07289_ ), .ZN(_00450_ ) );
OAI21_X1 _16210_ ( .A(_06883_ ), .B1(_00449_ ), .B2(_00450_ ), .ZN(_00451_ ) );
NAND3_X1 _16211_ ( .A1(_00447_ ), .A2(_06988_ ), .A3(_06993_ ), .ZN(_00452_ ) );
AND3_X1 _16212_ ( .A1(_07668_ ), .A2(_07669_ ), .A3(_07006_ ), .ZN(_00453_ ) );
AOI21_X1 _16213_ ( .A(_07006_ ), .B1(_07672_ ), .B2(_07673_ ), .ZN(_00454_ ) );
OAI21_X1 _16214_ ( .A(_07055_ ), .B1(_00453_ ), .B2(_00454_ ), .ZN(_00455_ ) );
NAND2_X1 _16215_ ( .A1(_07325_ ), .A2(_07257_ ), .ZN(_00456_ ) );
NAND3_X1 _16216_ ( .A1(_00455_ ), .A2(_07480_ ), .A3(_00456_ ), .ZN(_00457_ ) );
NAND3_X1 _16217_ ( .A1(_07742_ ), .A2(_07743_ ), .A3(_00426_ ), .ZN(_00458_ ) );
AND4_X1 _16218_ ( .A1(_00451_ ), .A2(_00452_ ), .A3(_00457_ ), .A4(_00458_ ), .ZN(_00459_ ) );
AND3_X1 _16219_ ( .A1(_00429_ ), .A2(_00428_ ), .A3(_07641_ ), .ZN(_00460_ ) );
OR3_X1 _16220_ ( .A1(_00460_ ), .A2(_00430_ ), .A3(_06880_ ), .ZN(_00461_ ) );
OR3_X1 _16221_ ( .A1(_05352_ ), .A2(_05353_ ), .A3(_05468_ ), .ZN(_00462_ ) );
OR3_X1 _16222_ ( .A1(_05350_ ), .A2(_05351_ ), .A3(_07065_ ), .ZN(_00463_ ) );
OR2_X1 _16223_ ( .A1(_05353_ ), .A2(_07129_ ), .ZN(_00464_ ) );
AND3_X1 _16224_ ( .A1(_00462_ ), .A2(_00463_ ), .A3(_00464_ ), .ZN(_00465_ ) );
NAND3_X1 _16225_ ( .A1(_00459_ ), .A2(_00461_ ), .A3(_00465_ ), .ZN(_00466_ ) );
AOI21_X1 _16226_ ( .A(_00446_ ), .B1(_00466_ ), .B2(_07756_ ), .ZN(_00467_ ) );
OAI21_X1 _16227_ ( .A(_08006_ ), .B1(_06103_ ), .B2(_07788_ ), .ZN(_00468_ ) );
OAI21_X1 _16228_ ( .A(_00441_ ), .B1(_00467_ ), .B2(_00468_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _16229_ ( .A1(_06137_ ), .A2(_08008_ ), .ZN(_00469_ ) );
OAI22_X1 _16230_ ( .A1(_06129_ ), .A2(_06788_ ), .B1(_03210_ ), .B2(_07945_ ), .ZN(_00470_ ) );
AND2_X1 _16231_ ( .A1(_07612_ ), .A2(_04654_ ), .ZN(_00471_ ) );
OR3_X1 _16232_ ( .A1(_00471_ ), .A2(_04677_ ), .A3(_05458_ ), .ZN(_00472_ ) );
OAI21_X1 _16233_ ( .A(_04677_ ), .B1(_00471_ ), .B2(_05458_ ), .ZN(_00473_ ) );
AND3_X1 _16234_ ( .A1(_00472_ ), .A2(_06795_ ), .A3(_00473_ ), .ZN(_00474_ ) );
OAI21_X1 _16235_ ( .A(_07816_ ), .B1(_00470_ ), .B2(_00474_ ), .ZN(_00475_ ) );
NAND2_X1 _16236_ ( .A1(_00475_ ), .A2(_05601_ ), .ZN(_00476_ ) );
AND3_X1 _16237_ ( .A1(_07362_ ), .A2(_07054_ ), .A3(_07364_ ), .ZN(_00477_ ) );
NAND2_X1 _16238_ ( .A1(_00477_ ), .A2(_06987_ ), .ZN(_00478_ ) );
NAND3_X1 _16239_ ( .A1(_00418_ ), .A2(_00419_ ), .A3(_00478_ ), .ZN(_00479_ ) );
NAND3_X1 _16240_ ( .A1(_07287_ ), .A2(_06942_ ), .A3(_06934_ ), .ZN(_00480_ ) );
NOR2_X1 _16241_ ( .A1(_00480_ ), .A2(_06932_ ), .ZN(_00481_ ) );
OAI21_X1 _16242_ ( .A(_06883_ ), .B1(_00479_ ), .B2(_00481_ ), .ZN(_00482_ ) );
NAND3_X1 _16243_ ( .A1(_00477_ ), .A2(_06988_ ), .A3(_06993_ ), .ZN(_00483_ ) );
NAND2_X1 _16244_ ( .A1(_05371_ ), .A2(_07192_ ), .ZN(_00484_ ) );
OAI21_X1 _16245_ ( .A(_05129_ ), .B1(_07639_ ), .B2(_03184_ ), .ZN(_00485_ ) );
AND4_X1 _16246_ ( .A1(_00482_ ), .A2(_00483_ ), .A3(_00484_ ), .A4(_00485_ ), .ZN(_00486_ ) );
NOR2_X1 _16247_ ( .A1(_07626_ ), .A2(_07636_ ), .ZN(_00487_ ) );
NOR2_X1 _16248_ ( .A1(_00487_ ), .A2(_05367_ ), .ZN(_00488_ ) );
OR3_X1 _16249_ ( .A1(_00488_ ), .A2(_05364_ ), .A3(_05371_ ), .ZN(_00489_ ) );
OAI21_X1 _16250_ ( .A(_05371_ ), .B1(_00488_ ), .B2(_05364_ ), .ZN(_00490_ ) );
NAND3_X1 _16251_ ( .A1(_00489_ ), .A2(_06878_ ), .A3(_00490_ ), .ZN(_00491_ ) );
AOI211_X1 _16252_ ( .A(_06996_ ), .B(_07045_ ), .C1(_07772_ ), .C2(_07773_ ), .ZN(_00492_ ) );
NOR2_X1 _16253_ ( .A1(_08024_ ), .A2(_07255_ ), .ZN(_00493_ ) );
AOI21_X1 _16254_ ( .A(_07006_ ), .B1(_07035_ ), .B2(_07039_ ), .ZN(_00494_ ) );
OAI21_X1 _16255_ ( .A(_07055_ ), .B1(_00493_ ), .B2(_00494_ ), .ZN(_00495_ ) );
NAND2_X1 _16256_ ( .A1(_00495_ ), .A2(_07480_ ), .ZN(_00496_ ) );
AOI21_X1 _16257_ ( .A(_00496_ ), .B1(_07257_ ), .B2(_07382_ ), .ZN(_00497_ ) );
AOI211_X1 _16258_ ( .A(_00492_ ), .B(_00497_ ), .C1(_07640_ ), .C2(_07368_ ), .ZN(_00498_ ) );
NAND3_X1 _16259_ ( .A1(_00486_ ), .A2(_00491_ ), .A3(_00498_ ), .ZN(_00499_ ) );
AOI21_X1 _16260_ ( .A(_00476_ ), .B1(_00499_ ), .B2(_07077_ ), .ZN(_00500_ ) );
OAI21_X1 _16261_ ( .A(_08006_ ), .B1(_06124_ ), .B2(_07788_ ), .ZN(_00501_ ) );
OAI21_X1 _16262_ ( .A(_00469_ ), .B1(_00500_ ), .B2(_00501_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _16263_ ( .A1(_06156_ ), .A2(_08008_ ), .ZN(_00502_ ) );
OAI22_X1 _16264_ ( .A1(_06147_ ), .A2(_06788_ ), .B1(_02511_ ), .B2(_07945_ ), .ZN(_00503_ ) );
NOR2_X1 _16265_ ( .A1(_07612_ ), .A2(_04654_ ), .ZN(_00504_ ) );
NOR3_X1 _16266_ ( .A1(_00471_ ), .A2(_00504_ ), .A3(_07207_ ), .ZN(_00505_ ) );
OAI21_X1 _16267_ ( .A(_07816_ ), .B1(_00503_ ), .B2(_00505_ ), .ZN(_00506_ ) );
NAND2_X1 _16268_ ( .A1(_00506_ ), .A2(_05601_ ), .ZN(_00507_ ) );
INV_X1 _16269_ ( .A(_06887_ ), .ZN(_00508_ ) );
AOI211_X1 _16270_ ( .A(_07097_ ), .B(_07398_ ), .C1(_07055_ ), .C2(_00508_ ), .ZN(_00509_ ) );
NOR2_X1 _16271_ ( .A1(_07407_ ), .A2(_07415_ ), .ZN(_00510_ ) );
AOI211_X1 _16272_ ( .A(_00509_ ), .B(_07213_ ), .C1(_07234_ ), .C2(_00510_ ), .ZN(_00511_ ) );
NOR2_X1 _16273_ ( .A1(_00511_ ), .A2(_07544_ ), .ZN(_00512_ ) );
OAI21_X1 _16274_ ( .A(_06878_ ), .B1(_00487_ ), .B2(_05367_ ), .ZN(_00513_ ) );
AOI21_X1 _16275_ ( .A(_00513_ ), .B1(_05367_ ), .B2(_00487_ ), .ZN(_00514_ ) );
NAND2_X1 _16276_ ( .A1(_07805_ ), .A2(_07807_ ), .ZN(_00515_ ) );
NAND2_X1 _16277_ ( .A1(_00515_ ), .A2(_00426_ ), .ZN(_00516_ ) );
OR3_X1 _16278_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_05468_ ), .ZN(_00517_ ) );
OR3_X1 _16279_ ( .A1(_05362_ ), .A2(_05363_ ), .A3(_07065_ ), .ZN(_00518_ ) );
OR2_X1 _16280_ ( .A1(_05365_ ), .A2(_05130_ ), .ZN(_00519_ ) );
AND4_X1 _16281_ ( .A1(_00516_ ), .A2(_00517_ ), .A3(_00518_ ), .A4(_00519_ ), .ZN(_00520_ ) );
NAND3_X1 _16282_ ( .A1(_00382_ ), .A2(_00383_ ), .A3(_07024_ ), .ZN(_00521_ ) );
NAND3_X1 _16283_ ( .A1(_07180_ ), .A2(_07184_ ), .A3(_06981_ ), .ZN(_00522_ ) );
AND3_X1 _16284_ ( .A1(_00521_ ), .A2(_00522_ ), .A3(_07315_ ), .ZN(_00523_ ) );
AOI21_X1 _16285_ ( .A(_07315_ ), .B1(_07417_ ), .B2(_07418_ ), .ZN(_00524_ ) );
OR3_X1 _16286_ ( .A1(_00523_ ), .A2(_00524_ ), .A3(_07559_ ), .ZN(_00525_ ) );
NAND3_X1 _16287_ ( .A1(_00510_ ), .A2(_07234_ ), .A3(_06992_ ), .ZN(_00526_ ) );
NAND3_X1 _16288_ ( .A1(_00520_ ), .A2(_00525_ ), .A3(_00526_ ), .ZN(_00527_ ) );
OR3_X1 _16289_ ( .A1(_00512_ ), .A2(_00514_ ), .A3(_00527_ ), .ZN(_00528_ ) );
AOI21_X1 _16290_ ( .A(_00507_ ), .B1(_00528_ ), .B2(_07077_ ), .ZN(_00529_ ) );
OAI21_X1 _16291_ ( .A(_08006_ ), .B1(_06144_ ), .B2(_07788_ ), .ZN(_00530_ ) );
OAI21_X1 _16292_ ( .A(_00502_ ), .B1(_00529_ ), .B2(_00530_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _16293_ ( .A1(_06175_ ), .A2(_08008_ ), .ZN(_00531_ ) );
NAND3_X1 _16294_ ( .A1(_06791_ ), .A2(_04504_ ), .A3(_04529_ ), .ZN(_00532_ ) );
OAI21_X1 _16295_ ( .A(_00532_ ), .B1(_04528_ ), .B2(_05440_ ), .ZN(_00533_ ) );
AND2_X1 _16296_ ( .A1(_00533_ ), .A2(_04456_ ), .ZN(_00534_ ) );
OR3_X1 _16297_ ( .A1(_00534_ ), .A2(_04481_ ), .A3(_05436_ ), .ZN(_00535_ ) );
OAI21_X1 _16298_ ( .A(_04481_ ), .B1(_00534_ ), .B2(_05436_ ), .ZN(_00536_ ) );
AND3_X1 _16299_ ( .A1(_00535_ ), .A2(_06795_ ), .A3(_00536_ ), .ZN(_00537_ ) );
OAI22_X1 _16300_ ( .A1(_06167_ ), .A2(_06788_ ), .B1(_02562_ ), .B2(_07945_ ), .ZN(_00538_ ) );
OAI21_X1 _16301_ ( .A(_07816_ ), .B1(_00537_ ), .B2(_00538_ ), .ZN(_00539_ ) );
NAND2_X1 _16302_ ( .A1(_00539_ ), .A2(_06141_ ), .ZN(_00540_ ) );
NAND3_X1 _16303_ ( .A1(_06869_ ), .A2(_05302_ ), .A3(_05314_ ), .ZN(_00541_ ) );
INV_X1 _16304_ ( .A(_07630_ ), .ZN(_00542_ ) );
AOI21_X1 _16305_ ( .A(_05298_ ), .B1(_00541_ ), .B2(_00542_ ), .ZN(_00543_ ) );
INV_X1 _16306_ ( .A(_00543_ ), .ZN(_00544_ ) );
INV_X1 _16307_ ( .A(_07634_ ), .ZN(_00545_ ) );
AOI21_X1 _16308_ ( .A(_05328_ ), .B1(_00544_ ), .B2(_00545_ ), .ZN(_00546_ ) );
NOR3_X1 _16309_ ( .A1(_00543_ ), .A2(_05329_ ), .A3(_07634_ ), .ZN(_00547_ ) );
OAI21_X1 _16310_ ( .A(_07246_ ), .B1(_00546_ ), .B2(_00547_ ), .ZN(_00548_ ) );
OAI22_X1 _16311_ ( .A1(_07628_ ), .A2(_07190_ ), .B1(_05309_ ), .B2(_07130_ ), .ZN(_00549_ ) );
AOI21_X1 _16312_ ( .A(_00549_ ), .B1(_05328_ ), .B2(_07192_ ), .ZN(_00550_ ) );
NAND2_X1 _16313_ ( .A1(_07839_ ), .A2(_07840_ ), .ZN(_00551_ ) );
NAND2_X1 _16314_ ( .A1(_00551_ ), .A2(_07234_ ), .ZN(_00552_ ) );
AOI21_X1 _16315_ ( .A(_07544_ ), .B1(_07654_ ), .B2(_00552_ ), .ZN(_00553_ ) );
OR3_X1 _16316_ ( .A1(_07474_ ), .A2(_06987_ ), .A3(_07415_ ), .ZN(_00554_ ) );
NAND3_X1 _16317_ ( .A1(_07476_ ), .A2(_07477_ ), .A3(_07415_ ), .ZN(_00555_ ) );
NOR3_X1 _16318_ ( .A1(_00411_ ), .A2(_00412_ ), .A3(_06965_ ), .ZN(_00556_ ) );
AOI21_X1 _16319_ ( .A(_06951_ ), .B1(_07249_ ), .B2(_07250_ ), .ZN(_00557_ ) );
NOR2_X1 _16320_ ( .A1(_00556_ ), .A2(_00557_ ), .ZN(_00558_ ) );
OAI211_X1 _16321_ ( .A(_07234_ ), .B(_00555_ ), .C1(_00558_ ), .C2(_07257_ ), .ZN(_00559_ ) );
AOI21_X1 _16322_ ( .A(_07045_ ), .B1(_00554_ ), .B2(_00559_ ), .ZN(_00560_ ) );
AND3_X1 _16323_ ( .A1(_00551_ ), .A2(_07234_ ), .A3(_06992_ ), .ZN(_00561_ ) );
NOR3_X1 _16324_ ( .A1(_00553_ ), .A2(_00560_ ), .A3(_00561_ ), .ZN(_00562_ ) );
NAND3_X1 _16325_ ( .A1(_00548_ ), .A2(_00550_ ), .A3(_00562_ ), .ZN(_00563_ ) );
AOI21_X1 _16326_ ( .A(_00540_ ), .B1(_00563_ ), .B2(_07077_ ), .ZN(_00564_ ) );
OAI21_X1 _16327_ ( .A(_08006_ ), .B1(_06161_ ), .B2(_07788_ ), .ZN(_00565_ ) );
OAI21_X1 _16328_ ( .A(_00531_ ), .B1(_00564_ ), .B2(_00565_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _16329_ ( .A1(_06186_ ), .A2(_08008_ ), .ZN(_00566_ ) );
NOR2_X1 _16330_ ( .A1(_00533_ ), .A2(_04456_ ), .ZN(_00567_ ) );
NOR3_X1 _16331_ ( .A1(_00534_ ), .A2(_00567_ ), .A3(_07207_ ), .ZN(_00568_ ) );
NOR3_X1 _16332_ ( .A1(_06189_ ), .A2(_06165_ ), .A3(_06787_ ), .ZN(_00569_ ) );
AND3_X1 _16333_ ( .A1(_06797_ ), .A2(\ID_EX_imm [22] ), .A3(_06785_ ), .ZN(_00570_ ) );
NOR3_X1 _16334_ ( .A1(_00568_ ), .A2(_00569_ ), .A3(_00570_ ), .ZN(_00571_ ) );
OAI21_X1 _16335_ ( .A(_06141_ ), .B1(_00571_ ), .B2(_06803_ ), .ZN(_00572_ ) );
NAND3_X1 _16336_ ( .A1(_00541_ ), .A2(_05298_ ), .A3(_00542_ ), .ZN(_00573_ ) );
NAND3_X1 _16337_ ( .A1(_00544_ ), .A2(_07246_ ), .A3(_00573_ ), .ZN(_00574_ ) );
AND2_X1 _16338_ ( .A1(_05297_ ), .A2(_07192_ ), .ZN(_00575_ ) );
NOR3_X1 _16339_ ( .A1(_07633_ ), .A2(_05296_ ), .A3(_07190_ ), .ZN(_00576_ ) );
AOI21_X1 _16340_ ( .A(_07130_ ), .B1(_07633_ ), .B2(_05296_ ), .ZN(_00577_ ) );
NOR3_X1 _16341_ ( .A1(_00575_ ), .A2(_00576_ ), .A3(_00577_ ), .ZN(_00578_ ) );
OR3_X1 _16342_ ( .A1(_07674_ ), .A2(_07675_ ), .A3(_06983_ ), .ZN(_00579_ ) );
OAI211_X1 _16343_ ( .A(_06995_ ), .B(_00579_ ), .C1(_07522_ ), .C2(_07315_ ), .ZN(_00580_ ) );
OR3_X1 _16344_ ( .A1(_07524_ ), .A2(_06986_ ), .A3(_06984_ ), .ZN(_00581_ ) );
AOI21_X1 _16345_ ( .A(_07045_ ), .B1(_00580_ ), .B2(_00581_ ), .ZN(_00582_ ) );
AND2_X1 _16346_ ( .A1(_07866_ ), .A2(_06986_ ), .ZN(_00583_ ) );
NOR3_X1 _16347_ ( .A1(_07863_ ), .A2(_06934_ ), .A3(_07097_ ), .ZN(_00584_ ) );
OR3_X1 _16348_ ( .A1(_07213_ ), .A2(_00584_ ), .A3(_00583_ ), .ZN(_00585_ ) );
AOI221_X4 _16349_ ( .A(_00582_ ), .B1(_06992_ ), .B2(_00583_ ), .C1(_00585_ ), .C2(_06882_ ), .ZN(_00586_ ) );
NAND3_X1 _16350_ ( .A1(_00574_ ), .A2(_00578_ ), .A3(_00586_ ), .ZN(_00587_ ) );
AOI21_X1 _16351_ ( .A(_00572_ ), .B1(_00587_ ), .B2(_07077_ ), .ZN(_00588_ ) );
OAI21_X1 _16352_ ( .A(_06502_ ), .B1(_06188_ ), .B2(_05601_ ), .ZN(_00589_ ) );
OAI21_X1 _16353_ ( .A(_00566_ ), .B1(_00588_ ), .B2(_00589_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NAND3_X1 _16354_ ( .A1(_05670_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_05671_ ), .ZN(_00590_ ) );
NAND4_X1 _16355_ ( .A1(_06060_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_06061_ ), .A4(_06063_ ), .ZN(_00591_ ) );
NAND4_X1 _16356_ ( .A1(_06060_ ), .A2(_05679_ ), .A3(\mtvec [31] ), .A4(_06061_ ), .ZN(_00592_ ) );
AND4_X1 _16357_ ( .A1(_06230_ ), .A2(_06231_ ), .A3(_00591_ ), .A4(_00592_ ), .ZN(_00593_ ) );
OAI21_X1 _16358_ ( .A(_00590_ ), .B1(_00593_ ), .B2(_05682_ ), .ZN(_00594_ ) );
NAND2_X1 _16359_ ( .A1(_00594_ ), .A2(_08008_ ), .ZN(_00595_ ) );
OR2_X1 _16360_ ( .A1(_06223_ ), .A2(_06788_ ), .ZN(_00596_ ) );
AOI21_X1 _16361_ ( .A(_05450_ ), .B1(_07618_ ), .B2(_04607_ ), .ZN(_00597_ ) );
XNOR2_X1 _16362_ ( .A(_00597_ ), .B(_04630_ ), .ZN(_00598_ ) );
AOI22_X1 _16363_ ( .A1(_00598_ ), .A2(_07445_ ), .B1(\ID_EX_imm [31] ), .B2(_07087_ ), .ZN(_00599_ ) );
AOI21_X1 _16364_ ( .A(_06803_ ), .B1(_00596_ ), .B2(_00599_ ), .ZN(_00600_ ) );
AOI21_X1 _16365_ ( .A(_07682_ ), .B1(_02399_ ), .B2(_02400_ ), .ZN(_00601_ ) );
OR3_X1 _16366_ ( .A1(_07651_ ), .A2(_05140_ ), .A3(_00601_ ), .ZN(_00602_ ) );
OAI21_X1 _16367_ ( .A(_05140_ ), .B1(_07651_ ), .B2(_00601_ ), .ZN(_00603_ ) );
NAND3_X1 _16368_ ( .A1(_00602_ ), .A2(_06878_ ), .A3(_00603_ ), .ZN(_00604_ ) );
NOR3_X1 _16369_ ( .A1(_07472_ ), .A2(_07060_ ), .A3(_07557_ ), .ZN(_00605_ ) );
AOI221_X4 _16370_ ( .A(_00605_ ), .B1(_05137_ ), .B2(_05129_ ), .C1(_05140_ ), .C2(_05467_ ), .ZN(_00606_ ) );
NAND3_X1 _16371_ ( .A1(_07475_ ), .A2(_07478_ ), .A3(_00426_ ), .ZN(_00607_ ) );
OR2_X1 _16372_ ( .A1(_05138_ ), .A2(_07065_ ), .ZN(_00608_ ) );
NAND3_X1 _16373_ ( .A1(_00606_ ), .A2(_00607_ ), .A3(_00608_ ), .ZN(_00609_ ) );
OAI211_X1 _16374_ ( .A(_06976_ ), .B(_06939_ ), .C1(_03243_ ), .C2(_06975_ ), .ZN(_00610_ ) );
OAI21_X1 _16375_ ( .A(_00610_ ), .B1(_08020_ ), .B2(_07141_ ), .ZN(_00611_ ) );
MUX2_X1 _16376_ ( .A(_00611_ ), .B(_00410_ ), .S(_06965_ ), .Z(_00612_ ) );
MUX2_X1 _16377_ ( .A(_00558_ ), .B(_00612_ ), .S(_07054_ ), .Z(_00613_ ) );
OAI22_X1 _16378_ ( .A1(_07398_ ), .A2(_07397_ ), .B1(_07146_ ), .B2(_07472_ ), .ZN(_00614_ ) );
AOI221_X4 _16379_ ( .A(_00609_ ), .B1(_07480_ ), .B2(_00613_ ), .C1(_00614_ ), .C2(_06882_ ), .ZN(_00615_ ) );
AOI21_X1 _16380_ ( .A(_07076_ ), .B1(_00604_ ), .B2(_00615_ ), .ZN(_00616_ ) );
NOR3_X1 _16381_ ( .A1(_00600_ ), .A2(_05553_ ), .A3(_00616_ ), .ZN(_00617_ ) );
NAND2_X1 _16382_ ( .A1(_06237_ ), .A2(_05838_ ), .ZN(_00618_ ) );
NAND2_X1 _16383_ ( .A1(_00618_ ), .A2(_06563_ ), .ZN(_00619_ ) );
OAI21_X1 _16384_ ( .A(_00595_ ), .B1(_00617_ ), .B2(_00619_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
NOR4_X1 _16385_ ( .A1(_03592_ ), .A2(reset ), .A3(excp_written ), .A4(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ) );
NAND2_X1 _16386_ ( .A1(_03617_ ), .A2(IDU_valid_EXU ), .ZN(_00620_ ) );
OAI21_X1 _16387_ ( .A(_00620_ ), .B1(_03493_ ), .B2(_03547_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16388_ ( .A1(_03545_ ), .A2(_03547_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16389_ ( .A1(_03545_ ), .A2(_03547_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16390_ ( .A(_03542_ ), .ZN(_00621_ ) );
NOR4_X1 _16391_ ( .A1(_03545_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03322_ ), .A4(_00621_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16392_ ( .A1(_03959_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03322_ ), .A4(_03541_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16393_ ( .A(_04098_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16394_ ( .A(_00620_ ), .B1(_00621_ ), .B2(_03617_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16395_ ( .A1(_03542_ ), .A2(_03617_ ), .B1(_02187_ ), .B2(_03592_ ), .ZN(_00622_ ) );
INV_X1 _16396_ ( .A(loaduse_clear ), .ZN(_00623_ ) );
AOI221_X4 _16397_ ( .A(_00622_ ), .B1(\myidu.state [2] ), .B2(_00623_ ), .C1(_03492_ ), .C2(_04098_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
NAND3_X1 _16398_ ( .A1(_03361_ ), .A2(IDU_valid_EXU ), .A3(_06276_ ), .ZN(_00624_ ) );
NAND3_X1 _16399_ ( .A1(_03361_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_00625_ ) );
INV_X1 _16400_ ( .A(_03607_ ), .ZN(_00626_ ) );
OR3_X1 _16401_ ( .A1(_03611_ ), .A2(_03612_ ), .A3(_03613_ ), .ZN(_00627_ ) );
AOI22_X1 _16402_ ( .A1(_03455_ ), .A2(_03489_ ), .B1(_00626_ ), .B2(_00627_ ), .ZN(_00628_ ) );
AOI21_X1 _16403_ ( .A(_00626_ ), .B1(_03475_ ), .B2(_03317_ ), .ZN(_00629_ ) );
OR2_X1 _16404_ ( .A1(_00628_ ), .A2(_00629_ ), .ZN(_00630_ ) );
NAND3_X1 _16405_ ( .A1(_03542_ ), .A2(IDU_ready_IFU ), .A3(_03321_ ), .ZN(_00631_ ) );
OAI211_X1 _16406_ ( .A(_00624_ ), .B(_00625_ ), .C1(_00630_ ), .C2(_00631_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16407_ ( .A(_03361_ ), .B(_04143_ ), .C1(_03542_ ), .C2(_03617_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
OAI221_X1 _16408_ ( .A(_03540_ ), .B1(_03607_ ), .B2(_03614_ ), .C1(_03536_ ), .C2(_03537_ ), .ZN(_00632_ ) );
AOI21_X1 _16409_ ( .A(_00632_ ), .B1(_03455_ ), .B2(_03489_ ), .ZN(_00633_ ) );
NAND3_X1 _16410_ ( .A1(_00633_ ), .A2(IDU_ready_IFU ), .A3(_03361_ ), .ZN(_00634_ ) );
NAND3_X1 _16411_ ( .A1(_03361_ ), .A2(\myidu.state [2] ), .A3(_00623_ ), .ZN(_00635_ ) );
NAND4_X1 _16412_ ( .A1(_03542_ ), .A2(_00629_ ), .A3(IDU_ready_IFU ), .A4(_03321_ ), .ZN(_00636_ ) );
NAND3_X1 _16413_ ( .A1(_00634_ ), .A2(_00635_ ), .A3(_00636_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16414_ ( .A1(_03539_ ), .A2(IDU_ready_IFU ), .ZN(_00637_ ) );
NOR2_X1 _16415_ ( .A1(_03539_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00638_ ) );
NOR2_X1 _16416_ ( .A1(\myifu.state [0] ), .A2(\myifu.state [1] ), .ZN(_00639_ ) );
NOR4_X1 _16417_ ( .A1(_00637_ ), .A2(_00638_ ), .A3(reset ), .A4(_00639_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
CLKBUF_X2 _16418_ ( .A(_06342_ ), .Z(_00640_ ) );
OR3_X1 _16419_ ( .A1(_02205_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00641_ ) );
OAI21_X1 _16420_ ( .A(_00641_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06343_ ), .ZN(_00642_ ) );
MUX2_X1 _16421_ ( .A(\io_master_rdata [31] ), .B(_00642_ ), .S(_04080_ ), .Z(_00643_ ) );
AND2_X1 _16422_ ( .A1(_00643_ ), .A2(_06297_ ), .ZN(\myifu.data_in [31] ) );
OR3_X1 _16423_ ( .A1(_02205_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00644_ ) );
OAI211_X1 _16424_ ( .A(_02226_ ), .B(_00644_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06344_ ), .ZN(_00645_ ) );
OAI21_X1 _16425_ ( .A(_00645_ ), .B1(_02227_ ), .B2(\io_master_rdata [30] ), .ZN(_00646_ ) );
NOR2_X1 _16426_ ( .A1(_00646_ ), .A2(_06311_ ), .ZN(\myifu.data_in [30] ) );
CLKBUF_X2 _16427_ ( .A(_02227_ ), .Z(_00647_ ) );
OR2_X1 _16428_ ( .A1(_00647_ ), .A2(\io_master_rdata [21] ), .ZN(_00648_ ) );
CLKBUF_X2 _16429_ ( .A(_02231_ ), .Z(_00649_ ) );
CLKBUF_X2 _16430_ ( .A(_00640_ ), .Z(_00650_ ) );
OR3_X1 _16431_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00651_ ) );
BUF_X4 _16432_ ( .A(_06344_ ), .Z(_00652_ ) );
OAI211_X1 _16433_ ( .A(_02228_ ), .B(_00651_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00653_ ) );
AND3_X1 _16434_ ( .A1(_00648_ ), .A2(_00653_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [21] ) );
OR2_X1 _16435_ ( .A1(_02227_ ), .A2(\io_master_rdata [20] ), .ZN(_00654_ ) );
OR3_X1 _16436_ ( .A1(_02231_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00655_ ) );
OAI211_X1 _16437_ ( .A(_00647_ ), .B(_00655_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06344_ ), .ZN(_00656_ ) );
AND3_X1 _16438_ ( .A1(_00654_ ), .A2(_00656_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [20] ) );
OR2_X1 _16439_ ( .A1(_00647_ ), .A2(\io_master_rdata [19] ), .ZN(_00657_ ) );
OR3_X1 _16440_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00658_ ) );
OAI211_X1 _16441_ ( .A(_02228_ ), .B(_00658_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00659_ ) );
AND3_X1 _16442_ ( .A1(_00657_ ), .A2(_00659_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [19] ) );
OR2_X1 _16443_ ( .A1(_00647_ ), .A2(\io_master_rdata [18] ), .ZN(_00660_ ) );
OR3_X1 _16444_ ( .A1(_02231_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00661_ ) );
OAI211_X1 _16445_ ( .A(_02228_ ), .B(_00661_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00662_ ) );
AND3_X1 _16446_ ( .A1(_00660_ ), .A2(_00662_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [18] ) );
OR2_X1 _16447_ ( .A1(_00647_ ), .A2(\io_master_rdata [17] ), .ZN(_00663_ ) );
OR3_X1 _16448_ ( .A1(_02231_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00664_ ) );
OAI211_X1 _16449_ ( .A(_02228_ ), .B(_00664_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00665_ ) );
AND3_X1 _16450_ ( .A1(_00663_ ), .A2(_00665_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [17] ) );
OR2_X1 _16451_ ( .A1(_00647_ ), .A2(\io_master_rdata [16] ), .ZN(_00666_ ) );
OR3_X1 _16452_ ( .A1(_02231_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00667_ ) );
OAI211_X1 _16453_ ( .A(_02228_ ), .B(_00667_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00668_ ) );
AND3_X1 _16454_ ( .A1(_00666_ ), .A2(_00668_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16455_ ( .A1(_02205_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00669_ ) );
OAI211_X1 _16456_ ( .A(_02226_ ), .B(_00669_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06343_ ), .ZN(_00670_ ) );
OAI21_X1 _16457_ ( .A(_00670_ ), .B1(_02226_ ), .B2(\io_master_rdata [15] ), .ZN(_00671_ ) );
BUF_X4 _16458_ ( .A(_06311_ ), .Z(_00672_ ) );
NOR2_X1 _16459_ ( .A1(_00671_ ), .A2(_00672_ ), .ZN(\myifu.data_in [15] ) );
OR2_X1 _16460_ ( .A1(_02227_ ), .A2(\io_master_rdata [14] ), .ZN(_00673_ ) );
OR3_X1 _16461_ ( .A1(_02231_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00674_ ) );
OAI211_X1 _16462_ ( .A(_02227_ ), .B(_00674_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06344_ ), .ZN(_00675_ ) );
AND3_X1 _16463_ ( .A1(_00673_ ), .A2(_00675_ ), .A3(_02232_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16464_ ( .A1(_00647_ ), .A2(\io_master_rdata [13] ), .ZN(_00676_ ) );
OR3_X1 _16465_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00677_ ) );
OAI211_X1 _16466_ ( .A(_02228_ ), .B(_00677_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00678_ ) );
AND3_X1 _16467_ ( .A1(_00676_ ), .A2(_00678_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [13] ) );
BUF_X2 _16468_ ( .A(_02227_ ), .Z(_00679_ ) );
OR2_X1 _16469_ ( .A1(_00679_ ), .A2(\io_master_rdata [12] ), .ZN(_00680_ ) );
CLKBUF_X2 _16470_ ( .A(_00640_ ), .Z(_00681_ ) );
OR3_X1 _16471_ ( .A1(_02232_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00682_ ) );
OAI211_X1 _16472_ ( .A(_02229_ ), .B(_00682_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00683_ ) );
AND3_X1 _16473_ ( .A1(_00680_ ), .A2(_00683_ ), .A3(_06297_ ), .ZN(\myifu.data_in [12] ) );
MUX2_X1 _16474_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06344_ ), .Z(_00684_ ) );
OR3_X1 _16475_ ( .A1(_06253_ ), .A2(_06256_ ), .A3(_00684_ ), .ZN(_00685_ ) );
OAI21_X1 _16476_ ( .A(\io_master_rdata [29] ), .B1(_04076_ ), .B2(_04079_ ), .ZN(_00686_ ) );
AOI21_X1 _16477_ ( .A(_00672_ ), .B1(_00685_ ), .B2(_00686_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16478_ ( .A1(_00679_ ), .A2(\io_master_rdata [11] ), .ZN(_00687_ ) );
OR3_X1 _16479_ ( .A1(_02232_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00688_ ) );
OAI211_X1 _16480_ ( .A(_02229_ ), .B(_00688_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00689_ ) );
AND3_X1 _16481_ ( .A1(_00687_ ), .A2(_00689_ ), .A3(_06297_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16482_ ( .A1(_00647_ ), .A2(\io_master_rdata [10] ), .ZN(_00690_ ) );
OR3_X1 _16483_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00691_ ) );
OAI211_X1 _16484_ ( .A(_02228_ ), .B(_00691_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00692_ ) );
AND3_X1 _16485_ ( .A1(_00690_ ), .A2(_00692_ ), .A3(_06297_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16486_ ( .A1(_02228_ ), .A2(\io_master_rdata [9] ), .ZN(_00693_ ) );
OR3_X1 _16487_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00694_ ) );
OAI211_X1 _16488_ ( .A(_00679_ ), .B(_00694_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00695_ ) );
AND3_X1 _16489_ ( .A1(_00693_ ), .A2(_00695_ ), .A3(_06297_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16490_ ( .A1(_00679_ ), .A2(\io_master_rdata [8] ), .ZN(_00696_ ) );
OR3_X1 _16491_ ( .A1(_02232_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00697_ ) );
OAI211_X1 _16492_ ( .A(_02229_ ), .B(_00697_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00698_ ) );
AND3_X1 _16493_ ( .A1(_00696_ ), .A2(_00698_ ), .A3(_06297_ ), .ZN(\myifu.data_in [8] ) );
OR2_X2 _16494_ ( .A1(_02226_ ), .A2(\io_master_rdata [7] ), .ZN(_00699_ ) );
OR3_X1 _16495_ ( .A1(_02205_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00700_ ) );
OAI211_X2 _16496_ ( .A(_02226_ ), .B(_00700_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06343_ ), .ZN(_00701_ ) );
AND3_X1 _16497_ ( .A1(_00699_ ), .A2(_00701_ ), .A3(_06297_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16498_ ( .A1(_02205_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00702_ ) );
OAI211_X1 _16499_ ( .A(_02226_ ), .B(_00702_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06343_ ), .ZN(_00703_ ) );
OAI21_X1 _16500_ ( .A(_00703_ ), .B1(_02227_ ), .B2(\io_master_rdata [6] ), .ZN(_00704_ ) );
NOR2_X1 _16501_ ( .A1(_00704_ ), .A2(_06311_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16502_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00705_ ) );
OAI211_X1 _16503_ ( .A(_00679_ ), .B(_00705_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00706_ ) );
OAI21_X1 _16504_ ( .A(_00706_ ), .B1(_02229_ ), .B2(\io_master_rdata [5] ), .ZN(_00707_ ) );
NOR2_X1 _16505_ ( .A1(_00707_ ), .A2(_00672_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16506_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00708_ ) );
OAI211_X1 _16507_ ( .A(_02228_ ), .B(_00708_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00709_ ) );
OAI21_X1 _16508_ ( .A(_00709_ ), .B1(_00679_ ), .B2(\io_master_rdata [4] ), .ZN(_00710_ ) );
NOR2_X1 _16509_ ( .A1(_00710_ ), .A2(_00672_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16510_ ( .A1(_02232_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00711_ ) );
OAI211_X1 _16511_ ( .A(_02229_ ), .B(_00711_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00712_ ) );
OAI21_X1 _16512_ ( .A(_00712_ ), .B1(_02229_ ), .B2(\io_master_rdata [3] ), .ZN(_00713_ ) );
NOR2_X1 _16513_ ( .A1(_00713_ ), .A2(_00672_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16514_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00714_ ) );
OAI211_X1 _16515_ ( .A(_00679_ ), .B(_00714_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00715_ ) );
OAI21_X1 _16516_ ( .A(_00715_ ), .B1(_02229_ ), .B2(\io_master_rdata [2] ), .ZN(_00716_ ) );
NOR2_X1 _16517_ ( .A1(_00716_ ), .A2(_00672_ ), .ZN(\myifu.data_in [2] ) );
OR2_X1 _16518_ ( .A1(_02227_ ), .A2(\io_master_rdata [28] ), .ZN(_00717_ ) );
OR3_X1 _16519_ ( .A1(_02231_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00718_ ) );
OAI211_X1 _16520_ ( .A(_00647_ ), .B(_00718_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00652_ ), .ZN(_00719_ ) );
AND3_X1 _16521_ ( .A1(_00717_ ), .A2(_00719_ ), .A3(_02232_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16522_ ( .A1(_00649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00681_ ), .ZN(_00720_ ) );
OAI211_X1 _16523_ ( .A(_00679_ ), .B(_00720_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00721_ ) );
OAI21_X1 _16524_ ( .A(_00721_ ), .B1(_02229_ ), .B2(\io_master_rdata [1] ), .ZN(_00722_ ) );
NOR2_X1 _16525_ ( .A1(_00722_ ), .A2(_00672_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16526_ ( .A1(_00649_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00681_ ), .ZN(_00723_ ) );
OAI211_X1 _16527_ ( .A(_00679_ ), .B(_00723_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00724_ ) );
OAI21_X1 _16528_ ( .A(_00724_ ), .B1(\io_master_rdata [0] ), .B2(_00679_ ), .ZN(_00725_ ) );
NOR2_X1 _16529_ ( .A1(_00725_ ), .A2(_00672_ ), .ZN(\myifu.data_in [0] ) );
MUX2_X1 _16530_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06344_ ), .Z(_00726_ ) );
OR3_X1 _16531_ ( .A1(_06253_ ), .A2(_06256_ ), .A3(_00726_ ), .ZN(_00727_ ) );
OAI21_X1 _16532_ ( .A(\io_master_rdata [27] ), .B1(_04076_ ), .B2(_04079_ ), .ZN(_00728_ ) );
AOI21_X1 _16533_ ( .A(_06312_ ), .B1(_00727_ ), .B2(_00728_ ), .ZN(\myifu.data_in [27] ) );
OR3_X1 _16534_ ( .A1(_02231_ ), .A2(_01866_ ), .A3(_00650_ ), .ZN(_00729_ ) );
OAI211_X1 _16535_ ( .A(_06257_ ), .B(_00729_ ), .C1(_01853_ ), .C2(_00652_ ), .ZN(_00730_ ) );
OAI21_X1 _16536_ ( .A(\io_master_rdata [26] ), .B1(_04076_ ), .B2(_04079_ ), .ZN(_00731_ ) );
AOI21_X1 _16537_ ( .A(_06310_ ), .B1(_00730_ ), .B2(_00731_ ), .ZN(\myifu.data_in [26] ) );
MUX2_X1 _16538_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06344_ ), .Z(_00732_ ) );
OR3_X1 _16539_ ( .A1(_06253_ ), .A2(_06256_ ), .A3(_00732_ ), .ZN(_00733_ ) );
OAI21_X1 _16540_ ( .A(\io_master_rdata [25] ), .B1(_04076_ ), .B2(_04079_ ), .ZN(_00734_ ) );
AOI21_X1 _16541_ ( .A(_06310_ ), .B1(_00733_ ), .B2(_00734_ ), .ZN(\myifu.data_in [25] ) );
OR2_X1 _16542_ ( .A1(_02227_ ), .A2(\io_master_rdata [24] ), .ZN(_00735_ ) );
OR3_X1 _16543_ ( .A1(_02231_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00650_ ), .ZN(_00736_ ) );
OAI211_X1 _16544_ ( .A(_00647_ ), .B(_00736_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06344_ ), .ZN(_00737_ ) );
AND3_X1 _16545_ ( .A1(_00735_ ), .A2(_00737_ ), .A3(_02232_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16546_ ( .A1(_02205_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06342_ ), .ZN(_00738_ ) );
OAI211_X1 _16547_ ( .A(_02225_ ), .B(_00738_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06343_ ), .ZN(_00739_ ) );
OAI21_X1 _16548_ ( .A(_00739_ ), .B1(_02226_ ), .B2(\io_master_rdata [23] ), .ZN(_00740_ ) );
NOR2_X1 _16549_ ( .A1(_00740_ ), .A2(_00672_ ), .ZN(\myifu.data_in [23] ) );
OR3_X1 _16550_ ( .A1(_02205_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00640_ ), .ZN(_00741_ ) );
OAI211_X1 _16551_ ( .A(_02226_ ), .B(_00741_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06344_ ), .ZN(_00742_ ) );
OAI21_X1 _16552_ ( .A(_00742_ ), .B1(\io_master_rdata [22] ), .B2(_02226_ ), .ZN(_00743_ ) );
NOR2_X1 _16553_ ( .A1(_00743_ ), .A2(_00672_ ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16554_ ( .A(_00278_ ), .ZN(_00744_ ) );
NAND2_X1 _16555_ ( .A1(_00744_ ), .A2(_02268_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16556_ ( .A1(_04014_ ), .A2(fanout_net_9 ), .ZN(_00745_ ) );
INV_X1 _16557_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00746_ ) );
OAI21_X1 _16558_ ( .A(_02268_ ), .B1(_00745_ ), .B2(_00746_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16559_ ( .A1(_04021_ ), .A2(fanout_net_13 ), .ZN(_00747_ ) );
OAI21_X1 _16560_ ( .A(_02268_ ), .B1(_00747_ ), .B2(_00746_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16561_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .ZN(_00748_ ) );
OAI21_X1 _16562_ ( .A(_02268_ ), .B1(_00748_ ), .B2(_00746_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
OAI21_X1 _16563_ ( .A(\IF_ID_inst [8] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00749_ ) );
NOR2_X1 _16564_ ( .A1(_03481_ ), .A2(_03619_ ), .ZN(_00750_ ) );
AND2_X1 _16565_ ( .A1(_00750_ ), .A2(_03667_ ), .ZN(_00751_ ) );
INV_X1 _16566_ ( .A(_03654_ ), .ZN(_00752_ ) );
NAND3_X1 _16567_ ( .A1(_03627_ ), .A2(_03690_ ), .A3(_03381_ ), .ZN(_00753_ ) );
NAND4_X1 _16568_ ( .A1(_00752_ ), .A2(_03317_ ), .A3(_00753_ ), .A4(_03628_ ), .ZN(_00754_ ) );
NAND3_X1 _16569_ ( .A1(_03638_ ), .A2(_03650_ ), .A3(_03641_ ), .ZN(_00755_ ) );
NOR2_X1 _16570_ ( .A1(_00754_ ), .A2(_00755_ ), .ZN(_00756_ ) );
NAND3_X1 _16571_ ( .A1(_00751_ ), .A2(_00756_ ), .A3(_03806_ ), .ZN(_00757_ ) );
AND2_X1 _16572_ ( .A1(_00757_ ), .A2(_03806_ ), .ZN(_00758_ ) );
OAI221_X1 _16573_ ( .A(_00749_ ), .B1(_03549_ ), .B2(_03318_ ), .C1(_00758_ ), .C2(_03325_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
AND2_X1 _16574_ ( .A1(_03405_ ), .A2(\IF_ID_inst [31] ), .ZN(_00759_ ) );
INV_X1 _16575_ ( .A(_00759_ ), .ZN(_00760_ ) );
BUF_X4 _16576_ ( .A(_00760_ ), .Z(_00761_ ) );
NOR2_X1 _16577_ ( .A1(_03475_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_00762_ ) );
INV_X1 _16578_ ( .A(_00762_ ), .ZN(_00763_ ) );
OAI211_X1 _16579_ ( .A(_00761_ ), .B(_00763_ ), .C1(_00751_ ), .C2(_03319_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
OAI21_X1 _16580_ ( .A(\IF_ID_inst [31] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00764_ ) );
AND2_X1 _16581_ ( .A1(_00763_ ), .A2(_00764_ ), .ZN(_00765_ ) );
BUF_X4 _16582_ ( .A(_00765_ ), .Z(_00766_ ) );
BUF_X4 _16583_ ( .A(_03667_ ), .Z(_00767_ ) );
OAI211_X1 _16584_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03324_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16585_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03325_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16586_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03328_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
BUF_X4 _16587_ ( .A(_03475_ ), .Z(_00768_ ) );
OAI221_X1 _16588_ ( .A(_00764_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00768_ ), .C1(_03395_ ), .C2(_03406_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI221_X1 _16589_ ( .A(_00764_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00768_ ), .C1(_03416_ ), .C2(_03406_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI221_X1 _16590_ ( .A(_00764_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00768_ ), .C1(_03417_ ), .C2(_03406_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16591_ ( .A(_00764_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00768_ ), .C1(_03549_ ), .C2(_03406_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _16592_ ( .A(_00764_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00768_ ), .C1(_03410_ ), .C2(_03406_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16593_ ( .A(_00764_ ), .B1(_03431_ ), .B2(_03406_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .C2(_00768_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16594_ ( .A(_00764_ ), .B1(_03353_ ), .B2(_03406_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .C2(_00768_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16595_ ( .A(_00764_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_03475_ ), .C1(_03346_ ), .C2(_03406_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16596_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03329_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
AND3_X1 _16597_ ( .A1(_03482_ ), .A2(\IF_ID_inst [7] ), .A3(_03458_ ), .ZN(_00769_ ) );
AOI21_X1 _16598_ ( .A(_03319_ ), .B1(_03478_ ), .B2(_03479_ ), .ZN(_00770_ ) );
OR4_X1 _16599_ ( .A1(_03758_ ), .A2(_00762_ ), .A3(_00769_ ), .A4(_00770_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16600_ ( .A(_03773_ ), .ZN(_00771_ ) );
OAI221_X1 _16601_ ( .A(_00771_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_03475_ ), .C1(_00750_ ), .C2(_03324_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
OAI221_X1 _16602_ ( .A(_03767_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03475_ ), .C1(_00750_ ), .C2(_03329_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
OAI21_X1 _16603_ ( .A(\IF_ID_inst [28] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00772_ ) );
OAI221_X1 _16604_ ( .A(_00772_ ), .B1(_03330_ ), .B2(_03806_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .C2(_00768_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
OAI21_X1 _16605_ ( .A(\IF_ID_inst [27] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00773_ ) );
OAI221_X1 _16606_ ( .A(_00773_ ), .B1(_03331_ ), .B2(_03806_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00768_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
OAI21_X1 _16607_ ( .A(\IF_ID_inst [26] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00774_ ) );
OAI221_X1 _16608_ ( .A(_00774_ ), .B1(_03332_ ), .B2(_03806_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .C2(_00768_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16609_ ( .A(_03778_ ), .ZN(_00775_ ) );
OAI221_X1 _16610_ ( .A(_00775_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .B2(_03475_ ), .C1(_00750_ ), .C2(_03333_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16611_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03330_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16612_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03331_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16613_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03332_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16614_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03333_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16615_ ( .A(_00766_ ), .B(_00761_ ), .C1(_03335_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16616_ ( .A(_00766_ ), .B(_00760_ ), .C1(_03336_ ), .C2(_00767_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16617_ ( .A(_00765_ ), .B(_00760_ ), .C1(_03337_ ), .C2(_03667_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16618_ ( .A(\IF_ID_inst [11] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00776_ ) );
OAI221_X1 _16619_ ( .A(_00776_ ), .B1(_03395_ ), .B2(_03317_ ), .C1(_00758_ ), .C2(_03335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16620_ ( .A(\IF_ID_inst [10] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00777_ ) );
OAI221_X1 _16621_ ( .A(_00777_ ), .B1(_03416_ ), .B2(_03317_ ), .C1(_00758_ ), .C2(_03336_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16622_ ( .A(\IF_ID_inst [9] ), .B1(_03481_ ), .B2(_03619_ ), .ZN(_00778_ ) );
OAI221_X1 _16623_ ( .A(_00778_ ), .B1(_03417_ ), .B2(_03317_ ), .C1(_00758_ ), .C2(_03337_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16624_ ( .A1(_03480_ ), .A2(_03362_ ), .ZN(_00779_ ) );
OAI221_X1 _16625_ ( .A(_00779_ ), .B1(_03410_ ), .B2(_03317_ ), .C1(_00757_ ), .C2(_03328_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AND3_X1 _16626_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00780_ ) );
CLKBUF_X2 _16627_ ( .A(_04011_ ), .Z(_00781_ ) );
AND3_X1 _16628_ ( .A1(_00781_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00782_ ) );
BUF_X4 _16629_ ( .A(_06268_ ), .Z(_00783_ ) );
BUF_X4 _16630_ ( .A(_00783_ ), .Z(_00784_ ) );
AOI211_X1 _16631_ ( .A(_00780_ ), .B(_00782_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_00784_ ), .ZN(_00785_ ) );
NAND2_X1 _16632_ ( .A1(_00746_ ), .A2(\IF_ID_pc [2] ), .ZN(_00786_ ) );
BUF_X4 _16633_ ( .A(_00786_ ), .Z(_00787_ ) );
BUF_X4 _16634_ ( .A(_00787_ ), .Z(_00788_ ) );
NAND2_X1 _16635_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00789_ ) );
BUF_X4 _16636_ ( .A(_00789_ ), .Z(_00790_ ) );
BUF_X4 _16637_ ( .A(_00790_ ), .Z(_00791_ ) );
BUF_X4 _16638_ ( .A(_03799_ ), .Z(_00792_ ) );
BUF_X4 _16639_ ( .A(_00792_ ), .Z(_00793_ ) );
BUF_X4 _16640_ ( .A(_00793_ ), .Z(_00794_ ) );
NAND3_X1 _16641_ ( .A1(_00794_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00795_ ) );
NAND4_X1 _16642_ ( .A1(_00785_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_00795_ ), .ZN(_00796_ ) );
NOR2_X1 _16643_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00797_ ) );
BUF_X4 _16644_ ( .A(_00797_ ), .Z(_00798_ ) );
BUF_X4 _16645_ ( .A(_00798_ ), .Z(_00799_ ) );
BUF_X4 _16646_ ( .A(_04011_ ), .Z(_00800_ ) );
BUF_X4 _16647_ ( .A(_00800_ ), .Z(_00801_ ) );
NAND3_X1 _16648_ ( .A1(_00801_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00802_ ) );
NAND3_X1 _16649_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00803_ ) );
AND2_X1 _16650_ ( .A1(_00802_ ), .A2(_00803_ ), .ZN(_00804_ ) );
NAND2_X1 _16651_ ( .A1(_00786_ ), .A2(_00789_ ), .ZN(_00805_ ) );
BUF_X4 _16652_ ( .A(_00805_ ), .Z(_00806_ ) );
BUF_X4 _16653_ ( .A(_00806_ ), .Z(_00807_ ) );
BUF_X4 _16654_ ( .A(_04020_ ), .Z(_00808_ ) );
NAND3_X1 _16655_ ( .A1(_00808_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00809_ ) );
BUF_X4 _16656_ ( .A(_04012_ ), .Z(_00810_ ) );
BUF_X4 _16657_ ( .A(_00810_ ), .Z(_00811_ ) );
BUF_X4 _16658_ ( .A(_00792_ ), .Z(_00812_ ) );
NAND3_X1 _16659_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00813_ ) );
NAND4_X1 _16660_ ( .A1(_00804_ ), .A2(_00807_ ), .A3(_00809_ ), .A4(_00813_ ), .ZN(_00814_ ) );
NAND3_X1 _16661_ ( .A1(_00796_ ), .A2(_00799_ ), .A3(_00814_ ), .ZN(_00815_ ) );
XOR2_X1 _16662_ ( .A(\IF_ID_pc [2] ), .B(\myifu.tmp_offset [2] ), .Z(_00816_ ) );
NAND2_X1 _16663_ ( .A1(_03791_ ), .A2(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .ZN(_00817_ ) );
NOR2_X2 _16664_ ( .A1(_00816_ ), .A2(_00817_ ), .ZN(_00818_ ) );
AND2_X2 _16665_ ( .A1(_04090_ ), .A2(_00818_ ), .ZN(_00819_ ) );
INV_X1 _16666_ ( .A(_00819_ ), .ZN(_00820_ ) );
BUF_X4 _16667_ ( .A(_00820_ ), .Z(_00821_ ) );
NOR2_X1 _16668_ ( .A1(_00821_ ), .A2(\myifu.data_in [8] ), .ZN(_00822_ ) );
BUF_X4 _16669_ ( .A(_00819_ ), .Z(_00823_ ) );
OAI21_X1 _16670_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03788_ ), .ZN(_00824_ ) );
OAI21_X1 _16671_ ( .A(_00815_ ), .B1(_00822_ ), .B2(_00824_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16672_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00825_ ) );
AND3_X1 _16673_ ( .A1(_00781_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00826_ ) );
AOI211_X1 _16674_ ( .A(_00825_ ), .B(_00826_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00783_ ), .ZN(_00827_ ) );
NAND3_X1 _16675_ ( .A1(_00794_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00828_ ) );
NAND4_X1 _16676_ ( .A1(_00827_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_00828_ ), .ZN(_00829_ ) );
NAND3_X1 _16677_ ( .A1(_00801_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00830_ ) );
NAND3_X1 _16678_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00831_ ) );
AND2_X1 _16679_ ( .A1(_00830_ ), .A2(_00831_ ), .ZN(_00832_ ) );
NAND3_X1 _16680_ ( .A1(_00808_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00833_ ) );
NAND3_X1 _16681_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00834_ ) );
NAND4_X1 _16682_ ( .A1(_00832_ ), .A2(_00807_ ), .A3(_00833_ ), .A4(_00834_ ), .ZN(_00835_ ) );
NAND3_X1 _16683_ ( .A1(_00829_ ), .A2(_00799_ ), .A3(_00835_ ), .ZN(_00836_ ) );
NOR2_X1 _16684_ ( .A1(_00821_ ), .A2(\myifu.data_in [31] ), .ZN(_00837_ ) );
OAI21_X1 _16685_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03658_ ), .ZN(_00838_ ) );
OAI21_X1 _16686_ ( .A(_00836_ ), .B1(_00837_ ), .B2(_00838_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
AND3_X1 _16687_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00839_ ) );
AND3_X1 _16688_ ( .A1(_00781_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00840_ ) );
AOI211_X1 _16689_ ( .A(_00839_ ), .B(_00840_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_00783_ ), .ZN(_00841_ ) );
NAND3_X1 _16690_ ( .A1(_00794_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00842_ ) );
NAND4_X1 _16691_ ( .A1(_00841_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_00842_ ), .ZN(_00843_ ) );
NAND3_X1 _16692_ ( .A1(_00801_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00844_ ) );
NAND3_X1 _16693_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00845_ ) );
AND2_X1 _16694_ ( .A1(_00844_ ), .A2(_00845_ ), .ZN(_00846_ ) );
NAND3_X1 _16695_ ( .A1(_00808_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00847_ ) );
NAND3_X1 _16696_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00848_ ) );
NAND4_X1 _16697_ ( .A1(_00846_ ), .A2(_00807_ ), .A3(_00847_ ), .A4(_00848_ ), .ZN(_00849_ ) );
NAND3_X1 _16698_ ( .A1(_00843_ ), .A2(_00799_ ), .A3(_00849_ ), .ZN(_00850_ ) );
NOR2_X1 _16699_ ( .A1(_00821_ ), .A2(\myifu.data_in [30] ), .ZN(_00851_ ) );
OAI21_X1 _16700_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03774_ ), .ZN(_00852_ ) );
OAI21_X1 _16701_ ( .A(_00850_ ), .B1(_00851_ ), .B2(_00852_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
INV_X1 _16702_ ( .A(\myifu.state [2] ), .ZN(_00853_ ) );
BUF_X4 _16703_ ( .A(_00853_ ), .Z(_00854_ ) );
BUF_X2 _16704_ ( .A(_00820_ ), .Z(_00855_ ) );
AOI21_X1 _16705_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00856_ ) );
BUF_X4 _16706_ ( .A(_00819_ ), .Z(_00857_ ) );
NAND2_X1 _16707_ ( .A1(_00648_ ), .A2(_00653_ ), .ZN(_00858_ ) );
OAI21_X1 _16708_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_00858_ ), .ZN(_00859_ ) );
NAND2_X1 _16709_ ( .A1(_00856_ ), .A2(_00859_ ), .ZN(_00860_ ) );
AND3_X1 _16710_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00861_ ) );
AND3_X1 _16711_ ( .A1(_04013_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00862_ ) );
AOI211_X1 _16712_ ( .A(_00861_ ), .B(_00862_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_06269_ ), .ZN(_00863_ ) );
BUF_X2 _16713_ ( .A(_00786_ ), .Z(_00864_ ) );
BUF_X4 _16714_ ( .A(_00790_ ), .Z(_00865_ ) );
NAND3_X1 _16715_ ( .A1(_04021_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00866_ ) );
NAND4_X1 _16716_ ( .A1(_00863_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_00866_ ), .ZN(_00867_ ) );
BUF_X4 _16717_ ( .A(_00798_ ), .Z(_00868_ ) );
BUF_X4 _16718_ ( .A(_00800_ ), .Z(_00869_ ) );
NAND3_X1 _16719_ ( .A1(_00869_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00870_ ) );
NAND3_X1 _16720_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00871_ ) );
AND2_X1 _16721_ ( .A1(_00870_ ), .A2(_00871_ ), .ZN(_00872_ ) );
BUF_X2 _16722_ ( .A(_00805_ ), .Z(_00873_ ) );
BUF_X4 _16723_ ( .A(_00793_ ), .Z(_00874_ ) );
NAND3_X1 _16724_ ( .A1(_00874_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00875_ ) );
BUF_X4 _16725_ ( .A(_04020_ ), .Z(_00876_ ) );
NAND3_X1 _16726_ ( .A1(_04014_ ), .A2(_00876_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00877_ ) );
NAND4_X1 _16727_ ( .A1(_00872_ ), .A2(_00873_ ), .A3(_00875_ ), .A4(_00877_ ), .ZN(_00878_ ) );
NAND3_X1 _16728_ ( .A1(_00867_ ), .A2(_00868_ ), .A3(_00878_ ), .ZN(_00879_ ) );
NAND2_X1 _16729_ ( .A1(_00860_ ), .A2(_00879_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
NAND2_X1 _16730_ ( .A1(_00654_ ), .A2(_00656_ ), .ZN(_00880_ ) );
OAI211_X1 _16731_ ( .A(_04091_ ), .B(_00818_ ), .C1(_00880_ ), .C2(_06310_ ), .ZN(_00881_ ) );
NAND2_X1 _16732_ ( .A1(_00881_ ), .A2(\myifu.state [2] ), .ZN(_00882_ ) );
BUF_X4 _16733_ ( .A(_00820_ ), .Z(_00883_ ) );
AOI21_X1 _16734_ ( .A(_00882_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00883_ ), .ZN(_00884_ ) );
AND3_X1 _16735_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00885_ ) );
AND3_X1 _16736_ ( .A1(_04012_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00886_ ) );
AOI211_X1 _16737_ ( .A(_00885_ ), .B(_00886_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_06268_ ), .ZN(_00887_ ) );
NAND3_X1 _16738_ ( .A1(_00793_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00888_ ) );
NAND4_X1 _16739_ ( .A1(_00887_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_00888_ ), .ZN(_00889_ ) );
NAND3_X1 _16740_ ( .A1(_00800_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00890_ ) );
NAND3_X1 _16741_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00891_ ) );
AND2_X1 _16742_ ( .A1(_00890_ ), .A2(_00891_ ), .ZN(_00892_ ) );
NAND3_X1 _16743_ ( .A1(_04020_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00893_ ) );
NAND3_X1 _16744_ ( .A1(_00810_ ), .A2(_00792_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00894_ ) );
NAND4_X1 _16745_ ( .A1(_00892_ ), .A2(_00806_ ), .A3(_00893_ ), .A4(_00894_ ), .ZN(_00895_ ) );
AND3_X1 _16746_ ( .A1(_00889_ ), .A2(_00798_ ), .A3(_00895_ ), .ZN(_00896_ ) );
OR2_X1 _16747_ ( .A1(_00884_ ), .A2(_00896_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
AOI21_X1 _16748_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00897_ ) );
NAND2_X1 _16749_ ( .A1(_00657_ ), .A2(_00659_ ), .ZN(_00898_ ) );
OAI21_X1 _16750_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_00898_ ), .ZN(_00899_ ) );
NAND2_X1 _16751_ ( .A1(_00897_ ), .A2(_00899_ ), .ZN(_00900_ ) );
AND3_X1 _16752_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00901_ ) );
AND3_X1 _16753_ ( .A1(_04013_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00902_ ) );
AOI211_X1 _16754_ ( .A(_00901_ ), .B(_00902_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_06269_ ), .ZN(_00903_ ) );
NAND3_X1 _16755_ ( .A1(_04021_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00904_ ) );
NAND4_X1 _16756_ ( .A1(_00903_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_00904_ ), .ZN(_00905_ ) );
NAND3_X1 _16757_ ( .A1(_00869_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00906_ ) );
NAND3_X1 _16758_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00907_ ) );
AND2_X1 _16759_ ( .A1(_00906_ ), .A2(_00907_ ), .ZN(_00908_ ) );
NAND3_X1 _16760_ ( .A1(_00874_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00909_ ) );
NAND3_X1 _16761_ ( .A1(_04014_ ), .A2(_00876_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00910_ ) );
NAND4_X1 _16762_ ( .A1(_00908_ ), .A2(_00873_ ), .A3(_00909_ ), .A4(_00910_ ), .ZN(_00911_ ) );
NAND3_X1 _16763_ ( .A1(_00905_ ), .A2(_00868_ ), .A3(_00911_ ), .ZN(_00912_ ) );
NAND2_X1 _16764_ ( .A1(_00900_ ), .A2(_00912_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
NAND2_X1 _16765_ ( .A1(_00660_ ), .A2(_00662_ ), .ZN(_00913_ ) );
OAI211_X1 _16766_ ( .A(_04091_ ), .B(_00818_ ), .C1(_00913_ ), .C2(_06310_ ), .ZN(_00914_ ) );
NAND2_X1 _16767_ ( .A1(_00914_ ), .A2(\myifu.state [2] ), .ZN(_00915_ ) );
AOI21_X1 _16768_ ( .A(_00915_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00883_ ), .ZN(_00916_ ) );
AND3_X1 _16769_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00917_ ) );
AND3_X1 _16770_ ( .A1(_04012_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00918_ ) );
AOI211_X1 _16771_ ( .A(_00917_ ), .B(_00918_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_06268_ ), .ZN(_00919_ ) );
NAND3_X1 _16772_ ( .A1(_00793_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00920_ ) );
NAND4_X1 _16773_ ( .A1(_00919_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_00920_ ), .ZN(_00921_ ) );
NAND3_X1 _16774_ ( .A1(_00800_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00922_ ) );
NAND3_X1 _16775_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00923_ ) );
AND2_X1 _16776_ ( .A1(_00922_ ), .A2(_00923_ ), .ZN(_00924_ ) );
NAND3_X1 _16777_ ( .A1(_04020_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00925_ ) );
NAND3_X1 _16778_ ( .A1(_00810_ ), .A2(_00792_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00926_ ) );
NAND4_X1 _16779_ ( .A1(_00924_ ), .A2(_00806_ ), .A3(_00925_ ), .A4(_00926_ ), .ZN(_00927_ ) );
AND3_X1 _16780_ ( .A1(_00921_ ), .A2(_00798_ ), .A3(_00927_ ), .ZN(_00928_ ) );
OR2_X1 _16781_ ( .A1(_00916_ ), .A2(_00928_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
AOI21_X1 _16782_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00929_ ) );
NAND2_X1 _16783_ ( .A1(_00663_ ), .A2(_00665_ ), .ZN(_00930_ ) );
OAI21_X1 _16784_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_00930_ ), .ZN(_00931_ ) );
NAND2_X1 _16785_ ( .A1(_00929_ ), .A2(_00931_ ), .ZN(_00932_ ) );
AND3_X1 _16786_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00933_ ) );
AND3_X1 _16787_ ( .A1(_04013_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00934_ ) );
AOI211_X1 _16788_ ( .A(_00933_ ), .B(_00934_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_06269_ ), .ZN(_00935_ ) );
NAND3_X1 _16789_ ( .A1(_04021_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00936_ ) );
NAND4_X1 _16790_ ( .A1(_00935_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_00936_ ), .ZN(_00937_ ) );
NAND3_X1 _16791_ ( .A1(_00869_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00938_ ) );
NAND3_X1 _16792_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00939_ ) );
AND2_X1 _16793_ ( .A1(_00938_ ), .A2(_00939_ ), .ZN(_00940_ ) );
NAND3_X1 _16794_ ( .A1(_00874_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00941_ ) );
NAND3_X1 _16795_ ( .A1(_04014_ ), .A2(_00876_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00942_ ) );
NAND4_X1 _16796_ ( .A1(_00940_ ), .A2(_00873_ ), .A3(_00941_ ), .A4(_00942_ ), .ZN(_00943_ ) );
NAND3_X1 _16797_ ( .A1(_00937_ ), .A2(_00868_ ), .A3(_00943_ ), .ZN(_00944_ ) );
NAND2_X1 _16798_ ( .A1(_00932_ ), .A2(_00944_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NAND2_X1 _16799_ ( .A1(_00666_ ), .A2(_00668_ ), .ZN(_00945_ ) );
OAI211_X1 _16800_ ( .A(_04091_ ), .B(_00818_ ), .C1(_00945_ ), .C2(_06310_ ), .ZN(_00946_ ) );
NAND2_X1 _16801_ ( .A1(_00946_ ), .A2(\myifu.state [2] ), .ZN(_00947_ ) );
AOI21_X1 _16802_ ( .A(_00947_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00883_ ), .ZN(_00948_ ) );
AND3_X1 _16803_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00949_ ) );
AND3_X1 _16804_ ( .A1(_04012_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00950_ ) );
AOI211_X1 _16805_ ( .A(_00949_ ), .B(_00950_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_06268_ ), .ZN(_00951_ ) );
NAND3_X1 _16806_ ( .A1(_00793_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00952_ ) );
NAND4_X1 _16807_ ( .A1(_00951_ ), .A2(_00787_ ), .A3(_00789_ ), .A4(_00952_ ), .ZN(_00953_ ) );
NAND3_X1 _16808_ ( .A1(_00800_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00954_ ) );
NAND3_X1 _16809_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00955_ ) );
AND2_X1 _16810_ ( .A1(_00954_ ), .A2(_00955_ ), .ZN(_00956_ ) );
NAND3_X1 _16811_ ( .A1(_04020_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00957_ ) );
NAND3_X1 _16812_ ( .A1(_04013_ ), .A2(_00792_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00958_ ) );
NAND4_X1 _16813_ ( .A1(_00956_ ), .A2(_00806_ ), .A3(_00957_ ), .A4(_00958_ ), .ZN(_00959_ ) );
AND3_X1 _16814_ ( .A1(_00953_ ), .A2(_00798_ ), .A3(_00959_ ), .ZN(_00960_ ) );
OR2_X1 _16815_ ( .A1(_00948_ ), .A2(_00960_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
OAI211_X1 _16816_ ( .A(_04091_ ), .B(_00818_ ), .C1(_00671_ ), .C2(_06310_ ), .ZN(_00961_ ) );
NAND2_X1 _16817_ ( .A1(_00961_ ), .A2(\myifu.state [2] ), .ZN(_00962_ ) );
AOI21_X1 _16818_ ( .A(_00962_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00883_ ), .ZN(_00963_ ) );
AND3_X1 _16819_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00964_ ) );
AND3_X1 _16820_ ( .A1(_04012_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00965_ ) );
AOI211_X1 _16821_ ( .A(_00964_ ), .B(_00965_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_06268_ ), .ZN(_00966_ ) );
NAND3_X1 _16822_ ( .A1(_00793_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00967_ ) );
NAND4_X1 _16823_ ( .A1(_00966_ ), .A2(_00786_ ), .A3(_00789_ ), .A4(_00967_ ), .ZN(_00968_ ) );
NAND3_X1 _16824_ ( .A1(_00800_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00969_ ) );
NAND3_X1 _16825_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00970_ ) );
AND2_X1 _16826_ ( .A1(_00969_ ), .A2(_00970_ ), .ZN(_00971_ ) );
NAND3_X1 _16827_ ( .A1(_04020_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00972_ ) );
NAND3_X1 _16828_ ( .A1(_04013_ ), .A2(_00792_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00973_ ) );
NAND4_X1 _16829_ ( .A1(_00971_ ), .A2(_00806_ ), .A3(_00972_ ), .A4(_00973_ ), .ZN(_00974_ ) );
AND3_X1 _16830_ ( .A1(_00968_ ), .A2(_00797_ ), .A3(_00974_ ), .ZN(_00975_ ) );
OR2_X1 _16831_ ( .A1(_00963_ ), .A2(_00975_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
OR2_X1 _16832_ ( .A1(_00820_ ), .A2(\myifu.data_in [14] ), .ZN(_00976_ ) );
AOI21_X1 _16833_ ( .A(_00853_ ), .B1(_00883_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00977_ ) );
NAND2_X1 _16834_ ( .A1(_00976_ ), .A2(_00977_ ), .ZN(_00978_ ) );
AND3_X1 _16835_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00979_ ) );
AND3_X1 _16836_ ( .A1(_04013_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00980_ ) );
AOI211_X1 _16837_ ( .A(_00979_ ), .B(_00980_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_06269_ ), .ZN(_00981_ ) );
NAND3_X1 _16838_ ( .A1(_04021_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00982_ ) );
NAND4_X1 _16839_ ( .A1(_00981_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_00982_ ), .ZN(_00983_ ) );
NAND3_X1 _16840_ ( .A1(_00869_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00984_ ) );
NAND3_X1 _16841_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00985_ ) );
AND2_X1 _16842_ ( .A1(_00984_ ), .A2(_00985_ ), .ZN(_00986_ ) );
BUF_X4 _16843_ ( .A(_00806_ ), .Z(_00987_ ) );
NAND3_X1 _16844_ ( .A1(_00874_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00988_ ) );
NAND3_X1 _16845_ ( .A1(_04014_ ), .A2(_00876_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00989_ ) );
NAND4_X1 _16846_ ( .A1(_00986_ ), .A2(_00987_ ), .A3(_00988_ ), .A4(_00989_ ), .ZN(_00990_ ) );
NAND3_X1 _16847_ ( .A1(_00983_ ), .A2(_00868_ ), .A3(_00990_ ), .ZN(_00991_ ) );
NAND2_X1 _16848_ ( .A1(_00978_ ), .A2(_00991_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
AOI21_X1 _16849_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00992_ ) );
NAND2_X1 _16850_ ( .A1(_00676_ ), .A2(_00678_ ), .ZN(_00993_ ) );
OAI21_X1 _16851_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_00993_ ), .ZN(_00994_ ) );
NAND2_X1 _16852_ ( .A1(_00992_ ), .A2(_00994_ ), .ZN(_00995_ ) );
AND3_X1 _16853_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00996_ ) );
CLKBUF_X2 _16854_ ( .A(_04012_ ), .Z(_00997_ ) );
AND3_X1 _16855_ ( .A1(_00997_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00998_ ) );
AOI211_X1 _16856_ ( .A(_00996_ ), .B(_00998_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_06269_ ), .ZN(_00999_ ) );
NAND3_X1 _16857_ ( .A1(_04021_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_01000_ ) );
NAND4_X1 _16858_ ( .A1(_00999_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_01000_ ), .ZN(_01001_ ) );
NAND3_X1 _16859_ ( .A1(_00869_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_01002_ ) );
NAND3_X1 _16860_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_01003_ ) );
AND2_X1 _16861_ ( .A1(_01002_ ), .A2(_01003_ ), .ZN(_01004_ ) );
NAND3_X1 _16862_ ( .A1(_00874_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_01005_ ) );
BUF_X4 _16863_ ( .A(_00810_ ), .Z(_01006_ ) );
NAND3_X1 _16864_ ( .A1(_01006_ ), .A2(_00876_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_01007_ ) );
NAND4_X1 _16865_ ( .A1(_01004_ ), .A2(_00987_ ), .A3(_01005_ ), .A4(_01007_ ), .ZN(_01008_ ) );
NAND3_X1 _16866_ ( .A1(_01001_ ), .A2(_00868_ ), .A3(_01008_ ), .ZN(_01009_ ) );
NAND2_X1 _16867_ ( .A1(_00995_ ), .A2(_01009_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
AOI21_X1 _16868_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01010_ ) );
NAND2_X1 _16869_ ( .A1(_00680_ ), .A2(_00683_ ), .ZN(_01011_ ) );
OAI21_X1 _16870_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_01011_ ), .ZN(_01012_ ) );
NAND2_X1 _16871_ ( .A1(_01010_ ), .A2(_01012_ ), .ZN(_01013_ ) );
AND3_X1 _16872_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_01014_ ) );
AND3_X1 _16873_ ( .A1(_00997_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_01015_ ) );
AOI211_X1 _16874_ ( .A(_01014_ ), .B(_01015_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_06269_ ), .ZN(_01016_ ) );
BUF_X4 _16875_ ( .A(_00793_ ), .Z(_01017_ ) );
NAND3_X1 _16876_ ( .A1(_01017_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_01018_ ) );
NAND4_X1 _16877_ ( .A1(_01016_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_01018_ ), .ZN(_01019_ ) );
NAND3_X1 _16878_ ( .A1(_00869_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_01020_ ) );
NAND3_X1 _16879_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_01021_ ) );
AND2_X1 _16880_ ( .A1(_01020_ ), .A2(_01021_ ), .ZN(_01022_ ) );
NAND3_X1 _16881_ ( .A1(_00874_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_01023_ ) );
BUF_X4 _16882_ ( .A(_04020_ ), .Z(_01024_ ) );
NAND3_X1 _16883_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_01025_ ) );
NAND4_X1 _16884_ ( .A1(_01022_ ), .A2(_00987_ ), .A3(_01023_ ), .A4(_01025_ ), .ZN(_01026_ ) );
NAND3_X1 _16885_ ( .A1(_01019_ ), .A2(_00868_ ), .A3(_01026_ ), .ZN(_01027_ ) );
NAND2_X1 _16886_ ( .A1(_01013_ ), .A2(_01027_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
AND2_X1 _16887_ ( .A1(_00685_ ), .A2(_00686_ ), .ZN(_01028_ ) );
OAI211_X1 _16888_ ( .A(_04091_ ), .B(_00818_ ), .C1(_06311_ ), .C2(_01028_ ), .ZN(_01029_ ) );
OAI211_X1 _16889_ ( .A(_01029_ ), .B(\myifu.state [2] ), .C1(_00823_ ), .C2(_03768_ ), .ZN(_01030_ ) );
AND3_X1 _16890_ ( .A1(fanout_net_15 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_01031_ ) );
AND3_X1 _16891_ ( .A1(_00997_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_01032_ ) );
AOI211_X1 _16892_ ( .A(_01031_ ), .B(_01032_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_00784_ ), .ZN(_01033_ ) );
NAND3_X1 _16893_ ( .A1(_01017_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_01034_ ) );
NAND4_X1 _16894_ ( .A1(_01033_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_01034_ ), .ZN(_01035_ ) );
NAND3_X1 _16895_ ( .A1(_00869_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_01036_ ) );
NAND3_X1 _16896_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_01037_ ) );
AND2_X1 _16897_ ( .A1(_01036_ ), .A2(_01037_ ), .ZN(_01038_ ) );
NAND3_X1 _16898_ ( .A1(_00874_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_01039_ ) );
NAND3_X1 _16899_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_01040_ ) );
NAND4_X1 _16900_ ( .A1(_01038_ ), .A2(_00987_ ), .A3(_01039_ ), .A4(_01040_ ), .ZN(_01041_ ) );
NAND3_X1 _16901_ ( .A1(_01035_ ), .A2(_00868_ ), .A3(_01041_ ), .ZN(_01042_ ) );
NAND2_X1 _16902_ ( .A1(_01030_ ), .A2(_01042_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16903_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_01043_ ) );
AND3_X1 _16904_ ( .A1(_00781_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_01044_ ) );
AOI211_X1 _16905_ ( .A(_01043_ ), .B(_01044_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_00783_ ), .ZN(_01045_ ) );
NAND3_X1 _16906_ ( .A1(_00794_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_01046_ ) );
NAND4_X1 _16907_ ( .A1(_01045_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_01046_ ), .ZN(_01047_ ) );
NAND3_X1 _16908_ ( .A1(_00801_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_01048_ ) );
NAND3_X1 _16909_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_01049_ ) );
AND2_X1 _16910_ ( .A1(_01048_ ), .A2(_01049_ ), .ZN(_01050_ ) );
NAND3_X1 _16911_ ( .A1(_00808_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_01051_ ) );
NAND3_X1 _16912_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_01052_ ) );
NAND4_X1 _16913_ ( .A1(_01050_ ), .A2(_00807_ ), .A3(_01051_ ), .A4(_01052_ ), .ZN(_01053_ ) );
NAND3_X1 _16914_ ( .A1(_01047_ ), .A2(_00799_ ), .A3(_01053_ ), .ZN(_01054_ ) );
NOR2_X1 _16915_ ( .A1(_00821_ ), .A2(\myifu.data_in [11] ), .ZN(_01055_ ) );
OAI21_X1 _16916_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03804_ ), .ZN(_01056_ ) );
OAI21_X1 _16917_ ( .A(_01054_ ), .B1(_01055_ ), .B2(_01056_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
NAND2_X1 _16918_ ( .A1(_00690_ ), .A2(_00692_ ), .ZN(_01057_ ) );
OAI211_X1 _16919_ ( .A(_04091_ ), .B(_00818_ ), .C1(_01057_ ), .C2(_06310_ ), .ZN(_01058_ ) );
NAND2_X1 _16920_ ( .A1(_01058_ ), .A2(\myifu.state [2] ), .ZN(_01059_ ) );
AOI21_X1 _16921_ ( .A(_01059_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .B2(_00883_ ), .ZN(_01060_ ) );
AND3_X1 _16922_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_01061_ ) );
AND3_X1 _16923_ ( .A1(_04012_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_01062_ ) );
AOI211_X1 _16924_ ( .A(_01061_ ), .B(_01062_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_06268_ ), .ZN(_01063_ ) );
NAND3_X1 _16925_ ( .A1(_00793_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_01064_ ) );
NAND4_X1 _16926_ ( .A1(_01063_ ), .A2(_00786_ ), .A3(_00789_ ), .A4(_01064_ ), .ZN(_01065_ ) );
NAND3_X1 _16927_ ( .A1(_00800_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_01066_ ) );
NAND3_X1 _16928_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_01067_ ) );
AND2_X1 _16929_ ( .A1(_01066_ ), .A2(_01067_ ), .ZN(_01068_ ) );
NAND3_X1 _16930_ ( .A1(_04020_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_01069_ ) );
NAND3_X1 _16931_ ( .A1(_04013_ ), .A2(_00792_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_01070_ ) );
NAND4_X1 _16932_ ( .A1(_01068_ ), .A2(_00806_ ), .A3(_01069_ ), .A4(_01070_ ), .ZN(_01071_ ) );
AND3_X1 _16933_ ( .A1(_01065_ ), .A2(_00797_ ), .A3(_01071_ ), .ZN(_01072_ ) );
OR2_X1 _16934_ ( .A1(_01060_ ), .A2(_01072_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
AOI21_X1 _16935_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_01073_ ) );
NAND2_X1 _16936_ ( .A1(_00693_ ), .A2(_00695_ ), .ZN(_01074_ ) );
OAI21_X1 _16937_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_01074_ ), .ZN(_01075_ ) );
NAND2_X1 _16938_ ( .A1(_01073_ ), .A2(_01075_ ), .ZN(_01076_ ) );
AND3_X1 _16939_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_01077_ ) );
AND3_X1 _16940_ ( .A1(_00997_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_01078_ ) );
AOI211_X1 _16941_ ( .A(_01077_ ), .B(_01078_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_00784_ ), .ZN(_01079_ ) );
NAND3_X1 _16942_ ( .A1(_01017_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_01080_ ) );
NAND4_X1 _16943_ ( .A1(_01079_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_01080_ ), .ZN(_01081_ ) );
NAND3_X1 _16944_ ( .A1(_00869_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_01082_ ) );
NAND3_X1 _16945_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_01083_ ) );
AND2_X1 _16946_ ( .A1(_01082_ ), .A2(_01083_ ), .ZN(_01084_ ) );
NAND3_X1 _16947_ ( .A1(_00874_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_01085_ ) );
NAND3_X1 _16948_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_01086_ ) );
NAND4_X1 _16949_ ( .A1(_01084_ ), .A2(_00987_ ), .A3(_01085_ ), .A4(_01086_ ), .ZN(_01087_ ) );
NAND3_X1 _16950_ ( .A1(_01081_ ), .A2(_00868_ ), .A3(_01087_ ), .ZN(_01088_ ) );
NAND2_X1 _16951_ ( .A1(_01076_ ), .A2(_01088_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
AND3_X1 _16952_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_01089_ ) );
AND3_X1 _16953_ ( .A1(_00781_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_01090_ ) );
AOI211_X1 _16954_ ( .A(_01089_ ), .B(_01090_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_00783_ ), .ZN(_01091_ ) );
NAND3_X1 _16955_ ( .A1(_00794_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_01092_ ) );
NAND4_X1 _16956_ ( .A1(_01091_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_01092_ ), .ZN(_01093_ ) );
NAND3_X1 _16957_ ( .A1(_00810_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_01094_ ) );
NAND3_X1 _16958_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_01095_ ) );
AND2_X1 _16959_ ( .A1(_01094_ ), .A2(_01095_ ), .ZN(_01096_ ) );
NAND3_X1 _16960_ ( .A1(_00808_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_01097_ ) );
NAND3_X1 _16961_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_01098_ ) );
NAND4_X1 _16962_ ( .A1(_01096_ ), .A2(_00807_ ), .A3(_01097_ ), .A4(_01098_ ), .ZN(_01099_ ) );
NAND3_X1 _16963_ ( .A1(_01093_ ), .A2(_00799_ ), .A3(_01099_ ), .ZN(_01100_ ) );
NOR2_X1 _16964_ ( .A1(_00821_ ), .A2(\myifu.data_in [7] ), .ZN(_01101_ ) );
OAI21_X1 _16965_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03759_ ), .ZN(_01102_ ) );
OAI21_X1 _16966_ ( .A(_01100_ ), .B1(_01101_ ), .B2(_01102_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AND3_X1 _16967_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_01103_ ) );
AND3_X1 _16968_ ( .A1(_00781_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_01104_ ) );
AOI211_X1 _16969_ ( .A(_01103_ ), .B(_01104_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00783_ ), .ZN(_01105_ ) );
NAND3_X1 _16970_ ( .A1(_00876_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_01106_ ) );
NAND4_X1 _16971_ ( .A1(_01105_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_01106_ ), .ZN(_01107_ ) );
NAND3_X1 _16972_ ( .A1(_00810_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_01108_ ) );
NAND3_X1 _16973_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_01109_ ) );
AND2_X1 _16974_ ( .A1(_01108_ ), .A2(_01109_ ), .ZN(_01110_ ) );
NAND3_X1 _16975_ ( .A1(_00808_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_01111_ ) );
NAND3_X1 _16976_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_01112_ ) );
NAND4_X1 _16977_ ( .A1(_01110_ ), .A2(_00807_ ), .A3(_01111_ ), .A4(_01112_ ), .ZN(_01113_ ) );
NAND3_X1 _16978_ ( .A1(_01107_ ), .A2(_00798_ ), .A3(_01113_ ), .ZN(_01114_ ) );
NOR2_X1 _16979_ ( .A1(_00821_ ), .A2(\myifu.data_in [6] ), .ZN(_01115_ ) );
OAI21_X1 _16980_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03401_ ), .ZN(_01116_ ) );
OAI21_X1 _16981_ ( .A(_01114_ ), .B1(_01115_ ), .B2(_01116_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
AOI21_X1 _16982_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01117_ ) );
OAI21_X1 _16983_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_00707_ ), .ZN(_01118_ ) );
NAND2_X1 _16984_ ( .A1(_01117_ ), .A2(_01118_ ), .ZN(_01119_ ) );
AND3_X1 _16985_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_01120_ ) );
AND3_X1 _16986_ ( .A1(_00997_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_01121_ ) );
AOI211_X1 _16987_ ( .A(_01120_ ), .B(_01121_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00784_ ), .ZN(_01122_ ) );
NAND3_X1 _16988_ ( .A1(_01017_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_01123_ ) );
NAND4_X1 _16989_ ( .A1(_01122_ ), .A2(_00864_ ), .A3(_00865_ ), .A4(_01123_ ), .ZN(_01124_ ) );
NAND3_X1 _16990_ ( .A1(_00869_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_01125_ ) );
NAND3_X1 _16991_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_01126_ ) );
AND2_X1 _16992_ ( .A1(_01125_ ), .A2(_01126_ ), .ZN(_01127_ ) );
NAND3_X1 _16993_ ( .A1(_00874_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_01128_ ) );
NAND3_X1 _16994_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_01129_ ) );
NAND4_X1 _16995_ ( .A1(_01127_ ), .A2(_00987_ ), .A3(_01128_ ), .A4(_01129_ ), .ZN(_01130_ ) );
NAND3_X1 _16996_ ( .A1(_01124_ ), .A2(_00868_ ), .A3(_01130_ ), .ZN(_01131_ ) );
NAND2_X1 _16997_ ( .A1(_01119_ ), .A2(_01131_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
AOI21_X1 _16998_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01132_ ) );
OAI21_X1 _16999_ ( .A(_00857_ ), .B1(_06345_ ), .B2(_00710_ ), .ZN(_01133_ ) );
NAND2_X1 _17000_ ( .A1(_01132_ ), .A2(_01133_ ), .ZN(_01134_ ) );
AND3_X1 _17001_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_01135_ ) );
AND3_X1 _17002_ ( .A1(_00997_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_01136_ ) );
AOI211_X1 _17003_ ( .A(_01135_ ), .B(_01136_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00784_ ), .ZN(_01137_ ) );
NAND3_X1 _17004_ ( .A1(_01017_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_01138_ ) );
NAND4_X1 _17005_ ( .A1(_01137_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_01138_ ), .ZN(_01139_ ) );
NAND3_X1 _17006_ ( .A1(_00801_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_01140_ ) );
NAND3_X1 _17007_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_01141_ ) );
AND2_X1 _17008_ ( .A1(_01140_ ), .A2(_01141_ ), .ZN(_01142_ ) );
NAND3_X1 _17009_ ( .A1(_00874_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_01143_ ) );
NAND3_X1 _17010_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_01144_ ) );
NAND4_X1 _17011_ ( .A1(_01142_ ), .A2(_00987_ ), .A3(_01143_ ), .A4(_01144_ ), .ZN(_01145_ ) );
NAND3_X1 _17012_ ( .A1(_01139_ ), .A2(_00868_ ), .A3(_01145_ ), .ZN(_01146_ ) );
NAND2_X1 _17013_ ( .A1(_01134_ ), .A2(_01146_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _17014_ ( .A(_00854_ ), .B1(_00855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01147_ ) );
OAI21_X1 _17015_ ( .A(_00857_ ), .B1(_06311_ ), .B2(_00713_ ), .ZN(_01148_ ) );
NAND2_X1 _17016_ ( .A1(_01147_ ), .A2(_01148_ ), .ZN(_01149_ ) );
AND3_X1 _17017_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_01150_ ) );
AND3_X1 _17018_ ( .A1(_00997_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_01151_ ) );
AOI211_X1 _17019_ ( .A(_01150_ ), .B(_01151_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00784_ ), .ZN(_01152_ ) );
NAND3_X1 _17020_ ( .A1(_01017_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_01153_ ) );
NAND4_X1 _17021_ ( .A1(_01152_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_01153_ ), .ZN(_01154_ ) );
NAND3_X1 _17022_ ( .A1(_00801_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_01155_ ) );
NAND3_X1 _17023_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_01156_ ) );
AND2_X1 _17024_ ( .A1(_01155_ ), .A2(_01156_ ), .ZN(_01157_ ) );
NAND3_X1 _17025_ ( .A1(_00794_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_01158_ ) );
NAND3_X1 _17026_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_01159_ ) );
NAND4_X1 _17027_ ( .A1(_01157_ ), .A2(_00987_ ), .A3(_01158_ ), .A4(_01159_ ), .ZN(_01160_ ) );
NAND3_X1 _17028_ ( .A1(_01154_ ), .A2(_00799_ ), .A3(_01160_ ), .ZN(_01161_ ) );
NAND2_X1 _17029_ ( .A1(_01149_ ), .A2(_01161_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
AOI21_X1 _17030_ ( .A(_00854_ ), .B1(_00883_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01162_ ) );
OAI21_X1 _17031_ ( .A(_00819_ ), .B1(_06311_ ), .B2(_00716_ ), .ZN(_01163_ ) );
NAND2_X1 _17032_ ( .A1(_01162_ ), .A2(_01163_ ), .ZN(_01164_ ) );
AND3_X1 _17033_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_01165_ ) );
AND3_X1 _17034_ ( .A1(_00997_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_01166_ ) );
AOI211_X1 _17035_ ( .A(_01165_ ), .B(_01166_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_00784_ ), .ZN(_01167_ ) );
NAND3_X1 _17036_ ( .A1(_01017_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_01168_ ) );
NAND4_X1 _17037_ ( .A1(_01167_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_01168_ ), .ZN(_01169_ ) );
NAND3_X1 _17038_ ( .A1(_00801_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_01170_ ) );
NAND3_X1 _17039_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_01171_ ) );
AND2_X1 _17040_ ( .A1(_01170_ ), .A2(_01171_ ), .ZN(_01172_ ) );
NAND3_X1 _17041_ ( .A1(_00794_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_01173_ ) );
NAND3_X1 _17042_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_01174_ ) );
NAND4_X1 _17043_ ( .A1(_01172_ ), .A2(_00987_ ), .A3(_01173_ ), .A4(_01174_ ), .ZN(_01175_ ) );
NAND3_X1 _17044_ ( .A1(_01169_ ), .A2(_00799_ ), .A3(_01175_ ), .ZN(_01176_ ) );
NAND2_X1 _17045_ ( .A1(_01164_ ), .A2(_01176_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
AOI21_X1 _17046_ ( .A(_00853_ ), .B1(_00883_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01177_ ) );
OAI21_X1 _17047_ ( .A(_00819_ ), .B1(_06311_ ), .B2(_00722_ ), .ZN(_01178_ ) );
NAND2_X1 _17048_ ( .A1(_01177_ ), .A2(_01178_ ), .ZN(_01179_ ) );
AND3_X1 _17049_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01180_ ) );
AND3_X1 _17050_ ( .A1(_00997_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01181_ ) );
AOI211_X1 _17051_ ( .A(_01180_ ), .B(_01181_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_00784_ ), .ZN(_01182_ ) );
NAND3_X1 _17052_ ( .A1(_01017_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01183_ ) );
NAND4_X1 _17053_ ( .A1(_01182_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_01183_ ), .ZN(_01184_ ) );
NAND3_X1 _17054_ ( .A1(_00801_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01185_ ) );
NAND3_X1 _17055_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01186_ ) );
AND2_X1 _17056_ ( .A1(_01185_ ), .A2(_01186_ ), .ZN(_01187_ ) );
NAND3_X1 _17057_ ( .A1(_00794_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01188_ ) );
NAND3_X1 _17058_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01189_ ) );
NAND4_X1 _17059_ ( .A1(_01187_ ), .A2(_00987_ ), .A3(_01188_ ), .A4(_01189_ ), .ZN(_01190_ ) );
NAND3_X1 _17060_ ( .A1(_01184_ ), .A2(_00799_ ), .A3(_01190_ ), .ZN(_01191_ ) );
NAND2_X1 _17061_ ( .A1(_01179_ ), .A2(_01191_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
AND3_X1 _17062_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01192_ ) );
AND3_X1 _17063_ ( .A1(_00781_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01193_ ) );
AOI211_X1 _17064_ ( .A(_01192_ ), .B(_01193_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00783_ ), .ZN(_01194_ ) );
NAND3_X1 _17065_ ( .A1(_00876_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01195_ ) );
NAND4_X1 _17066_ ( .A1(_01194_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_01195_ ), .ZN(_01196_ ) );
NAND3_X1 _17067_ ( .A1(_00810_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01197_ ) );
NAND3_X1 _17068_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01198_ ) );
AND2_X1 _17069_ ( .A1(_01197_ ), .A2(_01198_ ), .ZN(_01199_ ) );
NAND3_X1 _17070_ ( .A1(_00808_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01200_ ) );
NAND3_X1 _17071_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01201_ ) );
NAND4_X1 _17072_ ( .A1(_01199_ ), .A2(_00807_ ), .A3(_01200_ ), .A4(_01201_ ), .ZN(_01202_ ) );
NAND3_X1 _17073_ ( .A1(_01196_ ), .A2(_00798_ ), .A3(_01202_ ), .ZN(_01203_ ) );
NOR2_X1 _17074_ ( .A1(_00821_ ), .A2(\myifu.data_in [28] ), .ZN(_01204_ ) );
OAI21_X1 _17075_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03825_ ), .ZN(_01205_ ) );
OAI21_X1 _17076_ ( .A(_01203_ ), .B1(_01204_ ), .B2(_01205_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
OAI211_X1 _17077_ ( .A(_04091_ ), .B(_00818_ ), .C1(_00725_ ), .C2(_06310_ ), .ZN(_01206_ ) );
NAND2_X1 _17078_ ( .A1(_01206_ ), .A2(\myifu.state [2] ), .ZN(_01207_ ) );
AOI21_X1 _17079_ ( .A(_01207_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00883_ ), .ZN(_01208_ ) );
AND3_X1 _17080_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01209_ ) );
AND3_X1 _17081_ ( .A1(_04012_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01210_ ) );
AOI211_X1 _17082_ ( .A(_01209_ ), .B(_01210_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_06268_ ), .ZN(_01211_ ) );
NAND3_X1 _17083_ ( .A1(_00793_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01212_ ) );
NAND4_X1 _17084_ ( .A1(_01211_ ), .A2(_00786_ ), .A3(_00789_ ), .A4(_01212_ ), .ZN(_01213_ ) );
NAND3_X1 _17085_ ( .A1(_00800_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01214_ ) );
NAND3_X1 _17086_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01215_ ) );
AND2_X1 _17087_ ( .A1(_01214_ ), .A2(_01215_ ), .ZN(_01216_ ) );
NAND3_X1 _17088_ ( .A1(_04020_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01217_ ) );
NAND3_X1 _17089_ ( .A1(_04013_ ), .A2(_00792_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01218_ ) );
NAND4_X1 _17090_ ( .A1(_01216_ ), .A2(_00806_ ), .A3(_01217_ ), .A4(_01218_ ), .ZN(_01219_ ) );
AND3_X1 _17091_ ( .A1(_01213_ ), .A2(_00797_ ), .A3(_01219_ ), .ZN(_01220_ ) );
OR2_X1 _17092_ ( .A1(_01208_ ), .A2(_01220_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
AND2_X1 _17093_ ( .A1(_00727_ ), .A2(_00728_ ), .ZN(_01221_ ) );
OAI211_X1 _17094_ ( .A(_04091_ ), .B(_00818_ ), .C1(_06311_ ), .C2(_01221_ ), .ZN(_01222_ ) );
OAI211_X1 _17095_ ( .A(_01222_ ), .B(\myifu.state [2] ), .C1(_00823_ ), .C2(_03817_ ), .ZN(_01223_ ) );
AND3_X1 _17096_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01224_ ) );
AND3_X1 _17097_ ( .A1(_00997_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01225_ ) );
AOI211_X1 _17098_ ( .A(_01224_ ), .B(_01225_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00784_ ), .ZN(_01226_ ) );
NAND3_X1 _17099_ ( .A1(_01017_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01227_ ) );
NAND4_X1 _17100_ ( .A1(_01226_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_01227_ ), .ZN(_01228_ ) );
NAND3_X1 _17101_ ( .A1(_00801_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01229_ ) );
NAND3_X1 _17102_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01230_ ) );
AND2_X1 _17103_ ( .A1(_01229_ ), .A2(_01230_ ), .ZN(_01231_ ) );
NAND3_X1 _17104_ ( .A1(_00794_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01232_ ) );
NAND3_X1 _17105_ ( .A1(_01006_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01233_ ) );
NAND4_X1 _17106_ ( .A1(_01231_ ), .A2(_00807_ ), .A3(_01232_ ), .A4(_01233_ ), .ZN(_01234_ ) );
NAND3_X1 _17107_ ( .A1(_01228_ ), .A2(_00799_ ), .A3(_01234_ ), .ZN(_01235_ ) );
NAND2_X1 _17108_ ( .A1(_01223_ ), .A2(_01235_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
AND3_X1 _17109_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01236_ ) );
AND3_X1 _17110_ ( .A1(_00781_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01237_ ) );
AOI211_X1 _17111_ ( .A(_01236_ ), .B(_01237_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_00783_ ), .ZN(_01238_ ) );
NAND3_X1 _17112_ ( .A1(_00876_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01239_ ) );
NAND4_X1 _17113_ ( .A1(_01238_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_01239_ ), .ZN(_01240_ ) );
NAND3_X1 _17114_ ( .A1(_00810_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01241_ ) );
NAND3_X1 _17115_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01242_ ) );
AND2_X1 _17116_ ( .A1(_01241_ ), .A2(_01242_ ), .ZN(_01243_ ) );
NAND3_X1 _17117_ ( .A1(_00808_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01244_ ) );
NAND3_X1 _17118_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01245_ ) );
NAND4_X1 _17119_ ( .A1(_01243_ ), .A2(_00807_ ), .A3(_01244_ ), .A4(_01245_ ), .ZN(_01246_ ) );
NAND3_X1 _17120_ ( .A1(_01240_ ), .A2(_00798_ ), .A3(_01246_ ), .ZN(_01247_ ) );
NOR2_X1 _17121_ ( .A1(_00821_ ), .A2(\myifu.data_in [26] ), .ZN(_01248_ ) );
OAI21_X1 _17122_ ( .A(\myifu.state [2] ), .B1(_00823_ ), .B2(_03811_ ), .ZN(_01249_ ) );
OAI21_X1 _17123_ ( .A(_01247_ ), .B1(_01248_ ), .B2(_01249_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
AND3_X1 _17124_ ( .A1(\IF_ID_pc [4] ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01250_ ) );
AND3_X1 _17125_ ( .A1(_00781_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01251_ ) );
AOI211_X1 _17126_ ( .A(_01250_ ), .B(_01251_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00783_ ), .ZN(_01252_ ) );
NAND3_X1 _17127_ ( .A1(_00876_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01253_ ) );
NAND4_X1 _17128_ ( .A1(_01252_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_01253_ ), .ZN(_01254_ ) );
NAND3_X1 _17129_ ( .A1(_00810_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01255_ ) );
NAND3_X1 _17130_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01256_ ) );
AND2_X1 _17131_ ( .A1(_01255_ ), .A2(_01256_ ), .ZN(_01257_ ) );
NAND3_X1 _17132_ ( .A1(_00808_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01258_ ) );
NAND3_X1 _17133_ ( .A1(_00811_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01259_ ) );
NAND4_X1 _17134_ ( .A1(_01257_ ), .A2(_00806_ ), .A3(_01258_ ), .A4(_01259_ ), .ZN(_01260_ ) );
NAND3_X1 _17135_ ( .A1(_01254_ ), .A2(_00798_ ), .A3(_01260_ ), .ZN(_01261_ ) );
NOR2_X1 _17136_ ( .A1(_00821_ ), .A2(\myifu.data_in [25] ), .ZN(_01262_ ) );
OAI21_X1 _17137_ ( .A(\myifu.state [2] ), .B1(_00857_ ), .B2(_03779_ ), .ZN(_01263_ ) );
OAI21_X1 _17138_ ( .A(_01261_ ), .B1(_01262_ ), .B2(_01263_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
AND3_X1 _17139_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01264_ ) );
AND3_X1 _17140_ ( .A1(_00800_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01265_ ) );
AOI211_X1 _17141_ ( .A(_01264_ ), .B(_01265_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_00783_ ), .ZN(_01266_ ) );
NAND3_X1 _17142_ ( .A1(_00876_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01267_ ) );
NAND4_X1 _17143_ ( .A1(_01266_ ), .A2(_00787_ ), .A3(_00790_ ), .A4(_01267_ ), .ZN(_01268_ ) );
NAND3_X1 _17144_ ( .A1(_00810_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01269_ ) );
NAND3_X1 _17145_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01270_ ) );
AND2_X1 _17146_ ( .A1(_01269_ ), .A2(_01270_ ), .ZN(_01271_ ) );
NAND3_X1 _17147_ ( .A1(_00808_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01272_ ) );
NAND3_X1 _17148_ ( .A1(_00869_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01273_ ) );
NAND4_X1 _17149_ ( .A1(_01271_ ), .A2(_00806_ ), .A3(_01272_ ), .A4(_01273_ ), .ZN(_01274_ ) );
NAND3_X1 _17150_ ( .A1(_01268_ ), .A2(_00798_ ), .A3(_01274_ ), .ZN(_01275_ ) );
AND2_X1 _17151_ ( .A1(_00855_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01276_ ) );
OAI21_X1 _17152_ ( .A(\myifu.state [2] ), .B1(_00821_ ), .B2(\myifu.data_in [24] ), .ZN(_01277_ ) );
OAI21_X1 _17153_ ( .A(_01275_ ), .B1(_01276_ ), .B2(_01277_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
AOI21_X1 _17154_ ( .A(_00853_ ), .B1(_00883_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01278_ ) );
OAI21_X1 _17155_ ( .A(_00819_ ), .B1(_06311_ ), .B2(_00740_ ), .ZN(_01279_ ) );
NAND2_X1 _17156_ ( .A1(_01278_ ), .A2(_01279_ ), .ZN(_01280_ ) );
AND3_X1 _17157_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01281_ ) );
AND3_X1 _17158_ ( .A1(_00781_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01282_ ) );
AOI211_X1 _17159_ ( .A(_01281_ ), .B(_01282_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_00784_ ), .ZN(_01283_ ) );
NAND3_X1 _17160_ ( .A1(_01017_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01284_ ) );
NAND4_X1 _17161_ ( .A1(_01283_ ), .A2(_00788_ ), .A3(_00791_ ), .A4(_01284_ ), .ZN(_01285_ ) );
NAND3_X1 _17162_ ( .A1(_00801_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01286_ ) );
NAND3_X1 _17163_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01287_ ) );
AND2_X1 _17164_ ( .A1(_01286_ ), .A2(_01287_ ), .ZN(_01288_ ) );
NAND3_X1 _17165_ ( .A1(_00794_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01289_ ) );
NAND3_X1 _17166_ ( .A1(_00811_ ), .A2(_01024_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01290_ ) );
NAND4_X1 _17167_ ( .A1(_01288_ ), .A2(_00807_ ), .A3(_01289_ ), .A4(_01290_ ), .ZN(_01291_ ) );
NAND3_X1 _17168_ ( .A1(_01285_ ), .A2(_00799_ ), .A3(_01291_ ), .ZN(_01292_ ) );
NAND2_X1 _17169_ ( .A1(_01280_ ), .A2(_01292_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
OAI211_X1 _17170_ ( .A(_04091_ ), .B(_00818_ ), .C1(_00743_ ), .C2(_02167_ ), .ZN(_01293_ ) );
NAND2_X1 _17171_ ( .A1(_01293_ ), .A2(\myifu.state [2] ), .ZN(_01294_ ) );
AOI21_X1 _17172_ ( .A(_01294_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .B2(_00820_ ), .ZN(_01295_ ) );
AND3_X1 _17173_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01296_ ) );
AND3_X1 _17174_ ( .A1(_04012_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01297_ ) );
AOI211_X1 _17175_ ( .A(_01296_ ), .B(_01297_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_06268_ ), .ZN(_01298_ ) );
NAND3_X1 _17176_ ( .A1(_00793_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01299_ ) );
NAND4_X1 _17177_ ( .A1(_01298_ ), .A2(_00786_ ), .A3(_00789_ ), .A4(_01299_ ), .ZN(_01300_ ) );
NAND3_X1 _17178_ ( .A1(_00800_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01301_ ) );
NAND3_X1 _17179_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01302_ ) );
AND2_X1 _17180_ ( .A1(_01301_ ), .A2(_01302_ ), .ZN(_01303_ ) );
NAND3_X1 _17181_ ( .A1(_00792_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01304_ ) );
NAND3_X1 _17182_ ( .A1(_04013_ ), .A2(_00792_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01305_ ) );
NAND4_X1 _17183_ ( .A1(_01303_ ), .A2(_00805_ ), .A3(_01304_ ), .A4(_01305_ ), .ZN(_01306_ ) );
AND3_X1 _17184_ ( .A1(_01300_ ), .A2(_00797_ ), .A3(_01306_ ), .ZN(_01307_ ) );
OR2_X1 _17185_ ( .A1(_01295_ ), .A2(_01307_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI211_X1 _17186_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_03539_ ), .C1(_03913_ ), .C2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _17187_ ( .A1(_04086_ ), .A2(_04089_ ), .A3(\myifu.state [2] ), .A4(_04092_ ), .ZN(_01308_ ) );
INV_X1 _17188_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01309_ ) );
AND4_X1 _17189_ ( .A1(_01309_ ), .A2(_02052_ ), .A3(\myifu.state [0] ), .A4(_02137_ ), .ZN(_01310_ ) );
NOR2_X1 _17190_ ( .A1(_01310_ ), .A2(_00637_ ), .ZN(_01311_ ) );
AOI21_X1 _17191_ ( .A(reset ), .B1(_01308_ ), .B2(_01311_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _17192_ ( .A1(_06258_ ), .A2(_02167_ ), .ZN(_01312_ ) );
INV_X1 _17193_ ( .A(_01312_ ), .ZN(_01313_ ) );
AND3_X1 _17194_ ( .A1(_01313_ ), .A2(_01309_ ), .A3(_02156_ ), .ZN(_01314_ ) );
AND2_X1 _17195_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01315_ ) );
OR4_X1 _17196_ ( .A1(reset ), .A2(_01314_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A4(_01315_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _17197_ ( .A1(_04094_ ), .A2(_01813_ ), .A3(\myifu.state [2] ), .ZN(_01316_ ) );
NAND2_X1 _17198_ ( .A1(_01312_ ), .A2(_02269_ ), .ZN(_01317_ ) );
NAND2_X1 _17199_ ( .A1(_01316_ ), .A2(_01317_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _17200_ ( .A1(_04086_ ), .A2(\myifu.state [2] ), .A3(_04089_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17201_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01318_ ) );
NOR3_X1 _17202_ ( .A1(_01318_ ), .A2(_00747_ ), .A3(_00873_ ), .ZN(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ) );
NOR3_X1 _17203_ ( .A1(_01318_ ), .A2(_00748_ ), .A3(_00873_ ), .ZN(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ) );
AND4_X1 _17204_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00873_ ), .ZN(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ) );
AND4_X1 _17205_ ( .A1(\IF_ID_pc [4] ), .A2(_06267_ ), .A3(_04021_ ), .A4(_00873_ ), .ZN(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ) );
NOR3_X1 _17206_ ( .A1(_01318_ ), .A2(_00745_ ), .A3(_00873_ ), .ZN(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ) );
AND4_X1 _17207_ ( .A1(_04014_ ), .A2(_06267_ ), .A3(\IF_ID_pc [3] ), .A4(_00873_ ), .ZN(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _17208_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06269_ ), .A3(_00873_ ), .ZN(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ) );
AND4_X1 _17209_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06269_ ), .A3(_00864_ ), .A4(_00865_ ), .ZN(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ) );
AND3_X1 _17210_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_04014_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ) );
AND3_X1 _17211_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_04021_ ), .ZN(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ) );
AND3_X1 _17212_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _17213_ ( .A1(_02268_ ), .A2(_06269_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ) );
AND2_X1 _17214_ ( .A1(_02138_ ), .A2(\myifu.state [0] ), .ZN(_01319_ ) );
AOI21_X1 _17215_ ( .A(_03539_ ), .B1(IDU_ready_IFU ), .B2(\myifu.to_reset ), .ZN(_01320_ ) );
AND2_X1 _17216_ ( .A1(_00639_ ), .A2(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01321_ ) );
OR4_X1 _17217_ ( .A1(_01319_ ), .A2(_01315_ ), .A3(_01320_ ), .A4(_01321_ ), .ZN(_01322_ ) );
AOI221_X1 _17218_ ( .A(_01322_ ), .B1(\myifu.state [0] ), .B2(_01313_ ), .C1(_04094_ ), .C2(_02191_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17219_ ( .A1(_03959_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03541_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17220_ ( .A(_03378_ ), .ZN(_01323_ ) );
AOI211_X1 _17221_ ( .A(_03617_ ), .B(_00621_ ), .C1(_03318_ ), .C2(_01323_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
OR4_X1 _17222_ ( .A1(reset ), .A2(_01321_ ), .A3(_01315_ ), .A4(_01320_ ), .ZN(_01324_ ) );
AOI21_X1 _17223_ ( .A(_01324_ ), .B1(_02139_ ), .B2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _17224_ ( .A(_06272_ ), .B(_04156_ ), .S(\mylsu.state [0] ), .Z(_01325_ ) );
NOR2_X1 _17225_ ( .A1(_06358_ ), .A2(_01325_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ) );
NOR3_X1 _17226_ ( .A1(_06358_ ), .A2(_04159_ ), .A3(_01325_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
AND2_X1 _17227_ ( .A1(_06357_ ), .A2(_04089_ ), .ZN(_01326_ ) );
AND2_X1 _17228_ ( .A1(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .A2(_03320_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
AND3_X1 _17229_ ( .A1(_02253_ ), .A2(_02244_ ), .A3(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .ZN(_01327_ ) );
INV_X1 _17230_ ( .A(_01327_ ), .ZN(_01328_ ) );
OAI22_X1 _17231_ ( .A1(_01326_ ), .A2(_06294_ ), .B1(_06261_ ), .B2(_01328_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _17232_ ( .A(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .B(_03338_ ), .C1(io_master_wready ), .C2(io_master_awready ), .ZN(_01329_ ) );
NOR4_X1 _17233_ ( .A1(_02264_ ), .A2(_02251_ ), .A3(_04100_ ), .A4(_01329_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
AND2_X1 _17234_ ( .A1(_02265_ ), .A2(\mylsu.state [0] ), .ZN(_01330_ ) );
AND2_X1 _17235_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01331_ ) );
NOR3_X1 _17236_ ( .A1(_06264_ ), .A2(_04109_ ), .A3(_01331_ ), .ZN(_01332_ ) );
NAND4_X1 _17237_ ( .A1(_01330_ ), .A2(io_master_awready ), .A3(_02256_ ), .A4(_01332_ ), .ZN(_01333_ ) );
OR4_X1 _17238_ ( .A1(reset ), .A2(_06353_ ), .A3(excp_written ), .A4(io_master_wready ), .ZN(_01334_ ) );
NAND2_X1 _17239_ ( .A1(_01333_ ), .A2(_01334_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
NAND4_X1 _17240_ ( .A1(_01330_ ), .A2(_06276_ ), .A3(_02256_ ), .A4(_01331_ ), .ZN(_01335_ ) );
AOI221_X4 _17241_ ( .A(_06365_ ), .B1(\mylsu.state [2] ), .B2(io_master_wready ), .C1(\mylsu.state [4] ), .C2(io_master_awready ), .ZN(_01336_ ) );
AOI21_X1 _17242_ ( .A(_04142_ ), .B1(_01335_ ), .B2(_01336_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
AND4_X1 _17243_ ( .A1(_02244_ ), .A2(_06288_ ), .A3(_02251_ ), .A4(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .ZN(_01337_ ) );
AOI21_X1 _17244_ ( .A(_01337_ ), .B1(_06261_ ), .B2(_01327_ ), .ZN(_01338_ ) );
NOR4_X1 _17245_ ( .A1(_06264_ ), .A2(_04109_ ), .A3(io_master_wready ), .A4(io_master_awready ), .ZN(_01339_ ) );
NAND3_X1 _17246_ ( .A1(_01330_ ), .A2(_02256_ ), .A3(_01339_ ), .ZN(_01340_ ) );
INV_X1 _17247_ ( .A(\mylsu.state [0] ), .ZN(_01341_ ) );
NAND4_X1 _17248_ ( .A1(_04100_ ), .A2(_04132_ ), .A3(_06292_ ), .A4(_06263_ ), .ZN(_01342_ ) );
OAI211_X1 _17249_ ( .A(_01338_ ), .B(_01340_ ), .C1(_01341_ ), .C2(_01342_ ), .ZN(_01343_ ) );
AND2_X1 _17250_ ( .A1(_02257_ ), .A2(_06287_ ), .ZN(_01344_ ) );
AND3_X1 _17251_ ( .A1(_02255_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A3(_03320_ ), .ZN(_01345_ ) );
NAND4_X1 _17252_ ( .A1(_01344_ ), .A2(_06276_ ), .A3(_06292_ ), .A4(_01345_ ), .ZN(_01346_ ) );
NAND4_X1 _17253_ ( .A1(_02242_ ), .A2(_02245_ ), .A3(_04112_ ), .A4(_06263_ ), .ZN(_01347_ ) );
AOI21_X1 _17254_ ( .A(_01341_ ), .B1(_01346_ ), .B2(_01347_ ), .ZN(_01348_ ) );
NAND4_X1 _17255_ ( .A1(_06357_ ), .A2(_04089_ ), .A3(\mylsu.state [3] ), .A4(_03338_ ), .ZN(_01349_ ) );
NAND3_X1 _17256_ ( .A1(_06364_ ), .A2(\mylsu.state [1] ), .A3(_03338_ ), .ZN(_01350_ ) );
NAND2_X1 _17257_ ( .A1(_01349_ ), .A2(_01350_ ), .ZN(_01351_ ) );
AND4_X1 _17258_ ( .A1(_06276_ ), .A2(_02264_ ), .A3(_06292_ ), .A4(_01345_ ), .ZN(_01352_ ) );
NAND2_X1 _17259_ ( .A1(_01352_ ), .A2(\mylsu.state [0] ), .ZN(_01353_ ) );
NAND2_X1 _17260_ ( .A1(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .A2(_04109_ ), .ZN(_01354_ ) );
NAND3_X1 _17261_ ( .A1(_03320_ ), .A2(\mylsu.state [0] ), .A3(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01355_ ) );
NAND4_X1 _17262_ ( .A1(_01353_ ), .A2(_03338_ ), .A3(_01354_ ), .A4(_01355_ ), .ZN(_01356_ ) );
OR4_X1 _17263_ ( .A1(_01343_ ), .A2(_01348_ ), .A3(_01351_ ), .A4(_01356_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND3_X1 _17264_ ( .A1(_06248_ ), .A2(\mylsu.state [0] ), .A3(io_master_wready ), .ZN(_01357_ ) );
NOR4_X1 _17265_ ( .A1(_06249_ ), .A2(_04109_ ), .A3(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A4(_01357_ ), .ZN(_01358_ ) );
NAND3_X1 _17266_ ( .A1(_02265_ ), .A2(_04158_ ), .A3(_01358_ ), .ZN(_01359_ ) );
NAND3_X1 _17267_ ( .A1(_04158_ ), .A2(\mylsu.state [4] ), .A3(_06248_ ), .ZN(_01360_ ) );
NAND2_X1 _17268_ ( .A1(_01359_ ), .A2(_01360_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
MUX2_X1 _17269_ ( .A(\LS_WB_wdata_csreg [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_04105_ ), .Z(_01361_ ) );
INV_X2 _17270_ ( .A(_04110_ ), .ZN(_01362_ ) );
OR2_X1 _17271_ ( .A1(_04101_ ), .A2(_01362_ ), .ZN(_01363_ ) );
BUF_X4 _17272_ ( .A(_01363_ ), .Z(_01364_ ) );
BUF_X4 _17273_ ( .A(_01364_ ), .Z(_01365_ ) );
MUX2_X1 _17274_ ( .A(_01361_ ), .B(\EX_LS_pc [21] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
AOI21_X1 _17275_ ( .A(\EX_LS_pc [20] ), .B1(_04103_ ), .B2(_04111_ ), .ZN(_01366_ ) );
MUX2_X1 _17276_ ( .A(\LS_WB_wdata_csreg [20] ), .B(\EX_LS_result_csreg_mem [20] ), .S(_04105_ ), .Z(_01367_ ) );
NOR3_X1 _17277_ ( .A1(_06279_ ), .A2(_01362_ ), .A3(_01367_ ), .ZN(_01368_ ) );
NOR2_X1 _17278_ ( .A1(_01366_ ), .A2(_01368_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
AOI21_X1 _17279_ ( .A(\EX_LS_pc [19] ), .B1(_04103_ ), .B2(_04111_ ), .ZN(_01369_ ) );
MUX2_X1 _17280_ ( .A(\LS_WB_wdata_csreg [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_04105_ ), .Z(_01370_ ) );
NOR3_X1 _17281_ ( .A1(_06279_ ), .A2(_01362_ ), .A3(_01370_ ), .ZN(_01371_ ) );
NOR2_X1 _17282_ ( .A1(_01369_ ), .A2(_01371_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _17283_ ( .A(\LS_WB_wdata_csreg [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_04105_ ), .Z(_01372_ ) );
MUX2_X1 _17284_ ( .A(_01372_ ), .B(\EX_LS_pc [18] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
OAI22_X1 _17285_ ( .A1(_06295_ ), .A2(_02281_ ), .B1(_04117_ ), .B2(_06397_ ), .ZN(_01373_ ) );
MUX2_X1 _17286_ ( .A(_01373_ ), .B(\EX_LS_pc [17] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _17287_ ( .A(\EX_LS_pc [16] ), .B1(_04103_ ), .B2(_04111_ ), .ZN(_01374_ ) );
MUX2_X1 _17288_ ( .A(\LS_WB_wdata_csreg [16] ), .B(\EX_LS_result_csreg_mem [16] ), .S(_04105_ ), .Z(_01375_ ) );
NOR3_X1 _17289_ ( .A1(_06279_ ), .A2(_01362_ ), .A3(_01375_ ), .ZN(_01376_ ) );
NOR2_X1 _17290_ ( .A1(_01374_ ), .A2(_01376_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
AOI21_X1 _17291_ ( .A(\EX_LS_pc [15] ), .B1(_04103_ ), .B2(_04111_ ), .ZN(_01377_ ) );
BUF_X4 _17292_ ( .A(_04110_ ), .Z(_01378_ ) );
NAND3_X1 _17293_ ( .A1(_04115_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_result_csreg_mem [15] ), .ZN(_01379_ ) );
OAI211_X1 _17294_ ( .A(_01378_ ), .B(_01379_ ), .C1(_02283_ ), .C2(_06295_ ), .ZN(_01380_ ) );
NOR2_X1 _17295_ ( .A1(_06279_ ), .A2(_01380_ ), .ZN(_01381_ ) );
NOR2_X1 _17296_ ( .A1(_01377_ ), .A2(_01381_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _17297_ ( .A(\EX_LS_pc [14] ), .B1(_04103_ ), .B2(_04111_ ), .ZN(_01382_ ) );
MUX2_X1 _17298_ ( .A(\LS_WB_wdata_csreg [14] ), .B(\EX_LS_result_csreg_mem [14] ), .S(_04105_ ), .Z(_01383_ ) );
NOR3_X1 _17299_ ( .A1(_06279_ ), .A2(_01362_ ), .A3(_01383_ ), .ZN(_01384_ ) );
NOR2_X1 _17300_ ( .A1(_01382_ ), .A2(_01384_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
BUF_X4 _17301_ ( .A(_04102_ ), .Z(_01385_ ) );
AOI21_X1 _17302_ ( .A(\EX_LS_pc [13] ), .B1(_01385_ ), .B2(_04111_ ), .ZN(_01386_ ) );
NAND3_X1 _17303_ ( .A1(_04115_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_result_csreg_mem [13] ), .ZN(_01387_ ) );
OAI211_X1 _17304_ ( .A(_01378_ ), .B(_01387_ ), .C1(_02285_ ), .C2(_06295_ ), .ZN(_01388_ ) );
NOR2_X1 _17305_ ( .A1(_06279_ ), .A2(_01388_ ), .ZN(_01389_ ) );
NOR2_X1 _17306_ ( .A1(_01386_ ), .A2(_01389_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
INV_X1 _17307_ ( .A(_04104_ ), .ZN(_01390_ ) );
BUF_X4 _17308_ ( .A(_01390_ ), .Z(_01391_ ) );
AOI221_X4 _17309_ ( .A(_01365_ ), .B1(\LS_WB_wdata_csreg [12] ), .B2(_01391_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [12] ), .ZN(_01392_ ) );
BUF_X4 _17310_ ( .A(_04110_ ), .Z(_01393_ ) );
AOI21_X1 _17311_ ( .A(\EX_LS_pc [12] ), .B1(_01385_ ), .B2(_01393_ ), .ZN(_01394_ ) );
NOR2_X1 _17312_ ( .A1(_01392_ ), .A2(_01394_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI221_X4 _17313_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [30] ), .B2(_01391_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [30] ), .ZN(_01395_ ) );
AOI21_X1 _17314_ ( .A(\EX_LS_pc [30] ), .B1(_01385_ ), .B2(_01393_ ), .ZN(_01396_ ) );
NOR2_X1 _17315_ ( .A1(_01395_ ), .A2(_01396_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
AOI221_X4 _17316_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [11] ), .B2(_01391_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [11] ), .ZN(_01397_ ) );
AOI21_X1 _17317_ ( .A(\EX_LS_pc [11] ), .B1(_01385_ ), .B2(_01393_ ), .ZN(_01398_ ) );
NOR2_X1 _17318_ ( .A1(_01397_ ), .A2(_01398_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _17319_ ( .A(\EX_LS_pc [10] ), .B1(_01385_ ), .B2(_04111_ ), .ZN(_01399_ ) );
MUX2_X1 _17320_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_04105_ ), .Z(_01400_ ) );
NOR3_X1 _17321_ ( .A1(_06279_ ), .A2(_01362_ ), .A3(_01400_ ), .ZN(_01401_ ) );
NOR2_X1 _17322_ ( .A1(_01399_ ), .A2(_01401_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
AOI21_X1 _17323_ ( .A(\EX_LS_pc [9] ), .B1(_01385_ ), .B2(_04111_ ), .ZN(_01402_ ) );
NAND3_X1 _17324_ ( .A1(_04115_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_result_csreg_mem [9] ), .ZN(_01403_ ) );
OAI211_X1 _17325_ ( .A(_01378_ ), .B(_01403_ ), .C1(_02290_ ), .C2(_06295_ ), .ZN(_01404_ ) );
NOR2_X1 _17326_ ( .A1(_06279_ ), .A2(_01404_ ), .ZN(_01405_ ) );
NOR2_X1 _17327_ ( .A1(_01402_ ), .A2(_01405_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
AOI221_X4 _17328_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [8] ), .B2(_01391_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [8] ), .ZN(_01406_ ) );
AOI21_X1 _17329_ ( .A(\EX_LS_pc [8] ), .B1(_04102_ ), .B2(_01393_ ), .ZN(_01407_ ) );
NOR2_X1 _17330_ ( .A1(_01406_ ), .A2(_01407_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
OAI22_X1 _17331_ ( .A1(_06295_ ), .A2(_02292_ ), .B1(_04117_ ), .B2(_06382_ ), .ZN(_01408_ ) );
MUX2_X1 _17332_ ( .A(_01408_ ), .B(\EX_LS_pc [7] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _17333_ ( .A1(_06295_ ), .A2(_02293_ ), .B1(_04117_ ), .B2(_06383_ ), .ZN(_01409_ ) );
MUX2_X1 _17334_ ( .A(_01409_ ), .B(\EX_LS_pc [6] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
AOI21_X1 _17335_ ( .A(\EX_LS_pc [5] ), .B1(_04102_ ), .B2(_01378_ ), .ZN(_01410_ ) );
OAI21_X1 _17336_ ( .A(_01378_ ), .B1(_01391_ ), .B2(_06370_ ), .ZN(_01411_ ) );
AOI21_X1 _17337_ ( .A(_01411_ ), .B1(\LS_WB_wdata_csreg [5] ), .B2(_01391_ ), .ZN(_01412_ ) );
AOI21_X1 _17338_ ( .A(_01410_ ), .B1(_04103_ ), .B2(_01412_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
OAI22_X1 _17339_ ( .A1(_06295_ ), .A2(_02295_ ), .B1(_04117_ ), .B2(_06371_ ), .ZN(_01413_ ) );
MUX2_X1 _17340_ ( .A(_01413_ ), .B(\EX_LS_pc [4] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
OAI22_X1 _17341_ ( .A1(_06295_ ), .A2(_02296_ ), .B1(_04117_ ), .B2(_06372_ ), .ZN(_01414_ ) );
MUX2_X1 _17342_ ( .A(_01414_ ), .B(\EX_LS_pc [3] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
AOI221_X4 _17343_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [2] ), .B2(_01390_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [2] ), .ZN(_01415_ ) );
AOI21_X1 _17344_ ( .A(_01415_ ), .B1(_06270_ ), .B2(_01365_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
AOI21_X1 _17345_ ( .A(\EX_LS_pc [29] ), .B1(_01385_ ), .B2(_04111_ ), .ZN(_01416_ ) );
MUX2_X1 _17346_ ( .A(\LS_WB_wdata_csreg [29] ), .B(\EX_LS_result_csreg_mem [29] ), .S(_04105_ ), .Z(_01417_ ) );
NOR3_X1 _17347_ ( .A1(_06279_ ), .A2(_01362_ ), .A3(_01417_ ), .ZN(_01418_ ) );
NOR2_X1 _17348_ ( .A1(_01416_ ), .A2(_01418_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
AOI21_X1 _17349_ ( .A(\EX_LS_pc [1] ), .B1(_04102_ ), .B2(_01378_ ), .ZN(_01419_ ) );
OAI21_X1 _17350_ ( .A(_01378_ ), .B1(_01391_ ), .B2(_06374_ ), .ZN(_01420_ ) );
AOI21_X1 _17351_ ( .A(_01420_ ), .B1(\LS_WB_wdata_csreg [1] ), .B2(_01391_ ), .ZN(_01421_ ) );
AOI21_X1 _17352_ ( .A(_01419_ ), .B1(_04103_ ), .B2(_01421_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
OAI22_X1 _17353_ ( .A1(_06295_ ), .A2(_02300_ ), .B1(_04117_ ), .B2(_06375_ ), .ZN(_01422_ ) );
MUX2_X1 _17354_ ( .A(_01422_ ), .B(\EX_LS_pc [0] ), .S(_01365_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
AOI221_X4 _17355_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [28] ), .B2(_01390_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [28] ), .ZN(_01423_ ) );
AOI21_X1 _17356_ ( .A(\EX_LS_pc [28] ), .B1(_04102_ ), .B2(_01393_ ), .ZN(_01424_ ) );
NOR2_X1 _17357_ ( .A1(_01423_ ), .A2(_01424_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI221_X4 _17358_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [27] ), .B2(_01390_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [27] ), .ZN(_01425_ ) );
AOI21_X1 _17359_ ( .A(\EX_LS_pc [27] ), .B1(_04102_ ), .B2(_01393_ ), .ZN(_01426_ ) );
NOR2_X1 _17360_ ( .A1(_01425_ ), .A2(_01426_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI21_X1 _17361_ ( .A(\EX_LS_pc [26] ), .B1(_01385_ ), .B2(_01393_ ), .ZN(_01427_ ) );
MUX2_X1 _17362_ ( .A(\LS_WB_wdata_csreg [26] ), .B(\EX_LS_result_csreg_mem [26] ), .S(_04104_ ), .Z(_01428_ ) );
NOR3_X1 _17363_ ( .A1(_04101_ ), .A2(_01362_ ), .A3(_01428_ ), .ZN(_01429_ ) );
NOR2_X1 _17364_ ( .A1(_01427_ ), .A2(_01429_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI21_X1 _17365_ ( .A(\EX_LS_pc [25] ), .B1(_01385_ ), .B2(_01393_ ), .ZN(_01430_ ) );
MUX2_X1 _17366_ ( .A(\LS_WB_wdata_csreg [25] ), .B(\EX_LS_result_csreg_mem [25] ), .S(_04104_ ), .Z(_01431_ ) );
NOR3_X1 _17367_ ( .A1(_04101_ ), .A2(_01362_ ), .A3(_01431_ ), .ZN(_01432_ ) );
NOR2_X1 _17368_ ( .A1(_01430_ ), .A2(_01432_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI221_X4 _17369_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [24] ), .B2(_01390_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [24] ), .ZN(_01433_ ) );
AOI21_X1 _17370_ ( .A(\EX_LS_pc [24] ), .B1(_04102_ ), .B2(_01393_ ), .ZN(_01434_ ) );
NOR2_X1 _17371_ ( .A1(_01433_ ), .A2(_01434_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _17372_ ( .A(\EX_LS_pc [23] ), .B1(_04102_ ), .B2(_01378_ ), .ZN(_01435_ ) );
OAI21_X1 _17373_ ( .A(_01378_ ), .B1(_01391_ ), .B2(_06408_ ), .ZN(_01436_ ) );
AOI21_X1 _17374_ ( .A(_01436_ ), .B1(\LS_WB_wdata_csreg [23] ), .B2(_01391_ ), .ZN(_01437_ ) );
AOI21_X1 _17375_ ( .A(_01435_ ), .B1(_04103_ ), .B2(_01437_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
AOI221_X4 _17376_ ( .A(_01364_ ), .B1(\LS_WB_wdata_csreg [22] ), .B2(_01390_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [22] ), .ZN(_01438_ ) );
AOI21_X1 _17377_ ( .A(\EX_LS_pc [22] ), .B1(_04102_ ), .B2(_01378_ ), .ZN(_01439_ ) );
NOR2_X1 _17378_ ( .A1(_01438_ ), .A2(_01439_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
AOI21_X1 _17379_ ( .A(\EX_LS_pc [31] ), .B1(_01385_ ), .B2(_01393_ ), .ZN(_01440_ ) );
MUX2_X1 _17380_ ( .A(\LS_WB_wdata_csreg [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_04104_ ), .Z(_01441_ ) );
NOR3_X1 _17381_ ( .A1(_04101_ ), .A2(_01362_ ), .A3(_01441_ ), .ZN(_01442_ ) );
NOR2_X1 _17382_ ( .A1(_01440_ ), .A2(_01442_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17383_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01443_ ) );
INV_X1 _17384_ ( .A(_01443_ ), .ZN(_01444_ ) );
OR3_X1 _17385_ ( .A1(_00671_ ), .A2(_06259_ ), .A3(_01444_ ), .ZN(_01445_ ) );
NAND3_X1 _17386_ ( .A1(_00643_ ), .A2(_02220_ ), .A3(_01444_ ), .ZN(_01446_ ) );
NAND2_X1 _17387_ ( .A1(_01445_ ), .A2(_01446_ ), .ZN(_01447_ ) );
AND2_X1 _17388_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01448_ ) );
INV_X1 _17389_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01449_ ) );
AND2_X1 _17390_ ( .A1(_01448_ ), .A2(_01449_ ), .ZN(_01450_ ) );
BUF_X4 _17391_ ( .A(_01450_ ), .Z(_01451_ ) );
INV_X1 _17392_ ( .A(_01451_ ), .ZN(_01452_ ) );
NOR2_X1 _17393_ ( .A1(_01447_ ), .A2(_01452_ ), .ZN(_01453_ ) );
AND2_X1 _17394_ ( .A1(_01449_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01454_ ) );
INV_X1 _17395_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_01455_ ) );
AND2_X2 _17396_ ( .A1(_01454_ ), .A2(_01455_ ), .ZN(_01456_ ) );
NAND2_X1 _17397_ ( .A1(_01455_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01457_ ) );
NOR2_X1 _17398_ ( .A1(_01457_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01458_ ) );
OR2_X1 _17399_ ( .A1(_01456_ ), .A2(_01458_ ), .ZN(_01459_ ) );
NOR2_X4 _17400_ ( .A1(_01453_ ), .A2(_01459_ ), .ZN(_01460_ ) );
BUF_X4 _17401_ ( .A(_01460_ ), .Z(_01461_ ) );
NAND3_X1 _17402_ ( .A1(_00648_ ), .A2(_00653_ ), .A3(\io_master_arid [1] ), .ZN(_01462_ ) );
AND2_X2 _17403_ ( .A1(_01448_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01463_ ) );
NOR2_X1 _17404_ ( .A1(_01462_ ), .A2(_01463_ ), .ZN(_01464_ ) );
OAI21_X1 _17405_ ( .A(_01461_ ), .B1(_01464_ ), .B2(_01451_ ), .ZN(_01465_ ) );
INV_X1 _17406_ ( .A(_01456_ ), .ZN(_01466_ ) );
BUF_X4 _17407_ ( .A(_01466_ ), .Z(_01467_ ) );
BUF_X4 _17408_ ( .A(_01467_ ), .Z(_01468_ ) );
NOR2_X1 _17409_ ( .A1(_00671_ ), .A2(_06260_ ), .ZN(_01469_ ) );
NOR2_X1 _17410_ ( .A1(_06307_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01470_ ) );
NOR2_X2 _17411_ ( .A1(_00740_ ), .A2(_06259_ ), .ZN(_01471_ ) );
NOR2_X1 _17412_ ( .A1(_06303_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01472_ ) );
AOI22_X1 _17413_ ( .A1(_01469_ ), .A2(_01470_ ), .B1(_01471_ ), .B2(_01472_ ), .ZN(_01473_ ) );
AND3_X4 _17414_ ( .A1(_00699_ ), .A2(_00701_ ), .A3(_02220_ ), .ZN(_01474_ ) );
NAND2_X1 _17415_ ( .A1(_01474_ ), .A2(_01443_ ), .ZN(_01475_ ) );
NAND4_X1 _17416_ ( .A1(_00643_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_02220_ ), .ZN(_01476_ ) );
AND3_X1 _17417_ ( .A1(_01473_ ), .A2(_01475_ ), .A3(_01476_ ), .ZN(_01477_ ) );
BUF_X4 _17418_ ( .A(_01477_ ), .Z(_01478_ ) );
BUF_X4 _17419_ ( .A(_01478_ ), .Z(_01479_ ) );
OAI21_X1 _17420_ ( .A(_01465_ ), .B1(_01468_ ), .B2(_01479_ ), .ZN(_01480_ ) );
MUX2_X1 _17421_ ( .A(\EX_LS_result_reg [21] ), .B(_01480_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
BUF_X4 _17422_ ( .A(_01451_ ), .Z(_01481_ ) );
NAND3_X1 _17423_ ( .A1(_00654_ ), .A2(_00656_ ), .A3(\io_master_arid [1] ), .ZN(_01482_ ) );
NOR2_X1 _17424_ ( .A1(_01482_ ), .A2(_01463_ ), .ZN(_01483_ ) );
OAI21_X1 _17425_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01483_ ), .ZN(_01484_ ) );
OAI21_X1 _17426_ ( .A(_01484_ ), .B1(_01468_ ), .B2(_01479_ ), .ZN(_01485_ ) );
MUX2_X1 _17427_ ( .A(\EX_LS_result_reg [20] ), .B(_01485_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _17428_ ( .A1(_00657_ ), .A2(_00659_ ), .A3(\io_master_arid [1] ), .ZN(_01486_ ) );
NOR2_X1 _17429_ ( .A1(_01486_ ), .A2(_01463_ ), .ZN(_01487_ ) );
OAI21_X1 _17430_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01487_ ), .ZN(_01488_ ) );
OAI21_X1 _17431_ ( .A(_01488_ ), .B1(_01468_ ), .B2(_01479_ ), .ZN(_01489_ ) );
MUX2_X1 _17432_ ( .A(\EX_LS_result_reg [19] ), .B(_01489_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _17433_ ( .A1(_00660_ ), .A2(_00662_ ), .A3(\io_master_arid [1] ), .ZN(_01490_ ) );
NOR2_X1 _17434_ ( .A1(_01490_ ), .A2(_01463_ ), .ZN(_01491_ ) );
OAI21_X1 _17435_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01491_ ), .ZN(_01492_ ) );
OAI21_X1 _17436_ ( .A(_01492_ ), .B1(_01468_ ), .B2(_01479_ ), .ZN(_01493_ ) );
MUX2_X1 _17437_ ( .A(\EX_LS_result_reg [18] ), .B(_01493_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _17438_ ( .A1(_00663_ ), .A2(_00665_ ), .A3(\io_master_arid [1] ), .ZN(_01494_ ) );
NOR2_X1 _17439_ ( .A1(_01494_ ), .A2(_01463_ ), .ZN(_01495_ ) );
OAI21_X1 _17440_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01495_ ), .ZN(_01496_ ) );
OAI21_X1 _17441_ ( .A(_01496_ ), .B1(_01468_ ), .B2(_01478_ ), .ZN(_01497_ ) );
MUX2_X1 _17442_ ( .A(\EX_LS_result_reg [17] ), .B(_01497_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _17443_ ( .A1(_00666_ ), .A2(_00668_ ), .A3(_02220_ ), .ZN(_01498_ ) );
NOR2_X1 _17444_ ( .A1(_01498_ ), .A2(_01463_ ), .ZN(_01499_ ) );
OAI21_X1 _17445_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01499_ ), .ZN(_01500_ ) );
OAI21_X1 _17446_ ( .A(_01500_ ), .B1(_01468_ ), .B2(_01478_ ), .ZN(_01501_ ) );
MUX2_X1 _17447_ ( .A(\EX_LS_result_reg [16] ), .B(_01501_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
BUF_X4 _17448_ ( .A(_01448_ ), .Z(_01502_ ) );
NOR3_X1 _17449_ ( .A1(_01456_ ), .A2(_01502_ ), .A3(_01458_ ), .ZN(_01503_ ) );
NAND2_X1 _17450_ ( .A1(_01469_ ), .A2(_01503_ ), .ZN(_01504_ ) );
NAND2_X1 _17451_ ( .A1(_01447_ ), .A2(_01502_ ), .ZN(_01505_ ) );
OAI211_X1 _17452_ ( .A(_01504_ ), .B(_01505_ ), .C1(_01479_ ), .C2(_01467_ ), .ZN(_01506_ ) );
MUX2_X1 _17453_ ( .A(\EX_LS_result_reg [15] ), .B(_01506_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
INV_X1 _17454_ ( .A(_01502_ ), .ZN(_01507_ ) );
NOR2_X1 _17455_ ( .A1(_01507_ ), .A2(_01443_ ), .ZN(_01508_ ) );
OR2_X1 _17456_ ( .A1(_06260_ ), .A2(_01508_ ), .ZN(_01509_ ) );
NOR2_X1 _17457_ ( .A1(_01509_ ), .A2(_01459_ ), .ZN(_01510_ ) );
NAND3_X1 _17458_ ( .A1(_00673_ ), .A2(_00675_ ), .A3(_01510_ ), .ZN(_01511_ ) );
NOR2_X1 _17459_ ( .A1(_00646_ ), .A2(_06300_ ), .ZN(_01512_ ) );
NAND2_X1 _17460_ ( .A1(_01512_ ), .A2(_01508_ ), .ZN(_01513_ ) );
OAI211_X1 _17461_ ( .A(_01511_ ), .B(_01513_ ), .C1(_01479_ ), .C2(_01467_ ), .ZN(_01514_ ) );
MUX2_X1 _17462_ ( .A(\EX_LS_result_reg [14] ), .B(_01514_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
NOR2_X1 _17463_ ( .A1(_01028_ ), .A2(_06301_ ), .ZN(_01515_ ) );
NAND2_X1 _17464_ ( .A1(_01515_ ), .A2(_01508_ ), .ZN(_01516_ ) );
NAND3_X1 _17465_ ( .A1(_00676_ ), .A2(_00678_ ), .A3(_01510_ ), .ZN(_01517_ ) );
OAI211_X1 _17466_ ( .A(_01516_ ), .B(_01517_ ), .C1(_01479_ ), .C2(_01467_ ), .ZN(_01518_ ) );
MUX2_X1 _17467_ ( .A(\EX_LS_result_reg [13] ), .B(_01518_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _17468_ ( .A1(_00680_ ), .A2(_00683_ ), .A3(_01510_ ), .ZN(_01519_ ) );
NAND4_X1 _17469_ ( .A1(_00717_ ), .A2(_00719_ ), .A3(\io_master_arid [1] ), .A4(_01508_ ), .ZN(_01520_ ) );
OAI211_X1 _17470_ ( .A(_01519_ ), .B(_01520_ ), .C1(_01479_ ), .C2(_01467_ ), .ZN(_01521_ ) );
MUX2_X1 _17471_ ( .A(\EX_LS_result_reg [12] ), .B(_01521_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
NOR3_X1 _17472_ ( .A1(_00646_ ), .A2(_06300_ ), .A3(_01502_ ), .ZN(_01522_ ) );
OAI21_X2 _17473_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01522_ ), .ZN(_01523_ ) );
OAI21_X1 _17474_ ( .A(_01523_ ), .B1(_01468_ ), .B2(_01478_ ), .ZN(_01524_ ) );
MUX2_X1 _17475_ ( .A(\EX_LS_result_reg [30] ), .B(_01524_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NOR2_X1 _17476_ ( .A1(_01477_ ), .A2(_01466_ ), .ZN(_01525_ ) );
NOR2_X1 _17477_ ( .A1(_01525_ ), .A2(_06273_ ), .ZN(_01526_ ) );
AND3_X1 _17478_ ( .A1(_00687_ ), .A2(_00689_ ), .A3(_01510_ ), .ZN(_01527_ ) );
NOR2_X1 _17479_ ( .A1(_01221_ ), .A2(_06301_ ), .ZN(_01528_ ) );
AOI21_X1 _17480_ ( .A(_01527_ ), .B1(_01508_ ), .B2(_01528_ ), .ZN(_01529_ ) );
AOI22_X1 _17481_ ( .A1(_01526_ ), .A2(_01529_ ), .B1(_06273_ ), .B2(_04830_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
AND2_X1 _17482_ ( .A1(_00730_ ), .A2(_00731_ ), .ZN(_01530_ ) );
NOR2_X1 _17483_ ( .A1(_01530_ ), .A2(_06300_ ), .ZN(_01531_ ) );
NAND2_X1 _17484_ ( .A1(_01531_ ), .A2(_01508_ ), .ZN(_01532_ ) );
NAND3_X1 _17485_ ( .A1(_00690_ ), .A2(_00692_ ), .A3(_01510_ ), .ZN(_01533_ ) );
OAI211_X1 _17486_ ( .A(_01532_ ), .B(_01533_ ), .C1(_01479_ ), .C2(_01467_ ), .ZN(_01534_ ) );
MUX2_X1 _17487_ ( .A(\EX_LS_result_reg [10] ), .B(_01534_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17488_ ( .A1(_00693_ ), .A2(_00695_ ), .A3(_01510_ ), .ZN(_01535_ ) );
AND2_X1 _17489_ ( .A1(_00733_ ), .A2(_00734_ ), .ZN(_01536_ ) );
NOR2_X1 _17490_ ( .A1(_01536_ ), .A2(_06301_ ), .ZN(_01537_ ) );
AOI21_X1 _17491_ ( .A(_01535_ ), .B1(_01508_ ), .B2(_01537_ ), .ZN(_01538_ ) );
AOI22_X1 _17492_ ( .A1(_01526_ ), .A2(_01538_ ), .B1(_06273_ ), .B2(_04922_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _17493_ ( .A1(_00696_ ), .A2(_00698_ ), .A3(_01510_ ), .ZN(_01539_ ) );
NAND4_X1 _17494_ ( .A1(_00735_ ), .A2(_00737_ ), .A3(\io_master_arid [1] ), .A4(_01508_ ), .ZN(_01540_ ) );
OAI211_X1 _17495_ ( .A(_01539_ ), .B(_01540_ ), .C1(_01479_ ), .C2(_01467_ ), .ZN(_01541_ ) );
MUX2_X1 _17496_ ( .A(\EX_LS_result_reg [8] ), .B(_01541_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
MUX2_X2 _17497_ ( .A(_01471_ ), .B(_01474_ ), .S(_01443_ ), .Z(_01542_ ) );
MUX2_X2 _17498_ ( .A(_01474_ ), .B(_01542_ ), .S(_01463_ ), .Z(_01543_ ) );
MUX2_X2 _17499_ ( .A(_01542_ ), .B(_01543_ ), .S(_01452_ ), .Z(_01544_ ) );
OAI21_X2 _17500_ ( .A(_01544_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01457_ ), .ZN(_01545_ ) );
OR3_X1 _17501_ ( .A1(_01477_ ), .A2(\mylsu.typ_tmp [2] ), .A3(_01457_ ), .ZN(_01546_ ) );
AOI21_X1 _17502_ ( .A(_01456_ ), .B1(_01545_ ), .B2(_01546_ ), .ZN(_01547_ ) );
OR2_X2 _17503_ ( .A1(_01547_ ), .A2(_01525_ ), .ZN(_01548_ ) );
MUX2_X2 _17504_ ( .A(\EX_LS_result_reg [7] ), .B(_01548_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
NOR4_X1 _17505_ ( .A1(_00743_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(_06303_ ), .A4(_06260_ ), .ZN(_01549_ ) );
NOR3_X1 _17506_ ( .A1(_00646_ ), .A2(_06260_ ), .A3(_01472_ ), .ZN(_01550_ ) );
OAI22_X1 _17507_ ( .A1(_01549_ ), .A2(_01550_ ), .B1(_06307_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01551_ ) );
NAND4_X1 _17508_ ( .A1(_00673_ ), .A2(_00675_ ), .A3(_02220_ ), .A4(_01470_ ), .ZN(_01552_ ) );
AOI21_X1 _17509_ ( .A(_01443_ ), .B1(_01551_ ), .B2(_01552_ ), .ZN(_01553_ ) );
NOR3_X1 _17510_ ( .A1(_00704_ ), .A2(_06260_ ), .A3(_01444_ ), .ZN(_01554_ ) );
OAI21_X1 _17511_ ( .A(_01456_ ), .B1(_01553_ ), .B2(_01554_ ), .ZN(_01555_ ) );
OAI21_X1 _17512_ ( .A(_01458_ ), .B1(_01553_ ), .B2(_01554_ ), .ZN(_01556_ ) );
NOR3_X1 _17513_ ( .A1(_00743_ ), .A2(_06260_ ), .A3(_01443_ ), .ZN(_01557_ ) );
OAI21_X1 _17514_ ( .A(_01463_ ), .B1(_01557_ ), .B2(_01554_ ), .ZN(_01558_ ) );
OR3_X1 _17515_ ( .A1(_00704_ ), .A2(_06260_ ), .A3(_01463_ ), .ZN(_01559_ ) );
AOI21_X1 _17516_ ( .A(_01451_ ), .B1(_01558_ ), .B2(_01559_ ), .ZN(_01560_ ) );
INV_X1 _17517_ ( .A(_01557_ ), .ZN(_01561_ ) );
INV_X1 _17518_ ( .A(_01554_ ), .ZN(_01562_ ) );
AOI21_X1 _17519_ ( .A(_01452_ ), .B1(_01561_ ), .B2(_01562_ ), .ZN(_01563_ ) );
OAI22_X1 _17520_ ( .A1(_01560_ ), .A2(_01563_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01457_ ), .ZN(_01564_ ) );
AND2_X1 _17521_ ( .A1(_01556_ ), .A2(_01564_ ), .ZN(_01565_ ) );
OAI21_X1 _17522_ ( .A(_01555_ ), .B1(_01565_ ), .B2(_01456_ ), .ZN(_01566_ ) );
MUX2_X1 _17523_ ( .A(\EX_LS_result_reg [6] ), .B(_01566_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NOR2_X1 _17524_ ( .A1(_01503_ ), .A2(_01443_ ), .ZN(_01567_ ) );
INV_X1 _17525_ ( .A(_01567_ ), .ZN(_01568_ ) );
AND2_X2 _17526_ ( .A1(_01459_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01569_ ) );
NOR2_X1 _17527_ ( .A1(_01568_ ), .A2(_01569_ ), .ZN(_01570_ ) );
AOI211_X1 _17528_ ( .A(_06272_ ), .B(_06300_ ), .C1(_00858_ ), .C2(_01570_ ), .ZN(_01571_ ) );
NAND2_X1 _17529_ ( .A1(_00707_ ), .A2(_01568_ ), .ZN(_01572_ ) );
NAND2_X1 _17530_ ( .A1(_01571_ ), .A2(_01572_ ), .ZN(_01573_ ) );
MUX2_X1 _17531_ ( .A(_01028_ ), .B(_00993_ ), .S(_06303_ ), .Z(_01574_ ) );
AOI21_X1 _17532_ ( .A(_01573_ ), .B1(_01569_ ), .B2(_01574_ ), .ZN(_01575_ ) );
AND2_X1 _17533_ ( .A1(_06272_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01576_ ) );
OR2_X1 _17534_ ( .A1(_01575_ ), .A2(_01576_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
AOI221_X4 _17535_ ( .A(_06272_ ), .B1(_00880_ ), .B2(_01570_ ), .C1(_00710_ ), .C2(_01568_ ), .ZN(_01577_ ) );
AND3_X1 _17536_ ( .A1(_00717_ ), .A2(_00719_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01578_ ) );
OAI21_X1 _17537_ ( .A(_01569_ ), .B1(_01011_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01579_ ) );
OAI211_X1 _17538_ ( .A(_01577_ ), .B(\io_master_arid [1] ), .C1(_01578_ ), .C2(_01579_ ), .ZN(_01580_ ) );
NAND2_X1 _17539_ ( .A1(_06273_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_01581_ ) );
NAND2_X1 _17540_ ( .A1(_01580_ ), .A2(_01581_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _17541_ ( .A1(_06273_ ), .A2(\EX_LS_result_reg [3] ), .ZN(_01582_ ) );
AOI211_X1 _17542_ ( .A(_06272_ ), .B(_06301_ ), .C1(_00898_ ), .C2(_01570_ ), .ZN(_01583_ ) );
NAND2_X1 _17543_ ( .A1(_00713_ ), .A2(_01568_ ), .ZN(_01584_ ) );
NAND2_X1 _17544_ ( .A1(_01583_ ), .A2(_01584_ ), .ZN(_01585_ ) );
NAND3_X1 _17545_ ( .A1(_00687_ ), .A2(_06303_ ), .A3(_00689_ ), .ZN(_01586_ ) );
NAND4_X1 _17546_ ( .A1(_02170_ ), .A2(_02184_ ), .A3(_02224_ ), .A4(_00726_ ), .ZN(_01587_ ) );
OAI211_X1 _17547_ ( .A(\mylsu.araddr_tmp [1] ), .B(_01587_ ), .C1(_02229_ ), .C2(\io_master_rdata [27] ), .ZN(_01588_ ) );
AND3_X1 _17548_ ( .A1(_01586_ ), .A2(_01569_ ), .A3(_01588_ ), .ZN(_01589_ ) );
OAI21_X1 _17549_ ( .A(_01582_ ), .B1(_01585_ ), .B2(_01589_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
AOI211_X1 _17550_ ( .A(_06272_ ), .B(_06300_ ), .C1(_00913_ ), .C2(_01570_ ), .ZN(_01590_ ) );
NAND2_X1 _17551_ ( .A1(_00716_ ), .A2(_01568_ ), .ZN(_01591_ ) );
NAND2_X1 _17552_ ( .A1(_01590_ ), .A2(_01591_ ), .ZN(_01592_ ) );
MUX2_X1 _17553_ ( .A(_01530_ ), .B(_01057_ ), .S(_06303_ ), .Z(_01593_ ) );
AOI21_X1 _17554_ ( .A(_01592_ ), .B1(_01569_ ), .B2(_01593_ ), .ZN(_01594_ ) );
AND2_X1 _17555_ ( .A1(_06272_ ), .A2(\EX_LS_result_reg [2] ), .ZN(_01595_ ) );
OR2_X1 _17556_ ( .A1(_01594_ ), .A2(_01595_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
AOI211_X1 _17557_ ( .A(_06300_ ), .B(_01502_ ), .C1(_00685_ ), .C2(_00686_ ), .ZN(_01596_ ) );
OAI21_X1 _17558_ ( .A(_01460_ ), .B1(_01481_ ), .B2(_01596_ ), .ZN(_01597_ ) );
OAI21_X1 _17559_ ( .A(_01597_ ), .B1(_01468_ ), .B2(_01478_ ), .ZN(_01598_ ) );
MUX2_X1 _17560_ ( .A(\EX_LS_result_reg [29] ), .B(_01598_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
AOI211_X1 _17561_ ( .A(_06271_ ), .B(_06300_ ), .C1(_00930_ ), .C2(_01570_ ), .ZN(_01599_ ) );
NAND2_X1 _17562_ ( .A1(_00722_ ), .A2(_01568_ ), .ZN(_01600_ ) );
NAND2_X1 _17563_ ( .A1(_01599_ ), .A2(_01600_ ), .ZN(_01601_ ) );
MUX2_X1 _17564_ ( .A(_01536_ ), .B(_01074_ ), .S(_06303_ ), .Z(_01602_ ) );
AOI21_X1 _17565_ ( .A(_01601_ ), .B1(_01569_ ), .B2(_01602_ ), .ZN(_01603_ ) );
AND2_X1 _17566_ ( .A1(_06272_ ), .A2(\EX_LS_result_reg [1] ), .ZN(_01604_ ) );
OR2_X1 _17567_ ( .A1(_01603_ ), .A2(_01604_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
AOI211_X1 _17568_ ( .A(_06272_ ), .B(_06301_ ), .C1(_00945_ ), .C2(_01570_ ), .ZN(_01605_ ) );
NAND2_X1 _17569_ ( .A1(_00725_ ), .A2(_01568_ ), .ZN(_01606_ ) );
NAND2_X1 _17570_ ( .A1(_01605_ ), .A2(_01606_ ), .ZN(_01607_ ) );
NAND3_X1 _17571_ ( .A1(_00735_ ), .A2(\mylsu.araddr_tmp [1] ), .A3(_00737_ ), .ZN(_01608_ ) );
NAND3_X1 _17572_ ( .A1(_00696_ ), .A2(_06303_ ), .A3(_00698_ ), .ZN(_01609_ ) );
AND3_X1 _17573_ ( .A1(_01608_ ), .A2(_01609_ ), .A3(_01569_ ), .ZN(_01610_ ) );
OAI22_X1 _17574_ ( .A1(_01607_ ), .A2(_01610_ ), .B1(\mylsu.state [3] ), .B2(_04954_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
AND4_X1 _17575_ ( .A1(_02220_ ), .A2(_00717_ ), .A3(_00719_ ), .A4(_01507_ ), .ZN(_01611_ ) );
OAI21_X1 _17576_ ( .A(_01460_ ), .B1(_01451_ ), .B2(_01611_ ), .ZN(_01612_ ) );
OAI21_X1 _17577_ ( .A(_01612_ ), .B1(_01468_ ), .B2(_01478_ ), .ZN(_01613_ ) );
MUX2_X1 _17578_ ( .A(\EX_LS_result_reg [28] ), .B(_01613_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
AOI211_X1 _17579_ ( .A(_06301_ ), .B(_01502_ ), .C1(_00727_ ), .C2(_00728_ ), .ZN(_01614_ ) );
OAI21_X1 _17580_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01614_ ), .ZN(_01615_ ) );
AOI22_X1 _17581_ ( .A1(_01526_ ), .A2(_01615_ ), .B1(_06273_ ), .B2(_04702_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
AOI211_X1 _17582_ ( .A(_06300_ ), .B(_01502_ ), .C1(_00730_ ), .C2(_00731_ ), .ZN(_01616_ ) );
OAI21_X1 _17583_ ( .A(_01460_ ), .B1(_01451_ ), .B2(_01616_ ), .ZN(_01617_ ) );
OAI21_X1 _17584_ ( .A(_01617_ ), .B1(_01468_ ), .B2(_01478_ ), .ZN(_01618_ ) );
MUX2_X1 _17585_ ( .A(\EX_LS_result_reg [26] ), .B(_01618_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
AOI211_X1 _17586_ ( .A(_06301_ ), .B(_01502_ ), .C1(_00733_ ), .C2(_00734_ ), .ZN(_01619_ ) );
OAI21_X1 _17587_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01619_ ), .ZN(_01620_ ) );
AOI22_X1 _17588_ ( .A1(_01526_ ), .A2(_01620_ ), .B1(_06273_ ), .B2(_04655_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
AND4_X1 _17589_ ( .A1(_02220_ ), .A2(_00735_ ), .A3(_00737_ ), .A4(_01507_ ), .ZN(_01621_ ) );
OAI21_X1 _17590_ ( .A(_01460_ ), .B1(_01451_ ), .B2(_01621_ ), .ZN(_01622_ ) );
OAI21_X1 _17591_ ( .A(_01622_ ), .B1(_01467_ ), .B2(_01478_ ), .ZN(_01623_ ) );
MUX2_X1 _17592_ ( .A(\EX_LS_result_reg [24] ), .B(_01623_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _17593_ ( .A1(_00740_ ), .A2(_06301_ ), .A3(_01502_ ), .ZN(_01624_ ) );
OAI21_X1 _17594_ ( .A(_01461_ ), .B1(_01481_ ), .B2(_01624_ ), .ZN(_01625_ ) );
AOI22_X1 _17595_ ( .A1(_01526_ ), .A2(_01625_ ), .B1(_06273_ ), .B2(_04457_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _17596_ ( .A1(_00743_ ), .A2(_06300_ ), .A3(_01502_ ), .ZN(_01626_ ) );
OAI21_X1 _17597_ ( .A(_01460_ ), .B1(_01451_ ), .B2(_01626_ ), .ZN(_01627_ ) );
OAI21_X1 _17598_ ( .A(_01627_ ), .B1(_01467_ ), .B2(_01478_ ), .ZN(_01628_ ) );
MUX2_X1 _17599_ ( .A(\EX_LS_result_reg [22] ), .B(_01628_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17600_ ( .A1(_00643_ ), .A2(\io_master_arid [1] ), .A3(_01507_ ), .ZN(_01629_ ) );
OAI21_X1 _17601_ ( .A(_01460_ ), .B1(_01451_ ), .B2(_01629_ ), .ZN(_01630_ ) );
OAI21_X1 _17602_ ( .A(_01630_ ), .B1(_01467_ ), .B2(_01478_ ), .ZN(_01631_ ) );
MUX2_X1 _17603_ ( .A(\EX_LS_result_reg [31] ), .B(_01631_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17604_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(\LS_WB_waddr_reg [2] ), .ZN(_01632_ ) );
INV_X1 _17605_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01633_ ) );
INV_X1 _17606_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01634_ ) );
NAND3_X1 _17607_ ( .A1(_01632_ ), .A2(_01633_ ), .A3(_01634_ ), .ZN(_01635_ ) );
AND2_X1 _17608_ ( .A1(_01664_ ), .A2(LS_WB_wen_reg ), .ZN(_01636_ ) );
NAND2_X1 _17609_ ( .A1(_01635_ ), .A2(_01636_ ), .ZN(_01637_ ) );
BUF_X4 _17610_ ( .A(_01637_ ), .Z(_01638_ ) );
INV_X1 _17611_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01639_ ) );
INV_X1 _17612_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01640_ ) );
AOI21_X1 _17613_ ( .A(_01638_ ), .B1(_01639_ ), .B2(_01640_ ), .ZN(_01641_ ) );
NOR4_X1 _17614_ ( .A1(_01641_ ), .A2(_01633_ ), .A3(_01634_ ), .A4(_01638_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
AOI21_X1 _17615_ ( .A(_01638_ ), .B1(_01633_ ), .B2(_01634_ ), .ZN(_01642_ ) );
NOR2_X1 _17616_ ( .A1(_01637_ ), .A2(_01639_ ), .ZN(_01643_ ) );
NOR4_X1 _17617_ ( .A1(_01642_ ), .A2(_01643_ ), .A3(_01640_ ), .A4(_01638_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
NOR2_X1 _17618_ ( .A1(_01637_ ), .A2(_01633_ ), .ZN(_01644_ ) );
AND4_X1 _17619_ ( .A1(_01640_ ), .A2(_01644_ ), .A3(_01643_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR2_X1 _17620_ ( .A1(_01638_ ), .A2(_01640_ ), .ZN(_01645_ ) );
NOR4_X1 _17621_ ( .A1(_01642_ ), .A2(_01645_ ), .A3(_01639_ ), .A4(_01638_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
NOR2_X1 _17622_ ( .A1(_01638_ ), .A2(_01634_ ), .ZN(_01646_ ) );
AND4_X1 _17623_ ( .A1(_01640_ ), .A2(_01646_ ), .A3(_01643_ ), .A4(_01633_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
CLKBUF_X1 _17624_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17625_ ( .A1(_01641_ ), .A2(_01644_ ), .A3(_01634_ ), .A4(_01638_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17626_ ( .A1(_01639_ ), .A2(_01646_ ), .A3(_01645_ ), .A4(_01633_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17627_ ( .A1(_01639_ ), .A2(_01644_ ), .A3(_01645_ ), .A4(_01634_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
AND4_X1 _17628_ ( .A1(_01639_ ), .A2(_01644_ ), .A3(_01645_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
NOR4_X1 _17629_ ( .A1(_01642_ ), .A2(_01639_ ), .A3(_01640_ ), .A4(_01638_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17630_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01646_ ), .A3(_01643_ ), .A4(_01633_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17631_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01644_ ), .A3(_01643_ ), .A4(_01634_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17632_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01646_ ), .A3(_01643_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17633_ ( .A1(_01640_ ), .A2(_01644_ ), .A3(_01643_ ), .A4(_01634_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17634_ ( .A1(_01641_ ), .A2(_01646_ ), .A3(_01633_ ), .A4(_01638_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17635_ ( .A1(_02142_ ), .A2(_01813_ ), .A3(_02150_ ), .ZN(_01647_ ) );
NAND2_X1 _17636_ ( .A1(_01647_ ), .A2(_03903_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17637_ ( .A(reset ), .B(_02142_ ), .C1(_02143_ ), .C2(_02202_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17638_ ( .A(_01635_ ), .Z(_01648_ ) );
CLKBUF_X2 _17639_ ( .A(_01636_ ), .Z(_01649_ ) );
AND3_X1 _17640_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17641_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17642_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17643_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17644_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17645_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17646_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17647_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17648_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17649_ ( .A1(_01648_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01649_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17650_ ( .A(_01635_ ), .Z(_01650_ ) );
CLKBUF_X2 _17651_ ( .A(_01636_ ), .Z(_01651_ ) );
AND3_X1 _17652_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17653_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17654_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17655_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17656_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17657_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17658_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17659_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17660_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17661_ ( .A1(_01650_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01651_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17662_ ( .A(_01635_ ), .Z(_01652_ ) );
CLKBUF_X2 _17663_ ( .A(_01636_ ), .Z(_01653_ ) );
AND3_X1 _17664_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17665_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17666_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17667_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17668_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17669_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17670_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17671_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17672_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17673_ ( .A1(_01652_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01653_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17674_ ( .A1(_01635_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01636_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17675_ ( .A1(_01635_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01636_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_D ) );
AND3_X1 _17676_ ( .A1(_01813_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17677_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01654_ ) );
AND2_X1 _17678_ ( .A1(_01654_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01655_ ) );
INV_X1 _17679_ ( .A(_01655_ ), .ZN(_01656_ ) );
NOR2_X1 _17680_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01657_ ) );
OAI211_X1 _17681_ ( .A(_01664_ ), .B(\mysc.state [0] ), .C1(_01656_ ), .C2(_01657_ ), .ZN(_01658_ ) );
INV_X1 _17682_ ( .A(_01658_ ), .ZN(_01659_ ) );
OR3_X1 _17683_ ( .A1(_01659_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17684_ ( .A1(_01656_ ), .A2(reset ), .A3(_01657_ ), .ZN(_01660_ ) );
NAND2_X1 _17685_ ( .A1(_01660_ ), .A2(\mysc.state [0] ), .ZN(_01661_ ) );
OR3_X1 _17686_ ( .A1(_04141_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01662_ ) );
NAND2_X1 _17687_ ( .A1(_01661_ ), .A2(_01662_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17688_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_08077_ ) );
CLKGATE_X1 _17689_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_08078_ ) );
CLKGATE_X1 _17690_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_08079_ ) );
CLKGATE_X1 _17691_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08080_ ) );
CLKGATE_X1 _17692_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08081_ ) );
CLKGATE_X1 _17693_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08082_ ) );
CLKGATE_X1 _17694_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08083_ ) );
CLKGATE_X1 _17695_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_08084_ ) );
CLKGATE_X1 _17696_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_08085_ ) );
CLKGATE_X1 _17697_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_08086_ ) );
CLKGATE_X1 _17698_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_08087_ ) );
CLKGATE_X1 _17699_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08088_ ) );
CLKGATE_X1 _17700_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08089_ ) );
CLKGATE_X1 _17701_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08090_ ) );
CLKGATE_X1 _17702_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_08091_ ) );
CLKGATE_X1 _17703_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_08092_ ) );
CLKGATE_X1 _17704_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_08093_ ) );
CLKGATE_X1 _17705_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08094_ ) );
CLKGATE_X1 _17706_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_08095_ ) );
CLKGATE_X1 _17707_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ), .GCK(_08096_ ) );
CLKGATE_X1 _17708_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .GCK(_08097_ ) );
CLKGATE_X1 _17709_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08098_ ) );
CLKGATE_X1 _17710_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_08099_ ) );
CLKGATE_X1 _17711_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_08100_ ) );
CLKGATE_X1 _17712_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_08101_ ) );
CLKGATE_X1 _17713_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_08102_ ) );
CLKGATE_X1 _17714_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_08103_ ) );
CLKGATE_X1 _17715_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_08104_ ) );
CLKGATE_X1 _17716_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_08105_ ) );
CLKGATE_X1 _17717_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_08106_ ) );
CLKGATE_X1 _17718_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_08107_ ) );
CLKGATE_X1 _17719_ ( .CK(clock ), .E(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ), .GCK(_08108_ ) );
CLKGATE_X1 _17720_ ( .CK(clock ), .E(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ), .GCK(_08109_ ) );
CLKGATE_X1 _17721_ ( .CK(clock ), .E(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ), .GCK(_08110_ ) );
CLKGATE_X1 _17722_ ( .CK(clock ), .E(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ), .GCK(_08111_ ) );
CLKGATE_X1 _17723_ ( .CK(clock ), .E(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ), .GCK(_08112_ ) );
CLKGATE_X1 _17724_ ( .CK(clock ), .E(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ), .GCK(_08113_ ) );
CLKGATE_X1 _17725_ ( .CK(clock ), .E(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ), .GCK(_08114_ ) );
CLKGATE_X1 _17726_ ( .CK(clock ), .E(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ), .GCK(_08115_ ) );
CLKGATE_X1 _17727_ ( .CK(clock ), .E(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ), .GCK(_08116_ ) );
CLKGATE_X1 _17728_ ( .CK(clock ), .E(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ), .GCK(_08117_ ) );
CLKGATE_X1 _17729_ ( .CK(clock ), .E(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ), .GCK(_08118_ ) );
CLKGATE_X1 _17730_ ( .CK(clock ), .E(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ), .GCK(_08119_ ) );
CLKGATE_X1 _17731_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08120_ ) );
CLKGATE_X1 _17732_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08121_ ) );
CLKGATE_X1 _17733_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_08122_ ) );
CLKGATE_X1 _17734_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08123_ ) );
CLKGATE_X1 _17735_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08124_ ) );
CLKGATE_X1 _17736_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08125_ ) );
CLKGATE_X1 _17737_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08126_ ) );
CLKGATE_X1 _17738_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08127_ ) );
CLKGATE_X1 _17739_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_08128_ ) );
CLKGATE_X1 _17740_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08129_ ) );
CLKGATE_X1 _17741_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08130_ ) );
CLKGATE_X1 _17742_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08131_ ) );
CLKGATE_X1 _17743_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08132_ ) );
CLKGATE_X1 _17744_ ( .CK(clock ), .E(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08133_ ) );
CLKGATE_X1 _17745_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_08134_ ) );
CLKGATE_X1 _17746_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ), .GCK(_08135_ ) );
CLKGATE_X1 _17747_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08136_ ) );
CLKGATE_X1 _17748_ ( .CK(clock ), .E(\myec.state_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08137_ ) );
CLKGATE_X1 _17749_ ( .CK(clock ), .E(\mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ), .GCK(_08138_ ) );
CLKGATE_X1 _17750_ ( .CK(clock ), .E(\mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ), .GCK(_08139_ ) );
CLKGATE_X1 _17751_ ( .CK(clock ), .E(\mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ), .GCK(_08140_ ) );
CLKGATE_X1 _17752_ ( .CK(clock ), .E(\mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ), .GCK(_08141_ ) );
LOGIC1_X1 _17753_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17754_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00064_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00065_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08470_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08469_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08468_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08467_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08466_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08465_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08464_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08463_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08462_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08461_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08460_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08459_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08458_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08457_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08456_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08455_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08454_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08453_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08452_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08451_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08450_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08449_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08448_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08447_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08446_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08445_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08444_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08443_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08442_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08441_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08440_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08141_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08439_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08140_ ), .Q(\mtvec [31] ), .QN(_08438_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08140_ ), .Q(\mtvec [30] ), .QN(_08437_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08140_ ), .Q(\mtvec [21] ), .QN(_08436_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08140_ ), .Q(\mtvec [20] ), .QN(_08435_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08140_ ), .Q(\mtvec [19] ), .QN(_08434_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08140_ ), .Q(\mtvec [18] ), .QN(_08433_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08140_ ), .Q(\mtvec [17] ), .QN(_08432_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08140_ ), .Q(\mtvec [16] ), .QN(_08431_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08140_ ), .Q(\mtvec [15] ), .QN(_08430_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08140_ ), .Q(\mtvec [14] ), .QN(_08429_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08140_ ), .Q(\mtvec [13] ), .QN(_08428_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08140_ ), .Q(\mtvec [12] ), .QN(_08427_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08140_ ), .Q(\mtvec [29] ), .QN(_08426_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08140_ ), .Q(\mtvec [11] ), .QN(_08425_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08140_ ), .Q(\mtvec [10] ), .QN(_08424_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08140_ ), .Q(\mtvec [9] ), .QN(_08423_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08140_ ), .Q(\mtvec [8] ), .QN(_08422_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08140_ ), .Q(\mtvec [7] ), .QN(_08421_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08140_ ), .Q(\mtvec [6] ), .QN(_08420_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08140_ ), .Q(\mtvec [5] ), .QN(_08419_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08140_ ), .Q(\mtvec [4] ), .QN(_08418_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08140_ ), .Q(\mtvec [3] ), .QN(_08417_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08140_ ), .Q(\mtvec [2] ), .QN(_08416_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08140_ ), .Q(\mtvec [28] ), .QN(_08415_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08140_ ), .Q(\mtvec [1] ), .QN(_08414_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08140_ ), .Q(\mtvec [0] ), .QN(_08413_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08140_ ), .Q(\mtvec [27] ), .QN(_08412_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08140_ ), .Q(\mtvec [26] ), .QN(_08411_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08140_ ), .Q(\mtvec [25] ), .QN(_08410_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08140_ ), .Q(\mtvec [24] ), .QN(_08409_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08140_ ), .Q(\mtvec [23] ), .QN(_08408_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08140_ ), .Q(\mtvec [22] ), .QN(_08407_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08139_ ), .Q(\mepc [31] ), .QN(_08406_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08139_ ), .Q(\mepc [30] ), .QN(_08405_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08139_ ), .Q(\mepc [21] ), .QN(_08404_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08139_ ), .Q(\mepc [20] ), .QN(_08403_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08139_ ), .Q(\mepc [19] ), .QN(_08402_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08139_ ), .Q(\mepc [18] ), .QN(_08401_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08139_ ), .Q(\mepc [17] ), .QN(_08400_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08139_ ), .Q(\mepc [16] ), .QN(_08399_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08139_ ), .Q(\mepc [15] ), .QN(_08398_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08139_ ), .Q(\mepc [14] ), .QN(_08397_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08139_ ), .Q(\mepc [13] ), .QN(_08396_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08139_ ), .Q(\mepc [12] ), .QN(_08395_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08139_ ), .Q(\mepc [29] ), .QN(_08394_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08139_ ), .Q(\mepc [11] ), .QN(_08393_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08139_ ), .Q(\mepc [10] ), .QN(_08392_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08139_ ), .Q(\mepc [9] ), .QN(_08391_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08139_ ), .Q(\mepc [8] ), .QN(_08390_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08139_ ), .Q(\mepc [7] ), .QN(_08389_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08139_ ), .Q(\mepc [6] ), .QN(_08388_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08139_ ), .Q(\mepc [5] ), .QN(_08387_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08139_ ), .Q(\mepc [4] ), .QN(_08386_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08139_ ), .Q(\mepc [3] ), .QN(_08385_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08139_ ), .Q(\mepc [2] ), .QN(_08384_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08139_ ), .Q(\mepc [28] ), .QN(_08383_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08139_ ), .Q(\mepc [1] ), .QN(_08382_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08139_ ), .Q(\mepc [0] ), .QN(_08381_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08139_ ), .Q(\mepc [27] ), .QN(_08380_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08139_ ), .Q(\mepc [26] ), .QN(_08379_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08139_ ), .Q(\mepc [25] ), .QN(_08378_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08139_ ), .Q(\mepc [24] ), .QN(_08377_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08139_ ), .Q(\mepc [23] ), .QN(_08376_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08139_ ), .Q(\mepc [22] ), .QN(_08375_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q ( .D(_00097_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08374_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_1 ( .D(_00098_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08373_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_10 ( .D(_00099_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08372_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_11 ( .D(_00100_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08371_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_12 ( .D(_00101_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08370_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_13 ( .D(_00102_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08369_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_14 ( .D(_00103_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08368_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_15 ( .D(_00104_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08367_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_16 ( .D(_00105_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08366_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_17 ( .D(_00106_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08365_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_18 ( .D(_00107_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08364_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_19 ( .D(_00108_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08363_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_2 ( .D(_00109_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08362_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_20 ( .D(_00110_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08361_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_21 ( .D(_00111_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08360_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_22 ( .D(_00112_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08359_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_23 ( .D(_00113_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08358_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_24 ( .D(_00114_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08357_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_25 ( .D(_00115_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08356_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_26 ( .D(_00116_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08355_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_27 ( .D(_00117_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08354_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_28 ( .D(_00118_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08353_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_29 ( .D(_00119_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08352_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_3 ( .D(_00120_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08351_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_30 ( .D(_00121_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08350_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_31 ( .D(_00122_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08349_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_4 ( .D(_00123_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08348_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_5 ( .D(_00124_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08347_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_6 ( .D(_00125_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08346_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_7 ( .D(_00126_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08345_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_8 ( .D(_00127_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08344_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_9 ( .D(_00128_ ), .CK(_08138_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08471_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PP0__Q ( .D(_00129_ ), .CK(clock ), .Q(excp_written ), .QN(_08472_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08343_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08473_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08474_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08475_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08476_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08477_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08478_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08479_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08480_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08481_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08482_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08483_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08484_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08485_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08486_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08487_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08488_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08489_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08490_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08491_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08492_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08493_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08494_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08495_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08496_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08497_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08498_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08499_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08500_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08501_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08502_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08137_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08342_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00130_ ), .CK(_08136_ ), .Q(\myec.state [1] ), .QN(_08341_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00131_ ), .CK(_08136_ ), .Q(\myec.state [0] ), .QN(_08503_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PN0__Q ( .D(_00132_ ), .CK(clock ), .Q(check_quest ), .QN(_08504_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08340_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08505_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08506_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08507_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08508_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08509_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08510_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08511_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08512_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08513_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08514_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08339_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00133_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08338_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00134_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08337_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00135_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08336_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00136_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08335_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00137_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08334_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00138_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08333_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00139_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08332_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00140_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08331_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00141_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08330_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00142_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08329_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00143_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08328_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00144_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08327_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00145_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08326_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00146_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08325_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00147_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08324_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00148_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08323_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00149_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08322_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00150_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08321_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00151_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08320_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00152_ ), .CK(_08135_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08319_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q ( .D(_00153_ ), .CK(_08134_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08318_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_1 ( .D(_00154_ ), .CK(_08134_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08317_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_2 ( .D(_00155_ ), .CK(_08134_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08316_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_3 ( .D(_00156_ ), .CK(_08134_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08315_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_4 ( .D(_00157_ ), .CK(_08134_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08314_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q ( .D(_00158_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [30] ), .QN(_08313_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_1 ( .D(_00159_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [29] ), .QN(_08312_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_10 ( .D(_00160_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [20] ), .QN(_08311_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_11 ( .D(_00161_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [19] ), .QN(_08310_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_12 ( .D(_00162_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [18] ), .QN(_08309_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_13 ( .D(_00163_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [17] ), .QN(_08308_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_14 ( .D(_00164_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [16] ), .QN(_08307_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_15 ( .D(_00165_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [15] ), .QN(_08306_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_16 ( .D(_00166_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [14] ), .QN(_08305_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_17 ( .D(_00167_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [13] ), .QN(_08304_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_18 ( .D(_00168_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [12] ), .QN(_08303_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_19 ( .D(_00169_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [11] ), .QN(_08302_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_2 ( .D(_00170_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [28] ), .QN(_08301_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_20 ( .D(_00171_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [10] ), .QN(_08300_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_21 ( .D(_00172_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [9] ), .QN(_08299_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_22 ( .D(_00173_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [8] ), .QN(_08298_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_23 ( .D(_00174_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [7] ), .QN(_08297_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_24 ( .D(_00175_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [6] ), .QN(_08296_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_25 ( .D(_00176_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [5] ), .QN(_08295_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_26 ( .D(_00177_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [4] ), .QN(_08294_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_27 ( .D(_00178_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [3] ), .QN(_08293_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_28 ( .D(_00179_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [2] ), .QN(_08292_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_29 ( .D(_00180_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [1] ), .QN(_08291_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_3 ( .D(_00181_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [27] ), .QN(_08290_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_30 ( .D(_00182_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [0] ), .QN(_08289_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_4 ( .D(_00183_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [26] ), .QN(_08288_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_5 ( .D(_00184_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [25] ), .QN(_08287_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_6 ( .D(_00185_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [24] ), .QN(_08286_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_7 ( .D(_00186_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [23] ), .QN(_08285_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_8 ( .D(_00187_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [22] ), .QN(_08284_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_9 ( .D(_00188_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [21] ), .QN(_08283_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN1P__Q ( .D(_00189_ ), .CK(_08133_ ), .Q(\myexu.pc_jump [31] ), .QN(_08282_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q ( .D(_00190_ ), .CK(_08134_ ), .Q(\EX_LS_pc [31] ), .QN(_08281_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_1 ( .D(_00191_ ), .CK(_08134_ ), .Q(\EX_LS_pc [30] ), .QN(_08280_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_10 ( .D(_00192_ ), .CK(_08134_ ), .Q(\EX_LS_pc [21] ), .QN(_08279_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_11 ( .D(_00193_ ), .CK(_08134_ ), .Q(\EX_LS_pc [20] ), .QN(_08278_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_12 ( .D(_00194_ ), .CK(_08134_ ), .Q(\EX_LS_pc [19] ), .QN(_08277_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_13 ( .D(_00195_ ), .CK(_08134_ ), .Q(\EX_LS_pc [18] ), .QN(_08276_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_14 ( .D(_00196_ ), .CK(_08134_ ), .Q(\EX_LS_pc [17] ), .QN(_08275_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_15 ( .D(_00197_ ), .CK(_08134_ ), .Q(\EX_LS_pc [16] ), .QN(_08274_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_16 ( .D(_00198_ ), .CK(_08134_ ), .Q(\EX_LS_pc [15] ), .QN(_08273_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_17 ( .D(_00199_ ), .CK(_08134_ ), .Q(\EX_LS_pc [14] ), .QN(_08272_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_18 ( .D(_00200_ ), .CK(_08134_ ), .Q(\EX_LS_pc [13] ), .QN(_08271_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_19 ( .D(_00201_ ), .CK(_08134_ ), .Q(\EX_LS_pc [12] ), .QN(_08270_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_2 ( .D(_00202_ ), .CK(_08134_ ), .Q(\EX_LS_pc [29] ), .QN(_08269_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_20 ( .D(_00203_ ), .CK(_08134_ ), .Q(\EX_LS_pc [11] ), .QN(_08268_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_21 ( .D(_00204_ ), .CK(_08134_ ), .Q(\EX_LS_pc [10] ), .QN(_08267_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_22 ( .D(_00205_ ), .CK(_08134_ ), .Q(\EX_LS_pc [9] ), .QN(_08266_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_23 ( .D(_00206_ ), .CK(_08134_ ), .Q(\EX_LS_pc [8] ), .QN(_08265_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_24 ( .D(_00207_ ), .CK(_08134_ ), .Q(\EX_LS_pc [7] ), .QN(_08264_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_25 ( .D(_00208_ ), .CK(_08134_ ), .Q(\EX_LS_pc [6] ), .QN(_08263_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_26 ( .D(_00209_ ), .CK(_08134_ ), .Q(\EX_LS_pc [5] ), .QN(_08262_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_27 ( .D(_00210_ ), .CK(_08134_ ), .Q(\EX_LS_pc [4] ), .QN(_08261_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_28 ( .D(_00211_ ), .CK(_08134_ ), .Q(\EX_LS_pc [3] ), .QN(_08260_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_29 ( .D(_00212_ ), .CK(_08134_ ), .Q(\EX_LS_pc [2] ), .QN(_08259_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_3 ( .D(_00213_ ), .CK(_08134_ ), .Q(\EX_LS_pc [28] ), .QN(_08258_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_30 ( .D(_00214_ ), .CK(_08134_ ), .Q(\EX_LS_pc [1] ), .QN(_08257_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_31 ( .D(_00215_ ), .CK(_08134_ ), .Q(\EX_LS_pc [0] ), .QN(_08256_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_4 ( .D(_00216_ ), .CK(_08134_ ), .Q(\EX_LS_pc [27] ), .QN(_08255_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_5 ( .D(_00217_ ), .CK(_08134_ ), .Q(\EX_LS_pc [26] ), .QN(_08254_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_6 ( .D(_00218_ ), .CK(_08134_ ), .Q(\EX_LS_pc [25] ), .QN(_08253_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_7 ( .D(_00219_ ), .CK(_08134_ ), .Q(\EX_LS_pc [24] ), .QN(_08252_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_8 ( .D(_00220_ ), .CK(_08134_ ), .Q(\EX_LS_pc [23] ), .QN(_08251_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_9 ( .D(_00221_ ), .CK(_08134_ ), .Q(\EX_LS_pc [22] ), .QN(_08515_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08516_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08517_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08518_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08519_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08520_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08521_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08522_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08523_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08524_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08525_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08526_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08527_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08528_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08529_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08530_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08531_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08532_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08533_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08534_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08535_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08536_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08537_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08538_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08539_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08540_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08541_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08542_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08543_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08544_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08545_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08546_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08135_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08547_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08135_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PN0__Q ( .D(_00223_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q ( .D(_00222_ ), .CK(_08134_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_1 ( .D(_00224_ ), .CK(_08134_ ), .Q(\EX_LS_flag [1] ), .QN(_08250_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_2 ( .D(_00225_ ), .CK(_08134_ ), .Q(\EX_LS_flag [0] ), .QN(_08249_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_3 ( .D(_00226_ ), .CK(_08134_ ), .Q(\EX_LS_typ [4] ), .QN(_08248_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_4 ( .D(_00227_ ), .CK(_08134_ ), .Q(\EX_LS_typ [3] ), .QN(_08247_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_5 ( .D(_00228_ ), .CK(_08134_ ), .Q(\EX_LS_typ [2] ), .QN(_08246_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_6 ( .D(_00229_ ), .CK(_08134_ ), .Q(\EX_LS_typ [1] ), .QN(_08245_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_7 ( .D(_00230_ ), .CK(_08134_ ), .Q(\EX_LS_typ [0] ), .QN(_08244_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_08132_ ), .Q(\ID_EX_csr [11] ), .QN(_08243_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00232_ ), .CK(_08132_ ), .Q(\ID_EX_csr [10] ), .QN(_08242_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00233_ ), .CK(_08132_ ), .Q(\ID_EX_csr [1] ), .QN(_08241_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00234_ ), .CK(_08132_ ), .Q(\ID_EX_csr [0] ), .QN(_08240_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00235_ ), .CK(_08132_ ), .Q(\ID_EX_csr [9] ), .QN(_08239_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00236_ ), .CK(_08132_ ), .Q(\ID_EX_csr [8] ), .QN(_08238_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00237_ ), .CK(_08132_ ), .Q(\ID_EX_csr [7] ), .QN(_08237_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00238_ ), .CK(_08132_ ), .Q(\ID_EX_csr [6] ), .QN(_08236_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00239_ ), .CK(_08132_ ), .Q(\ID_EX_csr [5] ), .QN(_08235_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00240_ ), .CK(_08132_ ), .Q(\ID_EX_csr [4] ), .QN(_08234_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00241_ ), .CK(_08132_ ), .Q(\ID_EX_csr [3] ), .QN(_08233_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00242_ ), .CK(_08132_ ), .Q(\ID_EX_csr [2] ), .QN(_08232_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00243_ ), .CK(_08131_ ), .Q(exception_quest_IDU ), .QN(_08231_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00244_ ), .CK(_08130_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08129_ ), .Q(\ID_EX_imm [31] ), .QN(_08548_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08129_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08129_ ), .Q(\ID_EX_imm [21] ), .QN(_08549_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08129_ ), .Q(\ID_EX_imm [20] ), .QN(_08550_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08129_ ), .Q(\ID_EX_imm [19] ), .QN(_08551_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08129_ ), .Q(\ID_EX_imm [18] ), .QN(_08552_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08129_ ), .Q(\ID_EX_imm [17] ), .QN(_08553_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08129_ ), .Q(\ID_EX_imm [16] ), .QN(_08554_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08129_ ), .Q(\ID_EX_imm [15] ), .QN(_08555_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08129_ ), .Q(\ID_EX_imm [14] ), .QN(_08556_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08129_ ), .Q(\ID_EX_imm [13] ), .QN(_08557_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08129_ ), .Q(\ID_EX_imm [12] ), .QN(_08558_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08129_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08129_ ), .Q(\ID_EX_imm [11] ), .QN(_08559_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08129_ ), .Q(\ID_EX_imm [10] ), .QN(_08560_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08129_ ), .Q(\ID_EX_imm [9] ), .QN(_08561_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08129_ ), .Q(\ID_EX_imm [8] ), .QN(_08562_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08129_ ), .Q(\ID_EX_imm [7] ), .QN(_08563_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08129_ ), .Q(\ID_EX_imm [6] ), .QN(_08564_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08129_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08129_ ), .Q(\ID_EX_imm [4] ), .QN(_08565_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08129_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08129_ ), .Q(\ID_EX_imm [2] ), .QN(_08566_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08129_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08129_ ), .Q(\ID_EX_imm [1] ), .QN(_08567_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08129_ ), .Q(\ID_EX_imm [0] ), .QN(_08568_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08129_ ), .Q(\ID_EX_imm [27] ), .QN(_08569_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08129_ ), .Q(\ID_EX_imm [26] ), .QN(_08570_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08129_ ), .Q(\ID_EX_imm [25] ), .QN(_08571_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08129_ ), .Q(\ID_EX_imm [24] ), .QN(_08572_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08129_ ), .Q(\ID_EX_imm [23] ), .QN(_08573_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08129_ ), .Q(\ID_EX_imm [22] ), .QN(_08574_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08128_ ), .Q(\ID_EX_pc [31] ), .QN(_08575_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08128_ ), .Q(\ID_EX_pc [30] ), .QN(_08576_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08128_ ), .Q(\ID_EX_pc [21] ), .QN(_08577_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08128_ ), .Q(\ID_EX_pc [20] ), .QN(_08578_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08128_ ), .Q(\ID_EX_pc [19] ), .QN(_08579_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08128_ ), .Q(\ID_EX_pc [18] ), .QN(_08580_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08128_ ), .Q(\ID_EX_pc [17] ), .QN(_08581_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08128_ ), .Q(\ID_EX_pc [16] ), .QN(_08582_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08128_ ), .Q(\ID_EX_pc [15] ), .QN(_08583_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08128_ ), .Q(\ID_EX_pc [14] ), .QN(_08584_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08128_ ), .Q(\ID_EX_pc [13] ), .QN(_08585_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08128_ ), .Q(\ID_EX_pc [12] ), .QN(_08586_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08128_ ), .Q(\ID_EX_pc [29] ), .QN(_08587_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08128_ ), .Q(\ID_EX_pc [11] ), .QN(_08588_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08128_ ), .Q(\ID_EX_pc [10] ), .QN(_08589_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08128_ ), .Q(\ID_EX_pc [9] ), .QN(_08590_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08128_ ), .Q(\ID_EX_pc [8] ), .QN(_08591_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08128_ ), .Q(\ID_EX_pc [7] ), .QN(_08592_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08128_ ), .Q(\ID_EX_pc [6] ), .QN(_08593_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08128_ ), .Q(\ID_EX_pc [5] ), .QN(_08594_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08128_ ), .Q(\ID_EX_pc [4] ), .QN(_08595_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08128_ ), .Q(\ID_EX_pc [3] ), .QN(_08596_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08128_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08128_ ), .Q(\ID_EX_pc [28] ), .QN(_08597_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08128_ ), .Q(\ID_EX_pc [1] ), .QN(_08598_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08128_ ), .Q(\ID_EX_pc [0] ), .QN(_08599_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08128_ ), .Q(\ID_EX_pc [27] ), .QN(_08600_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08128_ ), .Q(\ID_EX_pc [26] ), .QN(_08601_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08128_ ), .Q(\ID_EX_pc [25] ), .QN(_08602_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08128_ ), .Q(\ID_EX_pc [24] ), .QN(_08603_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08128_ ), .Q(\ID_EX_pc [23] ), .QN(_08604_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08128_ ), .Q(\ID_EX_pc [22] ), .QN(_08230_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_08127_ ), .Q(\ID_EX_rd [4] ), .QN(_08229_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_08127_ ), .Q(\ID_EX_rd [3] ), .QN(_08228_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00247_ ), .CK(_08127_ ), .Q(\ID_EX_rd [2] ), .QN(_08227_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00248_ ), .CK(_08127_ ), .Q(\ID_EX_rd [1] ), .QN(_08226_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00249_ ), .CK(_08127_ ), .Q(\ID_EX_rd [0] ), .QN(_08225_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00250_ ), .CK(_08126_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08224_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00251_ ), .CK(_08126_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08223_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00253_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08221_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00252_ ), .CK(_08126_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08222_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00255_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08219_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00254_ ), .CK(_08126_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08220_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00257_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08217_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00256_ ), .CK(_08126_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08218_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00259_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08215_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00258_ ), .CK(_08125_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08216_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00260_ ), .CK(_08125_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08214_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00262_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08212_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00261_ ), .CK(_08125_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08213_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00264_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08210_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00263_ ), .CK(_08125_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08211_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00266_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08208_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00265_ ), .CK(_08125_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08209_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00268_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08206_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00267_ ), .CK(_08124_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08207_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00269_ ), .CK(_08123_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08205_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08606_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00270_ ), .CK(_08122_ ), .Q(\ID_EX_typ [7] ), .QN(_08605_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00271_ ), .CK(_08122_ ), .Q(\ID_EX_typ [6] ), .QN(_08204_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00272_ ), .CK(_08122_ ), .Q(\ID_EX_typ [5] ), .QN(_08203_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00273_ ), .CK(_08122_ ), .Q(\ID_EX_typ [4] ), .QN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00274_ ), .CK(_08122_ ), .Q(\ID_EX_typ [3] ), .QN(_08202_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00275_ ), .CK(_08122_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00276_ ), .CK(_08122_ ), .Q(\ID_EX_typ [1] ), .QN(_08201_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00277_ ), .CK(_08122_ ), .Q(\ID_EX_typ [0] ), .QN(_08607_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08121_ ), .Q(check_assert ), .QN(_08608_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08120_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08120_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08120_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08120_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08120_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08120_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08120_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08120_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08120_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08120_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08120_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08120_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08120_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08120_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08120_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08120_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08120_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08120_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08120_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08120_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08120_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08120_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08120_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08120_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08120_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08120_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08120_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08120_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08120_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08120_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08120_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08120_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08119_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08118_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08117_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08116_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08115_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08114_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08113_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08855_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08856_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08857_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08858_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08859_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08860_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08861_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08862_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08863_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08112_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08864_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08865_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08866_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08867_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08868_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08869_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08870_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08871_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08872_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08873_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08874_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08875_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08876_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08877_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08878_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08879_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08880_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08881_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08882_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08883_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08884_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08885_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08886_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08887_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08888_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08889_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08890_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08111_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08891_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08892_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08893_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08894_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08895_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08896_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08897_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08898_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08899_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08900_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08901_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08902_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08903_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08904_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08905_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08906_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08907_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08908_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08909_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08910_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08911_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08912_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08913_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08914_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08915_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08916_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08917_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08110_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08918_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08919_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08920_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08921_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08922_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08923_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08924_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08925_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08926_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08927_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08928_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08929_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08930_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08931_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08932_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08933_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08934_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08935_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08936_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08937_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08938_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08939_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08940_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08941_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08942_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08943_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08944_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08109_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08945_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08946_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08947_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08948_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08949_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08950_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08951_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08952_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08953_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08954_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08955_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08956_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08957_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08958_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08959_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08960_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08961_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08962_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08963_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08964_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08965_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08966_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08967_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08968_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08969_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08970_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08971_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08108_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08200_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00278_ ), .CK(_08107_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08199_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00279_ ), .CK(_08106_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08198_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00280_ ), .CK(_08105_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08972_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_08104_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08197_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00281_ ), .CK(_08103_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00282_ ), .CK(_08102_ ), .Q(\IF_ID_pc [30] ), .QN(_08196_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00283_ ), .CK(_08102_ ), .Q(\IF_ID_pc [21] ), .QN(_08195_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00284_ ), .CK(_08102_ ), .Q(\IF_ID_pc [20] ), .QN(_08194_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00285_ ), .CK(_08102_ ), .Q(\IF_ID_pc [19] ), .QN(_08193_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00286_ ), .CK(_08102_ ), .Q(\IF_ID_pc [18] ), .QN(_08192_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00287_ ), .CK(_08102_ ), .Q(\IF_ID_pc [17] ), .QN(_08191_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00288_ ), .CK(_08102_ ), .Q(\IF_ID_pc [16] ), .QN(_08190_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00289_ ), .CK(_08102_ ), .Q(\IF_ID_pc [15] ), .QN(_08189_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00290_ ), .CK(_08102_ ), .Q(\IF_ID_pc [14] ), .QN(_08188_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00291_ ), .CK(_08102_ ), .Q(\IF_ID_pc [13] ), .QN(_08187_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00292_ ), .CK(_08102_ ), .Q(\IF_ID_pc [12] ), .QN(_08186_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00293_ ), .CK(_08102_ ), .Q(\IF_ID_pc [29] ), .QN(_08185_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00294_ ), .CK(_08102_ ), .Q(\IF_ID_pc [11] ), .QN(_08184_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00295_ ), .CK(_08102_ ), .Q(\IF_ID_pc [10] ), .QN(_08183_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00296_ ), .CK(_08102_ ), .Q(\IF_ID_pc [9] ), .QN(_08182_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00297_ ), .CK(_08102_ ), .Q(\IF_ID_pc [8] ), .QN(_08181_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00298_ ), .CK(_08102_ ), .Q(\IF_ID_pc [7] ), .QN(_08180_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00299_ ), .CK(_08102_ ), .Q(\IF_ID_pc [6] ), .QN(_08179_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00300_ ), .CK(_08102_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00301_ ), .CK(_08102_ ), .Q(\IF_ID_pc [4] ), .QN(_08178_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00303_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08177_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00302_ ), .CK(_08102_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00305_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08175_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00304_ ), .CK(_08102_ ), .Q(\IF_ID_pc [2] ), .QN(_08176_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00306_ ), .CK(_08102_ ), .Q(\IF_ID_pc [28] ), .QN(_08174_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00307_ ), .CK(_08102_ ), .Q(\IF_ID_pc [1] ), .QN(_08173_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00308_ ), .CK(_08102_ ), .Q(\IF_ID_pc [27] ), .QN(_08172_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00309_ ), .CK(_08102_ ), .Q(\IF_ID_pc [26] ), .QN(_08171_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00310_ ), .CK(_08102_ ), .Q(\IF_ID_pc [25] ), .QN(_08170_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00311_ ), .CK(_08102_ ), .Q(\IF_ID_pc [24] ), .QN(_08169_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00312_ ), .CK(_08102_ ), .Q(\IF_ID_pc [23] ), .QN(_08168_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00313_ ), .CK(_08102_ ), .Q(\IF_ID_pc [22] ), .QN(_08167_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00314_ ), .CK(_08102_ ), .Q(\IF_ID_pc [31] ), .QN(_08166_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08974_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08165_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00315_ ), .CK(_08101_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08973_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00317_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00316_ ), .CK(_08100_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08164_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08975_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08976_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08977_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08978_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08979_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08980_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08981_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08982_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08983_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08984_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08985_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08986_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08987_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08988_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08989_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08990_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08991_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08992_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08993_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08994_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08995_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08996_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08997_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08998_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08999_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_09000_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_09001_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_09002_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_09003_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_09004_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_09005_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08099_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_09006_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_09007_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_09008_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_09009_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_09010_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_09011_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_09012_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_09013_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_09014_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_09015_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_09016_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_09017_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_09018_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_09019_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_09020_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_09021_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_09022_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_09023_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_09024_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_09025_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_09026_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_09027_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_09028_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_09029_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_09030_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_09031_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_09032_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_09033_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_09034_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_09035_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_09036_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_09037_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08098_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08163_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PN0P__Q ( .D(_00318_ ), .CK(_08097_ ), .Q(LS_WB_pc ), .QN(_08162_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PN0P__Q ( .D(_00319_ ), .CK(_08096_ ), .Q(\mylsu.previous_load_done ), .QN(_09038_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_09039_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_09040_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_09041_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(_09042_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_08099_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_08099_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_09043_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_08099_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08161_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00320_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08160_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00321_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08159_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00322_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08158_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00323_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08157_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00324_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08156_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00325_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08155_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00326_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08154_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00327_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08153_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00328_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08152_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00329_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08151_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00330_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08150_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00331_ ), .CK(_08099_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_09044_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_08099_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_09045_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_08099_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_09046_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_08099_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_09047_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_08099_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_09048_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_09049_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_09050_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_09051_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_09052_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_09053_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_09054_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_09055_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_09056_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_09057_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_09058_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_09059_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_09060_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_09061_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_09062_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_09063_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_09064_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_09065_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_09066_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_09067_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_09068_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_09069_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_09070_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_09071_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_09072_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_09073_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_09074_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_09075_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_09076_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_09077_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_09078_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_09079_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_08099_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_09080_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_09081_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_09082_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_09083_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_09084_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_09085_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_09086_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_09087_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_09088_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_09089_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_09090_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_09091_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_09092_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_09093_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_09094_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_09095_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_09096_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_09097_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_09098_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_09099_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_09100_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_09101_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_09102_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_09103_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_09104_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_09105_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_09106_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_09107_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_09108_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_09109_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_09110_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_09111_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_08095_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08149_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q ( .D(_00332_ ), .CK(_08094_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_08148_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_1 ( .D(_00333_ ), .CK(_08094_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08147_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_2 ( .D(_00334_ ), .CK(_08094_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08146_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_3 ( .D(_00335_ ), .CK(_08094_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08145_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_4 ( .D(_00336_ ), .CK(_08094_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08144_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_5 ( .D(_00337_ ), .CK(_08094_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08143_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PN0P__Q ( .D(_00338_ ), .CK(_08094_ ), .Q(LS_WB_wen_reg ), .QN(_09112_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_09113_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_09114_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08093_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08092_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08091_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08090_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08089_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08088_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08087_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08086_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08085_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08084_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08083_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08082_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08081_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08080_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08079_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_08078_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00339_ ), .CK(_08077_ ), .Q(loaduse_clear ), .QN(_09115_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_09116_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_09117_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08142_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(reset ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(excp_written ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_42 ) );

endmodule
