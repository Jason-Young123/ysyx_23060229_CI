//Generate the verilog at 2025-09-29T21:44:15 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire fc_disenable ;
wire io_master_awready_$_NOR__A_Y_$_OR__A_Y_$_OR__B_Y_$_ANDNOT__B_Y ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__B_A_$_ANDNOT__Y_A ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__B_Y_$_NOR__A_Y ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[0]_$_DFFE_PP__Q_E ;
wire \mycsreg.CSReg[1]_$_DFFE_PP__Q_E ;
wire \mycsreg.CSReg[2]_$_DFFE_PP__Q_E ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_E ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__A_Y ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__B_Y ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_B ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.inst_$_DFFE_PP__Q_10_D ;
wire \myifu.inst_$_DFFE_PP__Q_11_D ;
wire \myifu.inst_$_DFFE_PP__Q_12_D ;
wire \myifu.inst_$_DFFE_PP__Q_13_D ;
wire \myifu.inst_$_DFFE_PP__Q_14_D ;
wire \myifu.inst_$_DFFE_PP__Q_15_D ;
wire \myifu.inst_$_DFFE_PP__Q_16_D ;
wire \myifu.inst_$_DFFE_PP__Q_17_D ;
wire \myifu.inst_$_DFFE_PP__Q_18_D ;
wire \myifu.inst_$_DFFE_PP__Q_19_D ;
wire \myifu.inst_$_DFFE_PP__Q_1_D ;
wire \myifu.inst_$_DFFE_PP__Q_20_D ;
wire \myifu.inst_$_DFFE_PP__Q_21_D ;
wire \myifu.inst_$_DFFE_PP__Q_22_D ;
wire \myifu.inst_$_DFFE_PP__Q_23_D ;
wire \myifu.inst_$_DFFE_PP__Q_24_D ;
wire \myifu.inst_$_DFFE_PP__Q_25_D ;
wire \myifu.inst_$_DFFE_PP__Q_26_D ;
wire \myifu.inst_$_DFFE_PP__Q_27_D ;
wire \myifu.inst_$_DFFE_PP__Q_28_D ;
wire \myifu.inst_$_DFFE_PP__Q_29_D ;
wire \myifu.inst_$_DFFE_PP__Q_2_D ;
wire \myifu.inst_$_DFFE_PP__Q_30_D ;
wire \myifu.inst_$_DFFE_PP__Q_31_D ;
wire \myifu.inst_$_DFFE_PP__Q_3_D ;
wire \myifu.inst_$_DFFE_PP__Q_4_D ;
wire \myifu.inst_$_DFFE_PP__Q_5_D ;
wire \myifu.inst_$_DFFE_PP__Q_6_D ;
wire \myifu.inst_$_DFFE_PP__Q_7_D ;
wire \myifu.inst_$_DFFE_PP__Q_8_D ;
wire \myifu.inst_$_DFFE_PP__Q_9_D ;
wire \myifu.inst_$_DFFE_PP__Q_D ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_ORNOT__A_Y_$_NAND__A_Y_$_ANDNOT__B_Y ;
wire \myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_2_B_$_NOR__Y_B_$_OR__Y_B_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_Y ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_D ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_Y ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ORNOT__B_Y_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_D ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

INV_X1 _08668_ ( .A(fanout_net_1 ), .ZN(_01050_ ) );
BUF_X4 _08669_ ( .A(_01050_ ), .Z(_01051_ ) );
BUF_X2 _08670_ ( .A(_01051_ ), .Z(_01052_ ) );
AND3_X4 _08671_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01053_ ) );
AND3_X4 _08672_ ( .A1(_01053_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01054_ ) );
AND3_X4 _08673_ ( .A1(_01054_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01055_ ) );
AND3_X4 _08674_ ( .A1(_01055_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01056_ ) );
AND3_X4 _08675_ ( .A1(_01056_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01057_ ) );
AND3_X4 _08676_ ( .A1(_01057_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01058_ ) );
AND3_X4 _08677_ ( .A1(_01058_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01059_ ) );
AND3_X4 _08678_ ( .A1(_01059_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01060_ ) );
AND3_X4 _08679_ ( .A1(_01060_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01061_ ) );
AND3_X4 _08680_ ( .A1(_01061_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01062_ ) );
AND3_X4 _08681_ ( .A1(_01062_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01063_ ) );
AND3_X4 _08682_ ( .A1(_01063_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01064_ ) );
AND3_X4 _08683_ ( .A1(_01064_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01065_ ) );
AND2_X4 _08684_ ( .A1(_01065_ ), .A2(\myclint.mtime [27] ), .ZN(_01066_ ) );
AND2_X1 _08685_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01067_ ) );
AND2_X1 _08686_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01068_ ) );
AND4_X4 _08687_ ( .A1(\myclint.mtime [33] ), .A2(_01066_ ), .A3(_01067_ ), .A4(_01068_ ), .ZN(_01069_ ) );
AND3_X4 _08688_ ( .A1(_01069_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01070_ ) );
AND2_X4 _08689_ ( .A1(_01070_ ), .A2(\myclint.mtime [35] ), .ZN(_01071_ ) );
AND2_X1 _08690_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [39] ), .ZN(_01072_ ) );
AND2_X1 _08691_ ( .A1(\myclint.mtime [36] ), .A2(\myclint.mtime [37] ), .ZN(_01073_ ) );
AND3_X4 _08692_ ( .A1(_01071_ ), .A2(_01072_ ), .A3(_01073_ ), .ZN(_01074_ ) );
AND3_X4 _08693_ ( .A1(_01074_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01075_ ) );
AND2_X4 _08694_ ( .A1(_01075_ ), .A2(\myclint.mtime [42] ), .ZN(_01076_ ) );
AND2_X4 _08695_ ( .A1(_01076_ ), .A2(\myclint.mtime [43] ), .ZN(_01077_ ) );
AND2_X1 _08696_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01078_ ) );
AND3_X1 _08697_ ( .A1(_01078_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01079_ ) );
NAND2_X4 _08698_ ( .A1(_01077_ ), .A2(_01079_ ), .ZN(_01080_ ) );
AND2_X1 _08699_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01081_ ) );
INV_X1 _08700_ ( .A(_01081_ ), .ZN(_01082_ ) );
NOR2_X4 _08701_ ( .A1(_01080_ ), .A2(_01082_ ), .ZN(_01083_ ) );
AND2_X1 _08702_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01084_ ) );
AND2_X2 _08703_ ( .A1(_01083_ ), .A2(_01084_ ), .ZN(_01085_ ) );
AND2_X1 _08704_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01086_ ) );
AND2_X2 _08705_ ( .A1(_01085_ ), .A2(_01086_ ), .ZN(_01087_ ) );
AND2_X1 _08706_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01088_ ) );
AND2_X2 _08707_ ( .A1(_01087_ ), .A2(_01088_ ), .ZN(_01089_ ) );
AND2_X1 _08708_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01090_ ) );
AND2_X2 _08709_ ( .A1(_01089_ ), .A2(_01090_ ), .ZN(_01091_ ) );
AND2_X1 _08710_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01092_ ) );
AND2_X4 _08711_ ( .A1(_01091_ ), .A2(_01092_ ), .ZN(_01093_ ) );
NAND3_X4 _08712_ ( .A1(_01093_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01094_ ) );
NOR2_X2 _08713_ ( .A1(_01094_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01095_ ) );
OAI21_X1 _08714_ ( .A(_01052_ ), .B1(_01095_ ), .B2(\myclint.mtime [63] ), .ZN(_01096_ ) );
AND3_X4 _08715_ ( .A1(_01065_ ), .A2(\myclint.mtime [28] ), .A3(\myclint.mtime [27] ), .ZN(_01097_ ) );
AND2_X4 _08716_ ( .A1(_01097_ ), .A2(\myclint.mtime [29] ), .ZN(_01098_ ) );
AND2_X1 _08717_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01099_ ) );
AND3_X2 _08718_ ( .A1(_01098_ ), .A2(_01099_ ), .A3(_01067_ ), .ZN(_01100_ ) );
AND2_X4 _08719_ ( .A1(_01100_ ), .A2(\myclint.mtime [34] ), .ZN(_01101_ ) );
AND2_X4 _08720_ ( .A1(_01101_ ), .A2(\myclint.mtime [35] ), .ZN(_01102_ ) );
AND3_X2 _08721_ ( .A1(_01102_ ), .A2(_01072_ ), .A3(_01073_ ), .ZN(_01103_ ) );
NAND2_X4 _08722_ ( .A1(_01103_ ), .A2(\myclint.mtime [40] ), .ZN(_01104_ ) );
INV_X1 _08723_ ( .A(\myclint.mtime [42] ), .ZN(_01105_ ) );
INV_X1 _08724_ ( .A(\myclint.mtime [41] ), .ZN(_01106_ ) );
NOR3_X4 _08725_ ( .A1(_01104_ ), .A2(_01105_ ), .A3(_01106_ ), .ZN(_01107_ ) );
AND2_X4 _08726_ ( .A1(_01107_ ), .A2(\myclint.mtime [43] ), .ZN(_01108_ ) );
AND2_X2 _08727_ ( .A1(_01108_ ), .A2(_01079_ ), .ZN(_01109_ ) );
AND2_X4 _08728_ ( .A1(_01109_ ), .A2(_01081_ ), .ZN(_01110_ ) );
AND2_X2 _08729_ ( .A1(_01110_ ), .A2(_01084_ ), .ZN(_01111_ ) );
AND2_X2 _08730_ ( .A1(_01111_ ), .A2(_01086_ ), .ZN(_01112_ ) );
AND2_X2 _08731_ ( .A1(_01112_ ), .A2(_01088_ ), .ZN(_01113_ ) );
AND2_X2 _08732_ ( .A1(_01113_ ), .A2(_01090_ ), .ZN(_01114_ ) );
AND2_X2 _08733_ ( .A1(_01114_ ), .A2(_01092_ ), .ZN(_01115_ ) );
NAND3_X1 _08734_ ( .A1(_01115_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01116_ ) );
NOR2_X1 _08735_ ( .A1(_01116_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01117_ ) );
AOI21_X1 _08736_ ( .A(_01096_ ), .B1(\myclint.mtime [63] ), .B2(_01117_ ), .ZN(_00000_ ) );
AND2_X1 _08737_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_01118_ ) );
AND3_X1 _08738_ ( .A1(_01118_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01119_ ) );
AND4_X1 _08739_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01120_ ) );
AND2_X1 _08740_ ( .A1(_01119_ ), .A2(_01120_ ), .ZN(_01121_ ) );
AND2_X1 _08741_ ( .A1(\myclint.mtime [24] ), .A2(\myclint.mtime [25] ), .ZN(_01122_ ) );
AND3_X1 _08742_ ( .A1(_01122_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [27] ), .ZN(_01123_ ) );
AND4_X1 _08743_ ( .A1(_01067_ ), .A2(_01121_ ), .A3(_01068_ ), .A4(_01123_ ), .ZN(_01124_ ) );
AND2_X1 _08744_ ( .A1(_01053_ ), .A2(\myclint.mtime [3] ), .ZN(_01125_ ) );
AND4_X1 _08745_ ( .A1(\myclint.mtime [6] ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [5] ), .A4(\myclint.mtime [7] ), .ZN(_01126_ ) );
AND2_X1 _08746_ ( .A1(_01125_ ), .A2(_01126_ ), .ZN(_01127_ ) );
AND4_X1 _08747_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01128_ ) );
AND2_X1 _08748_ ( .A1(\myclint.mtime [10] ), .A2(\myclint.mtime [11] ), .ZN(_01129_ ) );
AND4_X1 _08749_ ( .A1(\myclint.mtime [8] ), .A2(_01128_ ), .A3(\myclint.mtime [9] ), .A4(_01129_ ), .ZN(_01130_ ) );
AND2_X2 _08750_ ( .A1(_01127_ ), .A2(_01130_ ), .ZN(_01131_ ) );
AND2_X1 _08751_ ( .A1(_01124_ ), .A2(_01131_ ), .ZN(_01132_ ) );
AND3_X1 _08752_ ( .A1(_01099_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01133_ ) );
AND3_X1 _08753_ ( .A1(_01133_ ), .A2(_01072_ ), .A3(_01073_ ), .ZN(_01134_ ) );
AND2_X1 _08754_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01135_ ) );
AND3_X1 _08755_ ( .A1(_01135_ ), .A2(\myclint.mtime [42] ), .A3(\myclint.mtime [43] ), .ZN(_01136_ ) );
AND3_X1 _08756_ ( .A1(_01134_ ), .A2(_01079_ ), .A3(_01136_ ), .ZN(_01137_ ) );
AND2_X1 _08757_ ( .A1(_01132_ ), .A2(_01137_ ), .ZN(_01138_ ) );
AND4_X1 _08758_ ( .A1(_01088_ ), .A2(_01086_ ), .A3(_01084_ ), .A4(_01081_ ), .ZN(_01139_ ) );
AND2_X1 _08759_ ( .A1(_01138_ ), .A2(_01139_ ), .ZN(_01140_ ) );
AND4_X1 _08760_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01141_ ) );
AND2_X1 _08761_ ( .A1(_01140_ ), .A2(_01141_ ), .ZN(_01142_ ) );
AND3_X1 _08762_ ( .A1(_01142_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01143_ ) );
XNOR2_X1 _08763_ ( .A(_01143_ ), .B(\myclint.mtime [62] ), .ZN(_01144_ ) );
NOR2_X1 _08764_ ( .A1(_01144_ ), .A2(fanout_net_1 ), .ZN(_00001_ ) );
INV_X1 _08765_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01145_ ) );
AND4_X1 _08766_ ( .A1(_01145_ ), .A2(_01110_ ), .A3(\myclint.mtime [53] ), .A4(_01084_ ), .ZN(_01146_ ) );
BUF_X4 _08767_ ( .A(_01051_ ), .Z(_01147_ ) );
BUF_X2 _08768_ ( .A(_01147_ ), .Z(_01148_ ) );
AND3_X1 _08769_ ( .A1(_01083_ ), .A2(_01145_ ), .A3(_01084_ ), .ZN(_01149_ ) );
OAI21_X1 _08770_ ( .A(_01148_ ), .B1(_01149_ ), .B2(\myclint.mtime [53] ), .ZN(_01150_ ) );
NOR2_X1 _08771_ ( .A1(_01146_ ), .A2(_01150_ ), .ZN(_00002_ ) );
AND2_X1 _08772_ ( .A1(_01084_ ), .A2(_01081_ ), .ZN(_01151_ ) );
AND2_X1 _08773_ ( .A1(_01138_ ), .A2(_01151_ ), .ZN(_01152_ ) );
XNOR2_X1 _08774_ ( .A(_01152_ ), .B(\myclint.mtime [52] ), .ZN(_01153_ ) );
NOR2_X1 _08775_ ( .A1(_01153_ ), .A2(fanout_net_1 ), .ZN(_00003_ ) );
NOR3_X1 _08776_ ( .A1(_01080_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01082_ ), .ZN(_01154_ ) );
OAI21_X1 _08777_ ( .A(_01052_ ), .B1(_01154_ ), .B2(\myclint.mtime [51] ), .ZN(_01155_ ) );
INV_X1 _08778_ ( .A(_01109_ ), .ZN(_01156_ ) );
NOR3_X1 _08779_ ( .A1(_01156_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01082_ ), .ZN(_01157_ ) );
AOI21_X1 _08780_ ( .A(_01155_ ), .B1(_01157_ ), .B2(\myclint.mtime [51] ), .ZN(_00004_ ) );
INV_X1 _08781_ ( .A(_01132_ ), .ZN(_01158_ ) );
INV_X1 _08782_ ( .A(_01137_ ), .ZN(_01159_ ) );
OR4_X1 _08783_ ( .A1(\myclint.mtime [50] ), .A2(_01158_ ), .A3(_01082_ ), .A4(_01159_ ), .ZN(_01160_ ) );
AND3_X1 _08784_ ( .A1(_01132_ ), .A2(_01081_ ), .A3(_01137_ ), .ZN(_01161_ ) );
INV_X1 _08785_ ( .A(_01161_ ), .ZN(_01162_ ) );
NAND2_X1 _08786_ ( .A1(_01162_ ), .A2(\myclint.mtime [50] ), .ZN(_01163_ ) );
AOI21_X1 _08787_ ( .A(fanout_net_1 ), .B1(_01160_ ), .B2(_01163_ ), .ZN(_00005_ ) );
INV_X1 _08788_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01164_ ) );
AND4_X1 _08789_ ( .A1(\myclint.mtime [49] ), .A2(_01108_ ), .A3(_01164_ ), .A4(_01079_ ), .ZN(_01165_ ) );
AND3_X1 _08790_ ( .A1(_01077_ ), .A2(_01164_ ), .A3(_01079_ ), .ZN(_01166_ ) );
OAI21_X1 _08791_ ( .A(_01148_ ), .B1(_01166_ ), .B2(\myclint.mtime [49] ), .ZN(_01167_ ) );
NOR2_X1 _08792_ ( .A1(_01165_ ), .A2(_01167_ ), .ZN(_00006_ ) );
INV_X1 _08793_ ( .A(_01124_ ), .ZN(_01168_ ) );
INV_X1 _08794_ ( .A(_01131_ ), .ZN(_01169_ ) );
OR4_X1 _08795_ ( .A1(\myclint.mtime [48] ), .A2(_01168_ ), .A3(_01159_ ), .A4(_01169_ ), .ZN(_01170_ ) );
OAI21_X1 _08796_ ( .A(\myclint.mtime [48] ), .B1(_01158_ ), .B2(_01159_ ), .ZN(_01171_ ) );
AOI21_X1 _08797_ ( .A(fanout_net_1 ), .B1(_01170_ ), .B2(_01171_ ), .ZN(_00007_ ) );
NAND3_X1 _08798_ ( .A1(_01076_ ), .A2(\myclint.mtime [43] ), .A3(_01078_ ), .ZN(_01172_ ) );
NOR2_X1 _08799_ ( .A1(_01172_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01173_ ) );
OAI21_X1 _08800_ ( .A(_01052_ ), .B1(_01173_ ), .B2(\myclint.mtime [47] ), .ZN(_01174_ ) );
NAND3_X1 _08801_ ( .A1(_01107_ ), .A2(\myclint.mtime [44] ), .A3(\myclint.mtime [43] ), .ZN(_01175_ ) );
INV_X1 _08802_ ( .A(\myclint.mtime [45] ), .ZN(_01176_ ) );
NOR3_X1 _08803_ ( .A1(_01175_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01176_ ), .ZN(_01177_ ) );
AOI21_X1 _08804_ ( .A(_01174_ ), .B1(_01177_ ), .B2(\myclint.mtime [47] ), .ZN(_00008_ ) );
AND2_X1 _08805_ ( .A1(_01132_ ), .A2(_01134_ ), .ZN(_01178_ ) );
AND3_X1 _08806_ ( .A1(_01178_ ), .A2(_01078_ ), .A3(_01136_ ), .ZN(_01179_ ) );
XNOR2_X1 _08807_ ( .A(_01179_ ), .B(\myclint.mtime [46] ), .ZN(_01180_ ) );
NOR2_X1 _08808_ ( .A1(_01180_ ), .A2(fanout_net_1 ), .ZN(_00009_ ) );
INV_X1 _08809_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01181_ ) );
NAND3_X1 _08810_ ( .A1(_01076_ ), .A2(_01181_ ), .A3(\myclint.mtime [43] ), .ZN(_01182_ ) );
AOI21_X1 _08811_ ( .A(fanout_net_1 ), .B1(_01182_ ), .B2(_01176_ ), .ZN(_01183_ ) );
NAND4_X1 _08812_ ( .A1(_01107_ ), .A2(\myclint.mtime [45] ), .A3(_01181_ ), .A4(\myclint.mtime [43] ), .ZN(_01184_ ) );
AND2_X1 _08813_ ( .A1(_01183_ ), .A2(_01184_ ), .ZN(_00010_ ) );
AND2_X1 _08814_ ( .A1(_01178_ ), .A2(_01136_ ), .ZN(_01185_ ) );
XNOR2_X1 _08815_ ( .A(_01185_ ), .B(\myclint.mtime [44] ), .ZN(_01186_ ) );
NOR2_X1 _08816_ ( .A1(_01186_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
INV_X1 _08817_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01187_ ) );
AND4_X1 _08818_ ( .A1(\myclint.mtime [61] ), .A2(_01114_ ), .A3(_01187_ ), .A4(_01092_ ), .ZN(_01188_ ) );
AND3_X1 _08819_ ( .A1(_01091_ ), .A2(_01187_ ), .A3(_01092_ ), .ZN(_01189_ ) );
OAI21_X1 _08820_ ( .A(_01148_ ), .B1(_01189_ ), .B2(\myclint.mtime [61] ), .ZN(_01190_ ) );
NOR2_X1 _08821_ ( .A1(_01188_ ), .A2(_01190_ ), .ZN(_00012_ ) );
BUF_X4 _08822_ ( .A(_01147_ ), .Z(_01191_ ) );
INV_X1 _08823_ ( .A(_01075_ ), .ZN(_01192_ ) );
NOR2_X1 _08824_ ( .A1(_01192_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01193_ ) );
OAI21_X1 _08825_ ( .A(_01191_ ), .B1(_01193_ ), .B2(\myclint.mtime [43] ), .ZN(_01194_ ) );
NOR3_X1 _08826_ ( .A1(_01104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01106_ ), .ZN(_01195_ ) );
AOI21_X1 _08827_ ( .A(_01194_ ), .B1(_01195_ ), .B2(\myclint.mtime [43] ), .ZN(_00013_ ) );
OAI21_X1 _08828_ ( .A(_01148_ ), .B1(_01075_ ), .B2(\myclint.mtime [42] ), .ZN(_01196_ ) );
NOR2_X1 _08829_ ( .A1(_01076_ ), .A2(_01196_ ), .ZN(_00014_ ) );
INV_X1 _08830_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01197_ ) );
NAND2_X1 _08831_ ( .A1(_01074_ ), .A2(_01197_ ), .ZN(_01198_ ) );
AOI21_X1 _08832_ ( .A(fanout_net_1 ), .B1(_01198_ ), .B2(_01106_ ), .ZN(_01199_ ) );
AND2_X1 _08833_ ( .A1(_01102_ ), .A2(_01073_ ), .ZN(_01200_ ) );
NAND4_X1 _08834_ ( .A1(_01200_ ), .A2(\myclint.mtime [41] ), .A3(_01197_ ), .A4(_01072_ ), .ZN(_01201_ ) );
AND2_X1 _08835_ ( .A1(_01199_ ), .A2(_01201_ ), .ZN(_00015_ ) );
XNOR2_X1 _08836_ ( .A(_01178_ ), .B(\myclint.mtime [40] ), .ZN(_01202_ ) );
NOR2_X1 _08837_ ( .A1(_01202_ ), .A2(fanout_net_1 ), .ZN(_00016_ ) );
NAND3_X1 _08838_ ( .A1(_01132_ ), .A2(_01073_ ), .A3(_01133_ ), .ZN(_01203_ ) );
OR3_X1 _08839_ ( .A1(_01203_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [39] ), .ZN(_01204_ ) );
OAI21_X1 _08840_ ( .A(\myclint.mtime [39] ), .B1(_01203_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01205_ ) );
AOI21_X1 _08841_ ( .A(fanout_net_1 ), .B1(_01204_ ), .B2(_01205_ ), .ZN(_00017_ ) );
OR2_X1 _08842_ ( .A1(_01203_ ), .A2(\myclint.mtime [38] ), .ZN(_01206_ ) );
NAND2_X1 _08843_ ( .A1(_01203_ ), .A2(\myclint.mtime [38] ), .ZN(_01207_ ) );
AOI21_X1 _08844_ ( .A(fanout_net_1 ), .B1(_01206_ ), .B2(_01207_ ), .ZN(_00018_ ) );
INV_X1 _08845_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01208_ ) );
AND4_X1 _08846_ ( .A1(\myclint.mtime [37] ), .A2(_01101_ ), .A3(_01208_ ), .A4(\myclint.mtime [35] ), .ZN(_01209_ ) );
AND3_X1 _08847_ ( .A1(_01070_ ), .A2(_01208_ ), .A3(\myclint.mtime [35] ), .ZN(_01210_ ) );
OAI21_X1 _08848_ ( .A(_01148_ ), .B1(_01210_ ), .B2(\myclint.mtime [37] ), .ZN(_01211_ ) );
NOR2_X1 _08849_ ( .A1(_01209_ ), .A2(_01211_ ), .ZN(_00019_ ) );
AND2_X1 _08850_ ( .A1(_01132_ ), .A2(_01133_ ), .ZN(_01212_ ) );
XNOR2_X1 _08851_ ( .A(_01212_ ), .B(\myclint.mtime [36] ), .ZN(_01213_ ) );
NOR2_X1 _08852_ ( .A1(_01213_ ), .A2(fanout_net_1 ), .ZN(_00020_ ) );
NAND3_X1 _08853_ ( .A1(_01124_ ), .A2(_01099_ ), .A3(_01131_ ), .ZN(_01214_ ) );
OR3_X1 _08854_ ( .A1(_01214_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [35] ), .ZN(_01215_ ) );
OAI21_X1 _08855_ ( .A(\myclint.mtime [35] ), .B1(_01214_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01216_ ) );
AOI21_X1 _08856_ ( .A(fanout_net_1 ), .B1(_01215_ ), .B2(_01216_ ), .ZN(_00021_ ) );
BUF_X2 _08857_ ( .A(_01147_ ), .Z(_01217_ ) );
NAND4_X1 _08858_ ( .A1(_01066_ ), .A2(\myclint.mtime [33] ), .A3(_01067_ ), .A4(_01068_ ), .ZN(_01218_ ) );
INV_X1 _08859_ ( .A(\myclint.mtime [32] ), .ZN(_01219_ ) );
NOR2_X1 _08860_ ( .A1(_01218_ ), .A2(_01219_ ), .ZN(_01220_ ) );
OAI21_X1 _08861_ ( .A(_01217_ ), .B1(_01220_ ), .B2(\myclint.mtime [34] ), .ZN(_01221_ ) );
NOR2_X1 _08862_ ( .A1(_01221_ ), .A2(_01070_ ), .ZN(_00022_ ) );
XNOR2_X1 _08863_ ( .A(_01142_ ), .B(\myclint.mtime [60] ), .ZN(_01222_ ) );
NOR2_X1 _08864_ ( .A1(_01222_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
AND2_X1 _08865_ ( .A1(_01066_ ), .A2(_01068_ ), .ZN(_01223_ ) );
INV_X1 _08866_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01224_ ) );
AND3_X1 _08867_ ( .A1(_01223_ ), .A2(_01224_ ), .A3(_01067_ ), .ZN(_01225_ ) );
OAI21_X1 _08868_ ( .A(_01217_ ), .B1(_01225_ ), .B2(\myclint.mtime [33] ), .ZN(_01226_ ) );
AND4_X1 _08869_ ( .A1(_01224_ ), .A2(_01098_ ), .A3(\myclint.mtime [33] ), .A4(_01067_ ), .ZN(_01227_ ) );
NOR2_X1 _08870_ ( .A1(_01226_ ), .A2(_01227_ ), .ZN(_00024_ ) );
OAI21_X1 _08871_ ( .A(\myclint.mtime [32] ), .B1(_01168_ ), .B2(_01169_ ), .ZN(_01228_ ) );
NAND3_X1 _08872_ ( .A1(_01124_ ), .A2(_01219_ ), .A3(_01131_ ), .ZN(_01229_ ) );
AOI21_X1 _08873_ ( .A(fanout_net_1 ), .B1(_01228_ ), .B2(_01229_ ), .ZN(_00025_ ) );
INV_X1 _08874_ ( .A(_01097_ ), .ZN(_01230_ ) );
INV_X1 _08875_ ( .A(\myclint.mtime [29] ), .ZN(_01231_ ) );
NOR3_X1 _08876_ ( .A1(_01230_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01231_ ), .ZN(_01232_ ) );
AND2_X1 _08877_ ( .A1(_01232_ ), .A2(\myclint.mtime [31] ), .ZN(_01233_ ) );
OAI21_X1 _08878_ ( .A(_01148_ ), .B1(_01232_ ), .B2(\myclint.mtime [31] ), .ZN(_01234_ ) );
NOR2_X1 _08879_ ( .A1(_01233_ ), .A2(_01234_ ), .ZN(_00026_ ) );
AND2_X1 _08880_ ( .A1(_01131_ ), .A2(_01121_ ), .ZN(_01235_ ) );
NAND3_X1 _08881_ ( .A1(_01235_ ), .A2(_01068_ ), .A3(_01123_ ), .ZN(_01236_ ) );
OR2_X1 _08882_ ( .A1(_01236_ ), .A2(\myclint.mtime [30] ), .ZN(_01237_ ) );
NAND2_X1 _08883_ ( .A1(_01236_ ), .A2(\myclint.mtime [30] ), .ZN(_01238_ ) );
AOI21_X1 _08884_ ( .A(fanout_net_1 ), .B1(_01237_ ), .B2(_01238_ ), .ZN(_00027_ ) );
INV_X1 _08885_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01239_ ) );
AND3_X1 _08886_ ( .A1(_01065_ ), .A2(_01239_ ), .A3(\myclint.mtime [27] ), .ZN(_01240_ ) );
AND2_X1 _08887_ ( .A1(_01240_ ), .A2(\myclint.mtime [29] ), .ZN(_01241_ ) );
BUF_X2 _08888_ ( .A(_01147_ ), .Z(_01242_ ) );
OAI21_X1 _08889_ ( .A(_01242_ ), .B1(_01240_ ), .B2(\myclint.mtime [29] ), .ZN(_01243_ ) );
NOR2_X1 _08890_ ( .A1(_01241_ ), .A2(_01243_ ), .ZN(_00028_ ) );
NAND2_X1 _08891_ ( .A1(_01235_ ), .A2(_01123_ ), .ZN(_01244_ ) );
XNOR2_X1 _08892_ ( .A(_01244_ ), .B(\myclint.mtime [28] ), .ZN(_01245_ ) );
CLKBUF_X2 _08893_ ( .A(_01147_ ), .Z(_01246_ ) );
AND2_X1 _08894_ ( .A1(_01245_ ), .A2(_01246_ ), .ZN(_00029_ ) );
NAND3_X1 _08895_ ( .A1(_01131_ ), .A2(_01122_ ), .A3(_01121_ ), .ZN(_01247_ ) );
OR3_X1 _08896_ ( .A1(_01247_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01248_ ) );
OAI21_X1 _08897_ ( .A(\myclint.mtime [27] ), .B1(_01247_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01249_ ) );
AOI21_X1 _08898_ ( .A(fanout_net_1 ), .B1(_01248_ ), .B2(_01249_ ), .ZN(_00030_ ) );
AND2_X1 _08899_ ( .A1(_01064_ ), .A2(\myclint.mtime [25] ), .ZN(_01250_ ) );
OAI21_X1 _08900_ ( .A(_01217_ ), .B1(_01250_ ), .B2(\myclint.mtime [26] ), .ZN(_01251_ ) );
NOR2_X1 _08901_ ( .A1(_01251_ ), .A2(_01065_ ), .ZN(_00031_ ) );
INV_X1 _08902_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01252_ ) );
AND3_X1 _08903_ ( .A1(_01063_ ), .A2(_01252_ ), .A3(\myclint.mtime [23] ), .ZN(_01253_ ) );
AND2_X1 _08904_ ( .A1(_01253_ ), .A2(\myclint.mtime [25] ), .ZN(_01254_ ) );
OAI21_X1 _08905_ ( .A(_01242_ ), .B1(_01253_ ), .B2(\myclint.mtime [25] ), .ZN(_01255_ ) );
NOR2_X1 _08906_ ( .A1(_01254_ ), .A2(_01255_ ), .ZN(_00032_ ) );
AND2_X1 _08907_ ( .A1(_01063_ ), .A2(\myclint.mtime [23] ), .ZN(_01256_ ) );
OAI21_X1 _08908_ ( .A(_01217_ ), .B1(_01256_ ), .B2(\myclint.mtime [24] ), .ZN(_01257_ ) );
NOR2_X1 _08909_ ( .A1(_01257_ ), .A2(_01064_ ), .ZN(_00033_ ) );
NAND3_X1 _08910_ ( .A1(_01138_ ), .A2(_01090_ ), .A3(_01139_ ), .ZN(_01258_ ) );
OR3_X1 _08911_ ( .A1(_01258_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [59] ), .ZN(_01259_ ) );
OAI21_X1 _08912_ ( .A(\myclint.mtime [59] ), .B1(_01258_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01260_ ) );
AOI21_X1 _08913_ ( .A(fanout_net_1 ), .B1(_01259_ ), .B2(_01260_ ), .ZN(_00034_ ) );
AND2_X1 _08914_ ( .A1(_01131_ ), .A2(_01119_ ), .ZN(_01261_ ) );
NAND3_X1 _08915_ ( .A1(_01261_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01262_ ) );
OR3_X1 _08916_ ( .A1(_01262_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01263_ ) );
OAI21_X1 _08917_ ( .A(\myclint.mtime [23] ), .B1(_01262_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01264_ ) );
AOI21_X1 _08918_ ( .A(fanout_net_1 ), .B1(_01263_ ), .B2(_01264_ ), .ZN(_00035_ ) );
BUF_X4 _08919_ ( .A(_01147_ ), .Z(_01265_ ) );
AND2_X1 _08920_ ( .A1(_01062_ ), .A2(\myclint.mtime [21] ), .ZN(_01266_ ) );
OAI21_X1 _08921_ ( .A(_01265_ ), .B1(_01266_ ), .B2(\myclint.mtime [22] ), .ZN(_01267_ ) );
NOR2_X1 _08922_ ( .A1(_01267_ ), .A2(_01063_ ), .ZN(_00036_ ) );
INV_X1 _08923_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01268_ ) );
AND3_X1 _08924_ ( .A1(_01061_ ), .A2(_01268_ ), .A3(\myclint.mtime [19] ), .ZN(_01269_ ) );
AND2_X1 _08925_ ( .A1(_01269_ ), .A2(\myclint.mtime [21] ), .ZN(_01270_ ) );
OAI21_X1 _08926_ ( .A(_01242_ ), .B1(_01269_ ), .B2(\myclint.mtime [21] ), .ZN(_01271_ ) );
NOR2_X1 _08927_ ( .A1(_01270_ ), .A2(_01271_ ), .ZN(_00037_ ) );
AND2_X1 _08928_ ( .A1(_01061_ ), .A2(\myclint.mtime [19] ), .ZN(_01272_ ) );
OAI21_X1 _08929_ ( .A(_01265_ ), .B1(_01272_ ), .B2(\myclint.mtime [20] ), .ZN(_01273_ ) );
NOR2_X1 _08930_ ( .A1(_01273_ ), .A2(_01062_ ), .ZN(_00038_ ) );
NAND3_X1 _08931_ ( .A1(_01131_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01274_ ) );
OR3_X1 _08932_ ( .A1(_01274_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01275_ ) );
OAI21_X1 _08933_ ( .A(\myclint.mtime [19] ), .B1(_01274_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01276_ ) );
AOI21_X1 _08934_ ( .A(fanout_net_1 ), .B1(_01275_ ), .B2(_01276_ ), .ZN(_00039_ ) );
AND2_X1 _08935_ ( .A1(_01060_ ), .A2(\myclint.mtime [17] ), .ZN(_01277_ ) );
OAI21_X1 _08936_ ( .A(_01265_ ), .B1(_01277_ ), .B2(\myclint.mtime [18] ), .ZN(_01278_ ) );
NOR2_X1 _08937_ ( .A1(_01278_ ), .A2(_01061_ ), .ZN(_00040_ ) );
INV_X1 _08938_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01279_ ) );
AND3_X1 _08939_ ( .A1(_01059_ ), .A2(_01279_ ), .A3(\myclint.mtime [15] ), .ZN(_01280_ ) );
AND2_X1 _08940_ ( .A1(_01280_ ), .A2(\myclint.mtime [17] ), .ZN(_01281_ ) );
OAI21_X1 _08941_ ( .A(_01242_ ), .B1(_01280_ ), .B2(\myclint.mtime [17] ), .ZN(_01282_ ) );
NOR2_X1 _08942_ ( .A1(_01281_ ), .A2(_01282_ ), .ZN(_00041_ ) );
AND2_X1 _08943_ ( .A1(_01059_ ), .A2(\myclint.mtime [15] ), .ZN(_01283_ ) );
OAI21_X1 _08944_ ( .A(_01265_ ), .B1(_01283_ ), .B2(\myclint.mtime [16] ), .ZN(_01284_ ) );
NOR2_X1 _08945_ ( .A1(_01284_ ), .A2(_01060_ ), .ZN(_00042_ ) );
AND3_X1 _08946_ ( .A1(_01129_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01285_ ) );
AND2_X1 _08947_ ( .A1(_01127_ ), .A2(_01285_ ), .ZN(_01286_ ) );
NAND3_X1 _08948_ ( .A1(_01286_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01287_ ) );
OR3_X1 _08949_ ( .A1(_01287_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01288_ ) );
OAI21_X1 _08950_ ( .A(\myclint.mtime [15] ), .B1(_01287_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01289_ ) );
AOI21_X1 _08951_ ( .A(fanout_net_1 ), .B1(_01288_ ), .B2(_01289_ ), .ZN(_00043_ ) );
AND2_X1 _08952_ ( .A1(_01058_ ), .A2(\myclint.mtime [13] ), .ZN(_01290_ ) );
OAI21_X1 _08953_ ( .A(_01265_ ), .B1(_01290_ ), .B2(\myclint.mtime [14] ), .ZN(_01291_ ) );
NOR2_X1 _08954_ ( .A1(_01291_ ), .A2(_01059_ ), .ZN(_00044_ ) );
OR2_X1 _08955_ ( .A1(_01258_ ), .A2(\myclint.mtime [58] ), .ZN(_01292_ ) );
NAND2_X1 _08956_ ( .A1(_01258_ ), .A2(\myclint.mtime [58] ), .ZN(_01293_ ) );
AOI21_X1 _08957_ ( .A(fanout_net_1 ), .B1(_01292_ ), .B2(_01293_ ), .ZN(_00045_ ) );
INV_X1 _08958_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01294_ ) );
AND3_X1 _08959_ ( .A1(_01057_ ), .A2(_01294_ ), .A3(\myclint.mtime [11] ), .ZN(_01295_ ) );
AND2_X1 _08960_ ( .A1(_01295_ ), .A2(\myclint.mtime [13] ), .ZN(_01296_ ) );
OAI21_X1 _08961_ ( .A(_01242_ ), .B1(_01295_ ), .B2(\myclint.mtime [13] ), .ZN(_01297_ ) );
NOR2_X1 _08962_ ( .A1(_01296_ ), .A2(_01297_ ), .ZN(_00046_ ) );
AND2_X1 _08963_ ( .A1(_01057_ ), .A2(\myclint.mtime [11] ), .ZN(_01298_ ) );
OAI21_X1 _08964_ ( .A(_01265_ ), .B1(_01298_ ), .B2(\myclint.mtime [12] ), .ZN(_01299_ ) );
NOR2_X1 _08965_ ( .A1(_01299_ ), .A2(_01058_ ), .ZN(_00047_ ) );
NAND3_X1 _08966_ ( .A1(_01127_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01300_ ) );
OR3_X1 _08967_ ( .A1(_01300_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_01301_ ) );
OAI21_X1 _08968_ ( .A(\myclint.mtime [11] ), .B1(_01300_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01302_ ) );
AOI21_X1 _08969_ ( .A(fanout_net_1 ), .B1(_01301_ ), .B2(_01302_ ), .ZN(_00048_ ) );
AND2_X1 _08970_ ( .A1(_01056_ ), .A2(\myclint.mtime [9] ), .ZN(_01303_ ) );
OAI21_X1 _08971_ ( .A(_01265_ ), .B1(_01303_ ), .B2(\myclint.mtime [10] ), .ZN(_01304_ ) );
NOR2_X1 _08972_ ( .A1(_01304_ ), .A2(_01057_ ), .ZN(_00049_ ) );
AND2_X1 _08973_ ( .A1(_01055_ ), .A2(\myclint.mtime [7] ), .ZN(_01305_ ) );
INV_X1 _08974_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01306_ ) );
AND3_X1 _08975_ ( .A1(_01305_ ), .A2(\myclint.mtime [9] ), .A3(_01306_ ), .ZN(_01307_ ) );
AOI21_X1 _08976_ ( .A(\myclint.mtime [9] ), .B1(_01305_ ), .B2(_01306_ ), .ZN(_01308_ ) );
NOR3_X1 _08977_ ( .A1(_01307_ ), .A2(_01308_ ), .A3(fanout_net_1 ), .ZN(_00050_ ) );
OAI21_X1 _08978_ ( .A(_01265_ ), .B1(_01305_ ), .B2(\myclint.mtime [8] ), .ZN(_01309_ ) );
NOR2_X1 _08979_ ( .A1(_01309_ ), .A2(_01056_ ), .ZN(_00051_ ) );
AND2_X1 _08980_ ( .A1(_01054_ ), .A2(\myclint.mtime [5] ), .ZN(_01310_ ) );
INV_X1 _08981_ ( .A(_01310_ ), .ZN(_01311_ ) );
OR3_X1 _08982_ ( .A1(_01311_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [7] ), .ZN(_01312_ ) );
OAI21_X1 _08983_ ( .A(\myclint.mtime [7] ), .B1(_01311_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01313_ ) );
AOI21_X1 _08984_ ( .A(fanout_net_1 ), .B1(_01312_ ), .B2(_01313_ ), .ZN(_00052_ ) );
OAI21_X1 _08985_ ( .A(_01265_ ), .B1(_01310_ ), .B2(\myclint.mtime [6] ), .ZN(_01314_ ) );
NOR2_X1 _08986_ ( .A1(_01314_ ), .A2(_01055_ ), .ZN(_00053_ ) );
INV_X1 _08987_ ( .A(_01125_ ), .ZN(_01315_ ) );
OR3_X1 _08988_ ( .A1(_01315_ ), .A2(\myclint.mtime [5] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01316_ ) );
OAI21_X1 _08989_ ( .A(\myclint.mtime [5] ), .B1(_01315_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01317_ ) );
AOI21_X1 _08990_ ( .A(fanout_net_1 ), .B1(_01316_ ), .B2(_01317_ ), .ZN(_00054_ ) );
OAI21_X1 _08991_ ( .A(_01265_ ), .B1(_01125_ ), .B2(\myclint.mtime [4] ), .ZN(_01318_ ) );
NOR2_X1 _08992_ ( .A1(_01318_ ), .A2(_01054_ ), .ZN(_00055_ ) );
INV_X1 _08993_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01319_ ) );
AND4_X1 _08994_ ( .A1(\myclint.mtime [57] ), .A2(_01112_ ), .A3(_01319_ ), .A4(_01088_ ), .ZN(_01320_ ) );
AND3_X1 _08995_ ( .A1(_01087_ ), .A2(_01319_ ), .A3(_01088_ ), .ZN(_01321_ ) );
OAI21_X1 _08996_ ( .A(_01242_ ), .B1(_01321_ ), .B2(\myclint.mtime [57] ), .ZN(_01322_ ) );
NOR2_X1 _08997_ ( .A1(_01320_ ), .A2(_01322_ ), .ZN(_00056_ ) );
AND2_X1 _08998_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01323_ ) );
INV_X1 _08999_ ( .A(_01323_ ), .ZN(_01324_ ) );
OR3_X1 _09000_ ( .A1(_01324_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01325_ ) );
OAI21_X1 _09001_ ( .A(\myclint.mtime [3] ), .B1(_01324_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01326_ ) );
AOI21_X1 _09002_ ( .A(fanout_net_1 ), .B1(_01325_ ), .B2(_01326_ ), .ZN(_00057_ ) );
AOI21_X1 _09003_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01327_ ) );
NOR3_X1 _09004_ ( .A1(_01053_ ), .A2(_01327_ ), .A3(fanout_net_1 ), .ZN(_00058_ ) );
NOR2_X1 _09005_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01328_ ) );
NOR3_X1 _09006_ ( .A1(_01323_ ), .A2(_01328_ ), .A3(fanout_net_1 ), .ZN(_00059_ ) );
CLKBUF_X2 _09007_ ( .A(_01147_ ), .Z(_01329_ ) );
AND2_X1 _09008_ ( .A1(_01329_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_00060_ ) );
XNOR2_X1 _09009_ ( .A(_01140_ ), .B(\myclint.mtime [56] ), .ZN(_01330_ ) );
NOR2_X1 _09010_ ( .A1(_01330_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
NAND2_X1 _09011_ ( .A1(_01085_ ), .A2(_01086_ ), .ZN(_01331_ ) );
NOR2_X1 _09012_ ( .A1(_01331_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01332_ ) );
OAI21_X1 _09013_ ( .A(_01191_ ), .B1(_01332_ ), .B2(\myclint.mtime [55] ), .ZN(_01333_ ) );
INV_X1 _09014_ ( .A(_01112_ ), .ZN(_01334_ ) );
NOR2_X1 _09015_ ( .A1(_01334_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01335_ ) );
AOI21_X1 _09016_ ( .A(_01333_ ), .B1(_01335_ ), .B2(\myclint.mtime [55] ), .ZN(_00062_ ) );
NAND3_X1 _09017_ ( .A1(_01138_ ), .A2(_01086_ ), .A3(_01151_ ), .ZN(_01336_ ) );
OR2_X1 _09018_ ( .A1(_01336_ ), .A2(\myclint.mtime [54] ), .ZN(_01337_ ) );
NAND2_X1 _09019_ ( .A1(_01336_ ), .A2(\myclint.mtime [54] ), .ZN(_01338_ ) );
AOI21_X1 _09020_ ( .A(fanout_net_2 ), .B1(_01337_ ), .B2(_01338_ ), .ZN(_00063_ ) );
MUX2_X1 _09021_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(fanout_net_38 ), .Z(_01339_ ) );
OR2_X1 _09022_ ( .A1(_01339_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01340_ ) );
INV_X16 _09023_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01341_ ) );
BUF_X4 _09024_ ( .A(_01341_ ), .Z(_01342_ ) );
MUX2_X1 _09025_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(fanout_net_38 ), .Z(_01343_ ) );
OAI21_X1 _09026_ ( .A(_01340_ ), .B1(_01342_ ), .B2(_01343_ ), .ZN(_01344_ ) );
INV_X1 _09027_ ( .A(\IF_ID_pc [27] ), .ZN(_01345_ ) );
MUX2_X1 _09028_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(fanout_net_38 ), .Z(_01346_ ) );
MUX2_X1 _09029_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(fanout_net_38 ), .Z(_01347_ ) );
MUX2_X2 _09030_ ( .A(_01346_ ), .B(_01347_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01348_ ) );
AOI22_X1 _09031_ ( .A1(_01344_ ), .A2(\IF_ID_pc [12] ), .B1(_01345_ ), .B2(_01348_ ), .ZN(_01349_ ) );
INV_X1 _09032_ ( .A(\IF_ID_pc [14] ), .ZN(_01350_ ) );
MUX2_X1 _09033_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(fanout_net_38 ), .Z(_01351_ ) );
MUX2_X1 _09034_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(fanout_net_38 ), .Z(_01352_ ) );
MUX2_X1 _09035_ ( .A(_01351_ ), .B(_01352_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01353_ ) );
INV_X32 _09036_ ( .A(fanout_net_38 ), .ZN(_01354_ ) );
BUF_X32 _09037_ ( .A(_01354_ ), .Z(_01355_ ) );
OR2_X1 _09038_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[1][23] ), .ZN(_01356_ ) );
OAI211_X1 _09039_ ( .A(_01356_ ), .B(_01341_ ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[0][23] ), .ZN(_01357_ ) );
OR2_X1 _09040_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[3][23] ), .ZN(_01358_ ) );
OAI211_X1 _09041_ ( .A(_01358_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[2][23] ), .ZN(_01359_ ) );
NAND2_X1 _09042_ ( .A1(_01357_ ), .A2(_01359_ ), .ZN(_01360_ ) );
INV_X1 _09043_ ( .A(_01360_ ), .ZN(_01361_ ) );
OAI221_X1 _09044_ ( .A(_01349_ ), .B1(_01350_ ), .B2(_01353_ ), .C1(\IF_ID_pc [28] ), .C2(_01361_ ), .ZN(_01362_ ) );
INV_X1 _09045_ ( .A(\IF_ID_pc [7] ), .ZN(_01363_ ) );
OR2_X4 _09046_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[1][2] ), .ZN(_01364_ ) );
OAI211_X2 _09047_ ( .A(_01364_ ), .B(_01341_ ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[0][2] ), .ZN(_01365_ ) );
OR2_X4 _09048_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[3][2] ), .ZN(_01366_ ) );
OAI211_X2 _09049_ ( .A(_01366_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[2][2] ), .ZN(_01367_ ) );
NAND2_X1 _09050_ ( .A1(_01365_ ), .A2(_01367_ ), .ZN(_01368_ ) );
AOI22_X1 _09051_ ( .A1(_01361_ ), .A2(\IF_ID_pc [28] ), .B1(_01363_ ), .B2(_01368_ ), .ZN(_01369_ ) );
INV_X1 _09052_ ( .A(\IF_ID_pc [20] ), .ZN(_01370_ ) );
MUX2_X1 _09053_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(fanout_net_38 ), .Z(_01371_ ) );
MUX2_X1 _09054_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(fanout_net_38 ), .Z(_01372_ ) );
MUX2_X1 _09055_ ( .A(_01371_ ), .B(_01372_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01373_ ) );
OAI221_X1 _09056_ ( .A(_01369_ ), .B1(_01370_ ), .B2(_01373_ ), .C1(_01363_ ), .C2(_01368_ ), .ZN(_01374_ ) );
MUX2_X1 _09057_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_38 ), .Z(_01375_ ) );
MUX2_X1 _09058_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_38 ), .Z(_01376_ ) );
MUX2_X2 _09059_ ( .A(_01375_ ), .B(_01376_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01377_ ) );
INV_X1 _09060_ ( .A(_01377_ ), .ZN(_01378_ ) );
INV_X1 _09061_ ( .A(\IF_ID_pc [24] ), .ZN(_01379_ ) );
OR2_X4 _09062_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[1][19] ), .ZN(_01380_ ) );
OAI211_X2 _09063_ ( .A(_01380_ ), .B(_01341_ ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[0][19] ), .ZN(_01381_ ) );
OR2_X1 _09064_ ( .A1(_01354_ ), .A2(\myifu.myicache.tag[3][19] ), .ZN(_01382_ ) );
OAI211_X1 _09065_ ( .A(_01382_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[2][19] ), .ZN(_01383_ ) );
NAND2_X1 _09066_ ( .A1(_01381_ ), .A2(_01383_ ), .ZN(_01384_ ) );
AOI22_X1 _09067_ ( .A1(_01378_ ), .A2(\IF_ID_pc [16] ), .B1(_01379_ ), .B2(_01384_ ), .ZN(_01385_ ) );
NAND2_X1 _09068_ ( .A1(_01373_ ), .A2(_01370_ ), .ZN(_01386_ ) );
OAI211_X2 _09069_ ( .A(_01385_ ), .B(_01386_ ), .C1(_01379_ ), .C2(_01384_ ), .ZN(_01387_ ) );
INV_X1 _09070_ ( .A(\IF_ID_pc [25] ), .ZN(_01388_ ) );
MUX2_X1 _09071_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(fanout_net_38 ), .Z(_01389_ ) );
MUX2_X1 _09072_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_38 ), .Z(_01390_ ) );
MUX2_X1 _09073_ ( .A(_01389_ ), .B(_01390_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01391_ ) );
MUX2_X1 _09074_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(fanout_net_38 ), .Z(_01392_ ) );
MUX2_X1 _09075_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(fanout_net_38 ), .Z(_01393_ ) );
MUX2_X2 _09076_ ( .A(_01392_ ), .B(_01393_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01394_ ) );
INV_X1 _09077_ ( .A(\IF_ID_pc [10] ), .ZN(_01395_ ) );
AOI22_X1 _09078_ ( .A1(_01388_ ), .A2(_01391_ ), .B1(_01394_ ), .B2(_01395_ ), .ZN(_01396_ ) );
MUX2_X1 _09079_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(fanout_net_38 ), .Z(_01397_ ) );
MUX2_X1 _09080_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(fanout_net_38 ), .Z(_01398_ ) );
MUX2_X2 _09081_ ( .A(_01397_ ), .B(_01398_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01399_ ) );
INV_X1 _09082_ ( .A(\IF_ID_pc [18] ), .ZN(_01400_ ) );
NAND2_X1 _09083_ ( .A1(_01399_ ), .A2(_01400_ ), .ZN(_01401_ ) );
INV_X1 _09084_ ( .A(\IF_ID_pc [23] ), .ZN(_01402_ ) );
OR2_X1 _09085_ ( .A1(_01354_ ), .A2(\myifu.myicache.tag[3][18] ), .ZN(_01403_ ) );
OAI211_X1 _09086_ ( .A(_01403_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[2][18] ), .ZN(_01404_ ) );
OR2_X1 _09087_ ( .A1(fanout_net_38 ), .A2(\myifu.myicache.tag[0][18] ), .ZN(_01405_ ) );
BUF_X2 _09088_ ( .A(_01354_ ), .Z(_01406_ ) );
OAI211_X1 _09089_ ( .A(_01405_ ), .B(_01341_ ), .C1(_01406_ ), .C2(\myifu.myicache.tag[1][18] ), .ZN(_01407_ ) );
NAND2_X1 _09090_ ( .A1(_01404_ ), .A2(_01407_ ), .ZN(_01408_ ) );
OAI211_X1 _09091_ ( .A(_01396_ ), .B(_01401_ ), .C1(_01402_ ), .C2(_01408_ ), .ZN(_01409_ ) );
NOR4_X2 _09092_ ( .A1(_01362_ ), .A2(_01374_ ), .A3(_01387_ ), .A4(_01409_ ), .ZN(_01410_ ) );
OR2_X1 _09093_ ( .A1(_01354_ ), .A2(\myifu.myicache.tag[1][3] ), .ZN(_01411_ ) );
OAI211_X1 _09094_ ( .A(_01411_ ), .B(_01341_ ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[0][3] ), .ZN(_01412_ ) );
OR2_X1 _09095_ ( .A1(fanout_net_38 ), .A2(\myifu.myicache.tag[2][3] ), .ZN(_01413_ ) );
OAI211_X1 _09096_ ( .A(_01413_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01406_ ), .C2(\myifu.myicache.tag[3][3] ), .ZN(_01414_ ) );
AOI21_X1 _09097_ ( .A(\IF_ID_pc [8] ), .B1(_01412_ ), .B2(_01414_ ), .ZN(_01415_ ) );
AOI21_X1 _09098_ ( .A(_01415_ ), .B1(_01350_ ), .B2(_01353_ ), .ZN(_01416_ ) );
MUX2_X1 _09099_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(fanout_net_38 ), .Z(_01417_ ) );
MUX2_X1 _09100_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(fanout_net_38 ), .Z(_01418_ ) );
MUX2_X1 _09101_ ( .A(_01417_ ), .B(_01418_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01419_ ) );
INV_X1 _09102_ ( .A(\IF_ID_pc [21] ), .ZN(_01420_ ) );
AOI22_X1 _09103_ ( .A1(_01419_ ), .A2(_01420_ ), .B1(_01408_ ), .B2(_01402_ ), .ZN(_01421_ ) );
NAND2_X1 _09104_ ( .A1(_01416_ ), .A2(_01421_ ), .ZN(_01422_ ) );
OAI22_X1 _09105_ ( .A1(_01378_ ), .A2(\IF_ID_pc [16] ), .B1(_01400_ ), .B2(_01399_ ), .ZN(_01423_ ) );
NOR2_X1 _09106_ ( .A1(_01419_ ), .A2(_01420_ ), .ZN(_01424_ ) );
AND3_X1 _09107_ ( .A1(_01412_ ), .A2(\IF_ID_pc [8] ), .A3(_01414_ ), .ZN(_01425_ ) );
NOR4_X1 _09108_ ( .A1(_01422_ ), .A2(_01423_ ), .A3(_01424_ ), .A4(_01425_ ), .ZN(_01426_ ) );
OR2_X1 _09109_ ( .A1(_01406_ ), .A2(\myifu.myicache.tag[3][0] ), .ZN(_01427_ ) );
OAI211_X1 _09110_ ( .A(_01427_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myifu.myicache.tag[2][0] ), .ZN(_01428_ ) );
INV_X1 _09111_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01429_ ) );
OR2_X1 _09112_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][0] ), .ZN(_01430_ ) );
OAI211_X1 _09113_ ( .A(_01430_ ), .B(_01342_ ), .C1(_01406_ ), .C2(\myifu.myicache.tag[1][0] ), .ZN(_01431_ ) );
AND3_X1 _09114_ ( .A1(_01428_ ), .A2(_01429_ ), .A3(_01431_ ), .ZN(_01432_ ) );
BUF_X32 _09115_ ( .A(_01354_ ), .Z(_01433_ ) );
OR2_X1 _09116_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[1][8] ), .ZN(_01434_ ) );
OAI211_X1 _09117_ ( .A(_01434_ ), .B(_01342_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][8] ), .ZN(_01435_ ) );
OR2_X1 _09118_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[3][8] ), .ZN(_01436_ ) );
OAI211_X1 _09119_ ( .A(_01436_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][8] ), .ZN(_01437_ ) );
AOI21_X1 _09120_ ( .A(\IF_ID_pc [13] ), .B1(_01435_ ), .B2(_01437_ ), .ZN(_01438_ ) );
AOI21_X1 _09121_ ( .A(_01429_ ), .B1(_01428_ ), .B2(_01431_ ), .ZN(_01439_ ) );
NOR3_X1 _09122_ ( .A1(_01432_ ), .A2(_01438_ ), .A3(_01439_ ), .ZN(_01440_ ) );
NOR2_X1 _09123_ ( .A1(_01348_ ), .A2(_01345_ ), .ZN(_01441_ ) );
OR2_X1 _09124_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[1][24] ), .ZN(_01442_ ) );
OAI211_X1 _09125_ ( .A(_01442_ ), .B(_01342_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][24] ), .ZN(_01443_ ) );
OR2_X1 _09126_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[3][24] ), .ZN(_01444_ ) );
OAI211_X1 _09127_ ( .A(_01444_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][24] ), .ZN(_01445_ ) );
AND3_X1 _09128_ ( .A1(_01443_ ), .A2(_01445_ ), .A3(\IF_ID_pc [29] ), .ZN(_01446_ ) );
AND3_X1 _09129_ ( .A1(_01435_ ), .A2(_01437_ ), .A3(\IF_ID_pc [13] ), .ZN(_01447_ ) );
AOI21_X1 _09130_ ( .A(\IF_ID_pc [29] ), .B1(_01443_ ), .B2(_01445_ ), .ZN(_01448_ ) );
NOR4_X1 _09131_ ( .A1(_01441_ ), .A2(_01446_ ), .A3(_01447_ ), .A4(_01448_ ), .ZN(_01449_ ) );
AND3_X2 _09132_ ( .A1(_01426_ ), .A2(_01440_ ), .A3(_01449_ ), .ZN(_01450_ ) );
AND2_X2 _09133_ ( .A1(_01410_ ), .A2(_01450_ ), .ZN(_01451_ ) );
OR2_X4 _09134_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[1][4] ), .ZN(_01452_ ) );
OAI211_X1 _09135_ ( .A(_01452_ ), .B(_01341_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][4] ), .ZN(_01453_ ) );
OR2_X1 _09136_ ( .A1(_01354_ ), .A2(\myifu.myicache.tag[3][4] ), .ZN(_01454_ ) );
OAI211_X1 _09137_ ( .A(_01454_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][4] ), .ZN(_01455_ ) );
NAND2_X1 _09138_ ( .A1(_01453_ ), .A2(_01455_ ), .ZN(_01456_ ) );
XNOR2_X1 _09139_ ( .A(_01456_ ), .B(\IF_ID_pc [9] ), .ZN(_01457_ ) );
MUX2_X1 _09140_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01458_ ) );
MUX2_X1 _09141_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01459_ ) );
MUX2_X1 _09142_ ( .A(_01458_ ), .B(_01459_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01460_ ) );
OR2_X4 _09143_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_01461_ ) );
OAI211_X4 _09144_ ( .A(_01461_ ), .B(_01342_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_01462_ ) );
OR2_X4 _09145_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[3][25] ), .ZN(_01463_ ) );
OAI211_X4 _09146_ ( .A(_01463_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][25] ), .ZN(_01464_ ) );
NAND3_X1 _09147_ ( .A1(_01462_ ), .A2(_01464_ ), .A3(\IF_ID_pc [30] ), .ZN(_01465_ ) );
AND3_X1 _09148_ ( .A1(_01457_ ), .A2(_01460_ ), .A3(_01465_ ), .ZN(_01466_ ) );
OR2_X1 _09149_ ( .A1(_01406_ ), .A2(\myifu.myicache.tag[1][21] ), .ZN(_01467_ ) );
OAI211_X1 _09150_ ( .A(_01467_ ), .B(_01342_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][21] ), .ZN(_01468_ ) );
OR2_X1 _09151_ ( .A1(_01406_ ), .A2(\myifu.myicache.tag[3][21] ), .ZN(_01469_ ) );
OAI211_X1 _09152_ ( .A(_01469_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][21] ), .ZN(_01470_ ) );
INV_X1 _09153_ ( .A(\IF_ID_pc [26] ), .ZN(_01471_ ) );
AND3_X1 _09154_ ( .A1(_01468_ ), .A2(_01470_ ), .A3(_01471_ ), .ZN(_01472_ ) );
AOI21_X1 _09155_ ( .A(_01471_ ), .B1(_01468_ ), .B2(_01470_ ), .ZN(_01473_ ) );
OR2_X1 _09156_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][17] ), .ZN(_01474_ ) );
OAI211_X1 _09157_ ( .A(_01474_ ), .B(_01342_ ), .C1(_01406_ ), .C2(\myifu.myicache.tag[1][17] ), .ZN(_01475_ ) );
OR2_X1 _09158_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][17] ), .ZN(_01476_ ) );
OAI211_X1 _09159_ ( .A(_01476_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01406_ ), .C2(\myifu.myicache.tag[3][17] ), .ZN(_01477_ ) );
INV_X1 _09160_ ( .A(\IF_ID_pc [22] ), .ZN(_01478_ ) );
AND3_X1 _09161_ ( .A1(_01475_ ), .A2(_01477_ ), .A3(_01478_ ), .ZN(_01479_ ) );
AOI21_X1 _09162_ ( .A(_01478_ ), .B1(_01475_ ), .B2(_01477_ ), .ZN(_01480_ ) );
OAI221_X1 _09163_ ( .A(_01466_ ), .B1(_01472_ ), .B2(_01473_ ), .C1(_01479_ ), .C2(_01480_ ), .ZN(_01481_ ) );
OR2_X4 _09164_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01482_ ) );
OAI211_X2 _09165_ ( .A(_01482_ ), .B(_01341_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01483_ ) );
OR2_X1 _09166_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][12] ), .ZN(_01484_ ) );
OAI211_X1 _09167_ ( .A(_01484_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01406_ ), .C2(\myifu.myicache.tag[3][12] ), .ZN(_01485_ ) );
NAND2_X1 _09168_ ( .A1(_01483_ ), .A2(_01485_ ), .ZN(_01486_ ) );
INV_X1 _09169_ ( .A(\IF_ID_pc [17] ), .ZN(_01487_ ) );
XNOR2_X1 _09170_ ( .A(_01486_ ), .B(_01487_ ), .ZN(_01488_ ) );
OR2_X4 _09171_ ( .A1(_01354_ ), .A2(\myifu.myicache.tag[3][26] ), .ZN(_01489_ ) );
OAI211_X2 _09172_ ( .A(_01489_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][26] ), .ZN(_01490_ ) );
INV_X1 _09173_ ( .A(\IF_ID_pc [31] ), .ZN(_01491_ ) );
OR2_X4 _09174_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][26] ), .ZN(_01492_ ) );
OAI211_X1 _09175_ ( .A(_01492_ ), .B(_01341_ ), .C1(_01433_ ), .C2(\myifu.myicache.tag[1][26] ), .ZN(_01493_ ) );
AND3_X2 _09176_ ( .A1(_01490_ ), .A2(_01491_ ), .A3(_01493_ ), .ZN(_01494_ ) );
AOI21_X1 _09177_ ( .A(_01491_ ), .B1(_01490_ ), .B2(_01493_ ), .ZN(_01495_ ) );
OR2_X4 _09178_ ( .A1(_01354_ ), .A2(\myifu.myicache.tag[3][1] ), .ZN(_01496_ ) );
OAI211_X2 _09179_ ( .A(_01496_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][1] ), .ZN(_01497_ ) );
INV_X1 _09180_ ( .A(\IF_ID_pc [6] ), .ZN(_01498_ ) );
OR2_X4 _09181_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_01499_ ) );
OAI211_X2 _09182_ ( .A(_01499_ ), .B(_01341_ ), .C1(_01433_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_01500_ ) );
AND3_X2 _09183_ ( .A1(_01497_ ), .A2(_01498_ ), .A3(_01500_ ), .ZN(_01501_ ) );
AOI21_X1 _09184_ ( .A(_01498_ ), .B1(_01497_ ), .B2(_01500_ ), .ZN(_01502_ ) );
OAI22_X1 _09185_ ( .A1(_01494_ ), .A2(_01495_ ), .B1(_01501_ ), .B2(_01502_ ), .ZN(_01503_ ) );
OR2_X4 _09186_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[1][10] ), .ZN(_01504_ ) );
OAI211_X1 _09187_ ( .A(_01504_ ), .B(_01342_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][10] ), .ZN(_01505_ ) );
OR2_X4 _09188_ ( .A1(_01355_ ), .A2(\myifu.myicache.tag[3][10] ), .ZN(_01506_ ) );
OAI211_X1 _09189_ ( .A(_01506_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][10] ), .ZN(_01507_ ) );
AND3_X1 _09190_ ( .A1(_01505_ ), .A2(_01507_ ), .A3(\IF_ID_pc [15] ), .ZN(_01508_ ) );
AOI21_X1 _09191_ ( .A(\IF_ID_pc [15] ), .B1(_01505_ ), .B2(_01507_ ), .ZN(_01509_ ) );
OR4_X2 _09192_ ( .A1(_01488_ ), .A2(_01503_ ), .A3(_01508_ ), .A4(_01509_ ), .ZN(_01510_ ) );
OR2_X1 _09193_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_01511_ ) );
OAI211_X1 _09194_ ( .A(_01511_ ), .B(_01342_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_01512_ ) );
OR2_X1 _09195_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[3][6] ), .ZN(_01513_ ) );
OAI211_X1 _09196_ ( .A(_01513_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][6] ), .ZN(_01514_ ) );
NAND2_X1 _09197_ ( .A1(_01512_ ), .A2(_01514_ ), .ZN(_01515_ ) );
XNOR2_X1 _09198_ ( .A(_01515_ ), .B(\IF_ID_pc [11] ), .ZN(_01516_ ) );
OAI221_X1 _09199_ ( .A(_01516_ ), .B1(\IF_ID_pc [12] ), .B2(_01344_ ), .C1(_01395_ ), .C2(_01394_ ), .ZN(_01517_ ) );
OR2_X4 _09200_ ( .A1(_01433_ ), .A2(\myifu.myicache.tag[3][14] ), .ZN(_01518_ ) );
OAI211_X2 _09201_ ( .A(_01518_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][14] ), .ZN(_01519_ ) );
OR2_X1 _09202_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][14] ), .ZN(_01520_ ) );
OAI211_X1 _09203_ ( .A(_01520_ ), .B(_01342_ ), .C1(_01406_ ), .C2(\myifu.myicache.tag[1][14] ), .ZN(_01521_ ) );
AND3_X1 _09204_ ( .A1(_01519_ ), .A2(\IF_ID_pc [19] ), .A3(_01521_ ), .ZN(_01522_ ) );
NOR2_X1 _09205_ ( .A1(_01391_ ), .A2(_01388_ ), .ZN(_01523_ ) );
AOI21_X1 _09206_ ( .A(\IF_ID_pc [19] ), .B1(_01519_ ), .B2(_01521_ ), .ZN(_01524_ ) );
AOI21_X2 _09207_ ( .A(\IF_ID_pc [30] ), .B1(_01462_ ), .B2(_01464_ ), .ZN(_01525_ ) );
OR4_X4 _09208_ ( .A1(_01522_ ), .A2(_01523_ ), .A3(_01524_ ), .A4(_01525_ ), .ZN(_01526_ ) );
NOR4_X4 _09209_ ( .A1(_01481_ ), .A2(_01510_ ), .A3(_01517_ ), .A4(_01526_ ), .ZN(_01527_ ) );
NAND2_X2 _09210_ ( .A1(_01451_ ), .A2(_01527_ ), .ZN(_01528_ ) );
AND2_X4 _09211_ ( .A1(_01528_ ), .A2(\myifu.state [0] ), .ZN(_01529_ ) );
INV_X1 _09212_ ( .A(\myifu.wen_$_SDFFE_PP0P__Q_D ), .ZN(_01530_ ) );
NOR2_X4 _09213_ ( .A1(_01529_ ), .A2(_01530_ ), .ZN(_01531_ ) );
NOR2_X1 _09214_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01532_ ) );
NOR2_X4 _09215_ ( .A1(_01531_ ), .A2(_01532_ ), .ZN(_01533_ ) );
NAND4_X1 _09216_ ( .A1(\mylsu.state [0] ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_01534_ ) );
INV_X1 _09217_ ( .A(EXU_valid_LSU ), .ZN(_01535_ ) );
NOR2_X1 _09218_ ( .A1(_01534_ ), .A2(_01535_ ), .ZN(_01536_ ) );
INV_X1 _09219_ ( .A(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__B_A_$_ANDNOT__Y_A ), .ZN(_01537_ ) );
NOR2_X1 _09220_ ( .A1(_01536_ ), .A2(_01537_ ), .ZN(_01538_ ) );
NOR2_X4 _09221_ ( .A1(_01533_ ), .A2(_01538_ ), .ZN(_01539_ ) );
BUF_X8 _09222_ ( .A(_01539_ ), .Z(_01540_ ) );
CLKBUF_X2 _09223_ ( .A(_01534_ ), .Z(_01541_ ) );
CLKBUF_X2 _09224_ ( .A(_01541_ ), .Z(_01542_ ) );
CLKBUF_X2 _09225_ ( .A(_01535_ ), .Z(_01543_ ) );
OR3_X1 _09226_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(_01543_ ), .ZN(_01544_ ) );
BUF_X4 _09227_ ( .A(_01536_ ), .Z(_01545_ ) );
BUF_X4 _09228_ ( .A(_01545_ ), .Z(_01546_ ) );
OAI211_X1 _09229_ ( .A(_01540_ ), .B(_01544_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01546_ ), .ZN(_01547_ ) );
BUF_X4 _09230_ ( .A(_01529_ ), .Z(_01548_ ) );
BUF_X4 _09231_ ( .A(_01530_ ), .Z(_01549_ ) );
OAI221_X1 _09232_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_01550_ ) );
AND2_X1 _09233_ ( .A1(_01547_ ), .A2(_01550_ ), .ZN(_01551_ ) );
BUF_X8 _09234_ ( .A(_01539_ ), .Z(_01552_ ) );
CLKBUF_X2 _09235_ ( .A(_01535_ ), .Z(_01553_ ) );
OR3_X1 _09236_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(_01553_ ), .ZN(_01554_ ) );
OAI211_X1 _09237_ ( .A(_01552_ ), .B(_01554_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01545_ ), .ZN(_01555_ ) );
BUF_X8 _09238_ ( .A(_01529_ ), .Z(_01556_ ) );
BUF_X4 _09239_ ( .A(_01530_ ), .Z(_01557_ ) );
OAI221_X1 _09240_ ( .A(\IF_ID_pc [24] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01558_ ) );
AND2_X1 _09241_ ( .A1(_01555_ ), .A2(_01558_ ), .ZN(_01559_ ) );
OR3_X1 _09242_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(_01553_ ), .ZN(_01560_ ) );
OAI211_X1 _09243_ ( .A(_01552_ ), .B(_01560_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01545_ ), .ZN(_01561_ ) );
OAI221_X1 _09244_ ( .A(\IF_ID_pc [28] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01562_ ) );
AND2_X2 _09245_ ( .A1(_01561_ ), .A2(_01562_ ), .ZN(_01563_ ) );
OR3_X1 _09246_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(_01535_ ), .ZN(_01564_ ) );
OAI211_X1 _09247_ ( .A(_01539_ ), .B(_01564_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01545_ ), .ZN(_01565_ ) );
OAI221_X1 _09248_ ( .A(\IF_ID_pc [26] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01566_ ) );
AND2_X1 _09249_ ( .A1(_01565_ ), .A2(_01566_ ), .ZN(_01567_ ) );
NAND4_X1 _09250_ ( .A1(_01551_ ), .A2(_01559_ ), .A3(_01563_ ), .A4(_01567_ ), .ZN(_01568_ ) );
OR3_X1 _09251_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(_01553_ ), .ZN(_01569_ ) );
OAI211_X1 _09252_ ( .A(_01540_ ), .B(_01569_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01546_ ), .ZN(_01570_ ) );
OAI221_X1 _09253_ ( .A(\IF_ID_pc [22] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_01571_ ) );
AND2_X1 _09254_ ( .A1(_01570_ ), .A2(_01571_ ), .ZN(_01572_ ) );
OR3_X1 _09255_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(_01553_ ), .ZN(_01573_ ) );
OAI211_X1 _09256_ ( .A(_01552_ ), .B(_01573_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01545_ ), .ZN(_01574_ ) );
OAI221_X1 _09257_ ( .A(\IF_ID_pc [16] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01575_ ) );
AND2_X1 _09258_ ( .A1(_01574_ ), .A2(_01575_ ), .ZN(_01576_ ) );
OR3_X1 _09259_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(_01553_ ), .ZN(_01577_ ) );
OAI211_X1 _09260_ ( .A(_01552_ ), .B(_01577_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01546_ ), .ZN(_01578_ ) );
OAI221_X1 _09261_ ( .A(\IF_ID_pc [21] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01579_ ) );
AND2_X1 _09262_ ( .A1(_01578_ ), .A2(_01579_ ), .ZN(_01580_ ) );
OR3_X1 _09263_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(_01535_ ), .ZN(_01581_ ) );
OAI211_X1 _09264_ ( .A(_01552_ ), .B(_01581_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01545_ ), .ZN(_01582_ ) );
OAI221_X1 _09265_ ( .A(\IF_ID_pc [19] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01583_ ) );
AND2_X1 _09266_ ( .A1(_01582_ ), .A2(_01583_ ), .ZN(_01584_ ) );
NAND4_X1 _09267_ ( .A1(_01572_ ), .A2(_01576_ ), .A3(_01580_ ), .A4(_01584_ ), .ZN(_01585_ ) );
NOR2_X1 _09268_ ( .A1(_01568_ ), .A2(_01585_ ), .ZN(_01586_ ) );
OR3_X1 _09269_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(_01543_ ), .ZN(_01587_ ) );
OAI211_X1 _09270_ ( .A(_01540_ ), .B(_01587_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01546_ ), .ZN(_01588_ ) );
OAI221_X1 _09271_ ( .A(\IF_ID_pc [23] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_01589_ ) );
AND2_X1 _09272_ ( .A1(_01588_ ), .A2(_01589_ ), .ZN(_01590_ ) );
OR3_X1 _09273_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(_01553_ ), .ZN(_01591_ ) );
OAI211_X1 _09274_ ( .A(_01552_ ), .B(_01591_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01546_ ), .ZN(_01592_ ) );
OAI221_X1 _09275_ ( .A(\IF_ID_pc [17] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_01593_ ) );
AND2_X2 _09276_ ( .A1(_01592_ ), .A2(_01593_ ), .ZN(_01594_ ) );
OR3_X1 _09277_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(_01553_ ), .ZN(_01595_ ) );
OAI211_X1 _09278_ ( .A(_01552_ ), .B(_01595_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01545_ ), .ZN(_01596_ ) );
OAI221_X1 _09279_ ( .A(\IF_ID_pc [20] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01597_ ) );
AND2_X2 _09280_ ( .A1(_01596_ ), .A2(_01597_ ), .ZN(_01598_ ) );
OR3_X1 _09281_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(_01535_ ), .ZN(_01599_ ) );
OAI211_X1 _09282_ ( .A(_01539_ ), .B(_01599_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01545_ ), .ZN(_01600_ ) );
OAI221_X1 _09283_ ( .A(\IF_ID_pc [18] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01601_ ) );
AND2_X1 _09284_ ( .A1(_01600_ ), .A2(_01601_ ), .ZN(_01602_ ) );
NAND4_X1 _09285_ ( .A1(_01590_ ), .A2(_01594_ ), .A3(_01598_ ), .A4(_01602_ ), .ZN(_01603_ ) );
OR3_X1 _09286_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(_01553_ ), .ZN(_01604_ ) );
OAI211_X1 _09287_ ( .A(_01552_ ), .B(_01604_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01546_ ), .ZN(_01605_ ) );
OAI221_X1 _09288_ ( .A(\IF_ID_pc [30] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_01606_ ) );
AND2_X1 _09289_ ( .A1(_01605_ ), .A2(_01606_ ), .ZN(_01607_ ) );
OR3_X1 _09290_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(_01553_ ), .ZN(_01608_ ) );
OAI211_X1 _09291_ ( .A(_01552_ ), .B(_01608_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01545_ ), .ZN(_01609_ ) );
OAI221_X1 _09292_ ( .A(\IF_ID_pc [29] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01610_ ) );
AND2_X1 _09293_ ( .A1(_01609_ ), .A2(_01610_ ), .ZN(_01611_ ) );
OR3_X1 _09294_ ( .A1(_01541_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(_01553_ ), .ZN(_01612_ ) );
OAI211_X1 _09295_ ( .A(_01552_ ), .B(_01612_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01545_ ), .ZN(_01613_ ) );
OAI221_X1 _09296_ ( .A(\IF_ID_pc [27] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01556_ ), .C2(_01557_ ), .ZN(_01614_ ) );
AND2_X1 _09297_ ( .A1(_01613_ ), .A2(_01614_ ), .ZN(_01615_ ) );
OR3_X1 _09298_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [25] ), .A3(_01543_ ), .ZN(_01616_ ) );
OAI211_X2 _09299_ ( .A(_01540_ ), .B(_01616_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_01546_ ), .ZN(_01617_ ) );
INV_X1 _09300_ ( .A(_01533_ ), .ZN(_01618_ ) );
OAI21_X2 _09301_ ( .A(_01617_ ), .B1(_01388_ ), .B2(_01618_ ), .ZN(\io_master_araddr [25] ) );
NAND4_X1 _09302_ ( .A1(_01607_ ), .A2(_01611_ ), .A3(_01615_ ), .A4(\io_master_araddr [25] ), .ZN(_01619_ ) );
NOR2_X1 _09303_ ( .A1(_01603_ ), .A2(_01619_ ), .ZN(_01620_ ) );
NAND3_X1 _09304_ ( .A1(_01586_ ), .A2(_01620_ ), .A3(\myclint.rvalid ), .ZN(_01621_ ) );
BUF_X2 _09305_ ( .A(_01540_ ), .Z(_01622_ ) );
CLKBUF_X2 _09306_ ( .A(_01622_ ), .Z(_01623_ ) );
BUF_X2 _09307_ ( .A(_01623_ ), .Z(\io_master_arid [1] ) );
NOR2_X1 _09308_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_01624_ ) );
AND3_X1 _09309_ ( .A1(_01528_ ), .A2(\myifu.state [0] ), .A3(_01624_ ), .ZN(_01625_ ) );
INV_X1 _09310_ ( .A(_01625_ ), .ZN(_01626_ ) );
AOI21_X1 _09311_ ( .A(_01532_ ), .B1(_01626_ ), .B2(\myifu.wen_$_SDFFE_PP0P__Q_D ), .ZN(_01627_ ) );
NOR2_X1 _09312_ ( .A1(\io_master_arid [1] ), .A2(_01627_ ), .ZN(_01628_ ) );
NOR2_X1 _09313_ ( .A1(_01621_ ), .A2(_01628_ ), .ZN(_01629_ ) );
INV_X1 _09314_ ( .A(\myclint.rvalid ), .ZN(_01630_ ) );
INV_X1 _09315_ ( .A(_01546_ ), .ZN(_01631_ ) );
OAI21_X1 _09316_ ( .A(_01631_ ), .B1(_01531_ ), .B2(_01532_ ), .ZN(_01632_ ) );
NAND2_X1 _09317_ ( .A1(_01051_ ), .A2(\myifu.state [0] ), .ZN(_01633_ ) );
NOR2_X1 _09318_ ( .A1(_01633_ ), .A2(\myidu.stall_quest_fencei ), .ZN(_01634_ ) );
OR3_X1 _09319_ ( .A1(_01531_ ), .A2(_01532_ ), .A3(_01634_ ), .ZN(_01635_ ) );
NAND4_X1 _09320_ ( .A1(_01586_ ), .A2(_01620_ ), .A3(_01632_ ), .A4(_01635_ ), .ZN(_01636_ ) );
AOI211_X1 _09321_ ( .A(fanout_net_2 ), .B(_01629_ ), .C1(_01630_ ), .C2(_01636_ ), .ZN(_00064_ ) );
INV_X1 _09322_ ( .A(\LS_WB_wen_csreg [1] ), .ZN(_01637_ ) );
CLKBUF_X2 _09323_ ( .A(_01637_ ), .Z(_01638_ ) );
AND2_X1 _09324_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00065_ ) );
AND2_X1 _09325_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [4] ), .ZN(_00066_ ) );
AND2_X1 _09326_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00067_ ) );
AND2_X1 _09327_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00068_ ) );
AND2_X1 _09328_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00069_ ) );
AND2_X1 _09329_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00070_ ) );
AND2_X1 _09330_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [20] ), .ZN(_00071_ ) );
AND2_X1 _09331_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [19] ), .ZN(_00072_ ) );
AND2_X1 _09332_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [18] ), .ZN(_00073_ ) );
AND2_X1 _09333_ ( .A1(_01638_ ), .A2(\LS_WB_wdata_csreg [17] ), .ZN(_00074_ ) );
CLKBUF_X2 _09334_ ( .A(_01637_ ), .Z(_01639_ ) );
AND2_X1 _09335_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00075_ ) );
AND2_X1 _09336_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00076_ ) );
AND2_X1 _09337_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [2] ), .ZN(_00077_ ) );
AND2_X1 _09338_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00078_ ) );
AND2_X1 _09339_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00079_ ) );
AND2_X1 _09340_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00080_ ) );
AND2_X1 _09341_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00081_ ) );
AND2_X1 _09342_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00082_ ) );
AND2_X1 _09343_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00083_ ) );
AND2_X1 _09344_ ( .A1(_01639_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00084_ ) );
CLKBUF_X2 _09345_ ( .A(_01637_ ), .Z(_01640_ ) );
AND2_X1 _09346_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00085_ ) );
AND2_X1 _09347_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [6] ), .ZN(_00086_ ) );
AND2_X1 _09348_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00087_ ) );
AND2_X1 _09349_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00088_ ) );
AND2_X1 _09350_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00089_ ) );
AND2_X1 _09351_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00090_ ) );
AND2_X1 _09352_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00091_ ) );
AND2_X1 _09353_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00092_ ) );
AND2_X1 _09354_ ( .A1(_01640_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00093_ ) );
INV_X1 _09355_ ( .A(check_quest ), .ZN(_01641_ ) );
NOR2_X1 _09356_ ( .A1(_01641_ ), .A2(check_assert ), .ZN(_01642_ ) );
INV_X1 _09357_ ( .A(IDU_valid_EXU ), .ZN(_01643_ ) );
NOR2_X1 _09358_ ( .A1(_01643_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
OAI21_X1 _09359_ ( .A(_01191_ ), .B1(_01642_ ), .B2(\myexu.state_$_ANDNOT__B_Y ), .ZN(_01644_ ) );
INV_X1 _09360_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_01645_ ) );
AND2_X1 _09361_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_01646_ ) );
INV_X1 _09362_ ( .A(\ID_EX_typ [5] ), .ZN(_01647_ ) );
NOR2_X1 _09363_ ( .A1(_01647_ ), .A2(\ID_EX_typ [6] ), .ZN(_01648_ ) );
AND2_X2 _09364_ ( .A1(_01648_ ), .A2(\ID_EX_typ [7] ), .ZN(_01649_ ) );
CLKBUF_X2 _09365_ ( .A(_01649_ ), .Z(_01650_ ) );
AOI221_X4 _09366_ ( .A(_01645_ ), .B1(\ID_EX_typ [7] ), .B2(_01646_ ), .C1(_01650_ ), .C2(fanout_net_8 ), .ZN(_01651_ ) );
INV_X1 _09367_ ( .A(_01649_ ), .ZN(_01652_ ) );
BUF_X4 _09368_ ( .A(_01652_ ), .Z(_01653_ ) );
BUF_X4 _09369_ ( .A(_01653_ ), .Z(_01654_ ) );
BUF_X4 _09370_ ( .A(_01654_ ), .Z(_01655_ ) );
INV_X1 _09371_ ( .A(\ID_EX_typ [7] ), .ZN(_01656_ ) );
NOR2_X1 _09372_ ( .A1(_01656_ ), .A2(\ID_EX_typ [6] ), .ZN(_01657_ ) );
AOI211_X1 _09373_ ( .A(_01641_ ), .B(check_assert ), .C1(_01657_ ), .C2(_01647_ ), .ZN(_01658_ ) );
INV_X1 _09374_ ( .A(\ID_EX_typ [6] ), .ZN(_01659_ ) );
AND4_X1 _09375_ ( .A1(\ID_EX_typ [7] ), .A2(_01659_ ), .A3(_01647_ ), .A4(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_01660_ ) );
OAI21_X1 _09376_ ( .A(_01655_ ), .B1(_01658_ ), .B2(_01660_ ), .ZN(_01661_ ) );
AOI21_X1 _09377_ ( .A(_01644_ ), .B1(_01651_ ), .B2(_01661_ ), .ZN(_00094_ ) );
INV_X32 _09378_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_01662_ ) );
OAI21_X4 _09379_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_01662_ ), .B2(\ID_EX_rs1 [1] ), .ZN(_01663_ ) );
NOR2_X1 _09380_ ( .A1(\EX_LS_dest_reg [4] ), .A2(\EX_LS_dest_reg [3] ), .ZN(_01664_ ) );
NOR3_X4 _09381_ ( .A1(\EX_LS_dest_reg [2] ), .A2(\EX_LS_dest_reg [1] ), .A3(\EX_LS_dest_reg [0] ), .ZN(_01665_ ) );
AOI221_X2 _09382_ ( .A(_01663_ ), .B1(\ID_EX_rs1 [1] ), .B2(_01662_ ), .C1(_01664_ ), .C2(_01665_ ), .ZN(_01666_ ) );
XNOR2_X1 _09383_ ( .A(\ID_EX_rs1 [3] ), .B(\EX_LS_dest_reg [3] ), .ZN(_01667_ ) );
XNOR2_X1 _09384_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .ZN(_01668_ ) );
XNOR2_X1 _09385_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .ZN(_01669_ ) );
XNOR2_X2 _09386_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_01670_ ) );
AND4_X2 _09387_ ( .A1(_01667_ ), .A2(_01668_ ), .A3(_01669_ ), .A4(_01670_ ), .ZN(_01671_ ) );
NAND2_X4 _09388_ ( .A1(_01666_ ), .A2(_01671_ ), .ZN(_01672_ ) );
INV_X32 _09389_ ( .A(\EX_LS_flag [0] ), .ZN(_01673_ ) );
NAND2_X4 _09390_ ( .A1(_01673_ ), .A2(\EX_LS_flag [1] ), .ZN(_01674_ ) );
INV_X8 _09391_ ( .A(\EX_LS_flag [2] ), .ZN(_01675_ ) );
NOR2_X4 _09392_ ( .A1(_01674_ ), .A2(_01675_ ), .ZN(_01676_ ) );
INV_X4 _09393_ ( .A(_01676_ ), .ZN(_01677_ ) );
NOR2_X2 _09394_ ( .A1(_01673_ ), .A2(\EX_LS_flag [1] ), .ZN(_01678_ ) );
INV_X1 _09395_ ( .A(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_01679_ ) );
AOI22_X2 _09396_ ( .A1(_01678_ ), .A2(_01679_ ), .B1(_01675_ ), .B2(\EX_LS_flag [0] ), .ZN(_01680_ ) );
AND2_X4 _09397_ ( .A1(_01677_ ), .A2(_01680_ ), .ZN(_01681_ ) );
NOR2_X1 _09398_ ( .A1(_01672_ ), .A2(_01681_ ), .ZN(_01682_ ) );
INV_X2 _09399_ ( .A(_01682_ ), .ZN(_01683_ ) );
INV_X32 _09400_ ( .A(fanout_net_12 ), .ZN(_01684_ ) );
BUF_X32 _09401_ ( .A(_01684_ ), .Z(_01685_ ) );
BUF_X8 _09402_ ( .A(_01685_ ), .Z(_01686_ ) );
BUF_X4 _09403_ ( .A(_01686_ ), .Z(_01687_ ) );
BUF_X2 _09404_ ( .A(_01687_ ), .Z(_01688_ ) );
BUF_X2 _09405_ ( .A(_01688_ ), .Z(_01689_ ) );
NOR2_X1 _09406_ ( .A1(_01689_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01690_ ) );
OAI21_X1 _09407_ ( .A(fanout_net_20 ), .B1(fanout_net_12 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01691_ ) );
NOR2_X1 _09408_ ( .A1(fanout_net_12 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01692_ ) );
INV_X1 _09409_ ( .A(fanout_net_20 ), .ZN(_01693_ ) );
BUF_X4 _09410_ ( .A(_01693_ ), .Z(_01694_ ) );
BUF_X4 _09411_ ( .A(_01694_ ), .Z(_01695_ ) );
BUF_X4 _09412_ ( .A(_01695_ ), .Z(_01696_ ) );
BUF_X4 _09413_ ( .A(_01696_ ), .Z(_01697_ ) );
BUF_X8 _09414_ ( .A(_01686_ ), .Z(_01698_ ) );
BUF_X2 _09415_ ( .A(_01698_ ), .Z(_01699_ ) );
BUF_X8 _09416_ ( .A(_01699_ ), .Z(_01700_ ) );
OAI21_X1 _09417_ ( .A(_01697_ ), .B1(_01700_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01701_ ) );
OAI221_X1 _09418_ ( .A(fanout_net_23 ), .B1(_01690_ ), .B2(_01691_ ), .C1(_01692_ ), .C2(_01701_ ), .ZN(_01702_ ) );
MUX2_X1 _09419_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01703_ ) );
MUX2_X1 _09420_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01704_ ) );
MUX2_X1 _09421_ ( .A(_01703_ ), .B(_01704_ ), .S(_01697_ ), .Z(_01705_ ) );
OAI211_X1 _09422_ ( .A(fanout_net_24 ), .B(_01702_ ), .C1(_01705_ ), .C2(fanout_net_23 ), .ZN(_01706_ ) );
MUX2_X1 _09423_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01707_ ) );
AND2_X1 _09424_ ( .A1(_01707_ ), .A2(_01697_ ), .ZN(_01708_ ) );
MUX2_X1 _09425_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01709_ ) );
AOI211_X1 _09426_ ( .A(fanout_net_23 ), .B(_01708_ ), .C1(fanout_net_20 ), .C2(_01709_ ), .ZN(_01710_ ) );
INV_X1 _09427_ ( .A(fanout_net_24 ), .ZN(_01711_ ) );
BUF_X4 _09428_ ( .A(_01711_ ), .Z(_01712_ ) );
BUF_X4 _09429_ ( .A(_01712_ ), .Z(_01713_ ) );
BUF_X4 _09430_ ( .A(_01713_ ), .Z(_01714_ ) );
MUX2_X1 _09431_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01715_ ) );
MUX2_X1 _09432_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01716_ ) );
MUX2_X1 _09433_ ( .A(_01715_ ), .B(_01716_ ), .S(fanout_net_20 ), .Z(_01717_ ) );
INV_X1 _09434_ ( .A(fanout_net_23 ), .ZN(_01718_ ) );
BUF_X4 _09435_ ( .A(_01718_ ), .Z(_01719_ ) );
BUF_X4 _09436_ ( .A(_01719_ ), .Z(_01720_ ) );
BUF_X4 _09437_ ( .A(_01720_ ), .Z(_01721_ ) );
BUF_X4 _09438_ ( .A(_01721_ ), .Z(_01722_ ) );
OAI21_X1 _09439_ ( .A(_01714_ ), .B1(_01717_ ), .B2(_01722_ ), .ZN(_01723_ ) );
OAI211_X2 _09440_ ( .A(_01683_ ), .B(_01706_ ), .C1(_01710_ ), .C2(_01723_ ), .ZN(_01724_ ) );
BUF_X8 _09441_ ( .A(_01672_ ), .Z(_01725_ ) );
BUF_X16 _09442_ ( .A(_01725_ ), .Z(_01726_ ) );
BUF_X16 _09443_ ( .A(_01726_ ), .Z(_01727_ ) );
BUF_X8 _09444_ ( .A(_01681_ ), .Z(_01728_ ) );
BUF_X16 _09445_ ( .A(_01728_ ), .Z(_01729_ ) );
BUF_X2 _09446_ ( .A(_01729_ ), .Z(_01730_ ) );
OR3_X1 _09447_ ( .A1(_01727_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_01730_ ), .ZN(_01731_ ) );
AND2_X2 _09448_ ( .A1(_01724_ ), .A2(_01731_ ), .ZN(_01732_ ) );
INV_X1 _09449_ ( .A(\ID_EX_imm [30] ), .ZN(_01733_ ) );
XNOR2_X1 _09450_ ( .A(_01732_ ), .B(_01733_ ), .ZN(_01734_ ) );
OR2_X1 _09451_ ( .A1(_01689_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01735_ ) );
BUF_X4 _09452_ ( .A(_01694_ ), .Z(_01736_ ) );
BUF_X4 _09453_ ( .A(_01736_ ), .Z(_01737_ ) );
BUF_X4 _09454_ ( .A(_01737_ ), .Z(_01738_ ) );
BUF_X4 _09455_ ( .A(_01738_ ), .Z(_01739_ ) );
OAI211_X1 _09456_ ( .A(_01735_ ), .B(_01739_ ), .C1(fanout_net_12 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01740_ ) );
OR2_X1 _09457_ ( .A1(_01689_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01741_ ) );
OAI211_X1 _09458_ ( .A(_01741_ ), .B(fanout_net_20 ), .C1(fanout_net_12 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01742_ ) );
NAND3_X1 _09459_ ( .A1(_01740_ ), .A2(_01742_ ), .A3(_01722_ ), .ZN(_01743_ ) );
MUX2_X1 _09460_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01744_ ) );
MUX2_X1 _09461_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01745_ ) );
MUX2_X1 _09462_ ( .A(_01744_ ), .B(_01745_ ), .S(_01739_ ), .Z(_01746_ ) );
BUF_X4 _09463_ ( .A(_01721_ ), .Z(_01747_ ) );
OAI211_X1 _09464_ ( .A(fanout_net_24 ), .B(_01743_ ), .C1(_01746_ ), .C2(_01747_ ), .ZN(_01748_ ) );
OR2_X1 _09465_ ( .A1(_01689_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01749_ ) );
OAI211_X1 _09466_ ( .A(_01749_ ), .B(fanout_net_20 ), .C1(fanout_net_12 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01750_ ) );
OR2_X1 _09467_ ( .A1(fanout_net_12 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01751_ ) );
OAI211_X1 _09468_ ( .A(_01751_ ), .B(_01739_ ), .C1(_01700_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01752_ ) );
NAND3_X1 _09469_ ( .A1(_01750_ ), .A2(_01722_ ), .A3(_01752_ ), .ZN(_01753_ ) );
MUX2_X1 _09470_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01754_ ) );
MUX2_X1 _09471_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01755_ ) );
MUX2_X1 _09472_ ( .A(_01754_ ), .B(_01755_ ), .S(_01739_ ), .Z(_01756_ ) );
OAI211_X1 _09473_ ( .A(_01714_ ), .B(_01753_ ), .C1(_01756_ ), .C2(_01747_ ), .ZN(_01757_ ) );
BUF_X4 _09474_ ( .A(_01728_ ), .Z(_01758_ ) );
BUF_X4 _09475_ ( .A(_01758_ ), .Z(_01759_ ) );
BUF_X2 _09476_ ( .A(_01759_ ), .Z(_01760_ ) );
BUF_X4 _09477_ ( .A(_01725_ ), .Z(_01761_ ) );
BUF_X2 _09478_ ( .A(_01761_ ), .Z(_01762_ ) );
OAI211_X1 _09479_ ( .A(_01748_ ), .B(_01757_ ), .C1(_01760_ ), .C2(_01762_ ), .ZN(_01763_ ) );
OR3_X1 _09480_ ( .A1(_01762_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_01760_ ), .ZN(_01764_ ) );
NAND2_X4 _09481_ ( .A1(_01763_ ), .A2(_01764_ ), .ZN(_01765_ ) );
XNOR2_X1 _09482_ ( .A(_01765_ ), .B(\ID_EX_imm [28] ), .ZN(_01766_ ) );
CLKBUF_X2 _09483_ ( .A(_01686_ ), .Z(_01767_ ) );
OR2_X1 _09484_ ( .A1(_01767_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01768_ ) );
OAI211_X1 _09485_ ( .A(_01768_ ), .B(_01696_ ), .C1(fanout_net_12 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01769_ ) );
BUF_X4 _09486_ ( .A(_01719_ ), .Z(_01770_ ) );
BUF_X4 _09487_ ( .A(_01770_ ), .Z(_01771_ ) );
OR2_X1 _09488_ ( .A1(fanout_net_12 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01772_ ) );
OAI211_X1 _09489_ ( .A(_01772_ ), .B(fanout_net_20 ), .C1(_01699_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01773_ ) );
NAND3_X1 _09490_ ( .A1(_01769_ ), .A2(_01771_ ), .A3(_01773_ ), .ZN(_01774_ ) );
MUX2_X1 _09491_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01775_ ) );
MUX2_X1 _09492_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01776_ ) );
BUF_X4 _09493_ ( .A(_01695_ ), .Z(_01777_ ) );
MUX2_X1 _09494_ ( .A(_01775_ ), .B(_01776_ ), .S(_01777_ ), .Z(_01778_ ) );
BUF_X4 _09495_ ( .A(_01720_ ), .Z(_01779_ ) );
OAI211_X1 _09496_ ( .A(_01713_ ), .B(_01774_ ), .C1(_01778_ ), .C2(_01779_ ), .ZN(_01780_ ) );
OR2_X1 _09497_ ( .A1(_01767_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01781_ ) );
OAI211_X1 _09498_ ( .A(_01781_ ), .B(_01696_ ), .C1(fanout_net_12 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01782_ ) );
OR2_X1 _09499_ ( .A1(fanout_net_12 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01783_ ) );
OAI211_X1 _09500_ ( .A(_01783_ ), .B(fanout_net_20 ), .C1(_01699_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01784_ ) );
NAND3_X1 _09501_ ( .A1(_01782_ ), .A2(fanout_net_23 ), .A3(_01784_ ), .ZN(_01785_ ) );
MUX2_X1 _09502_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01786_ ) );
MUX2_X1 _09503_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01787_ ) );
MUX2_X1 _09504_ ( .A(_01786_ ), .B(_01787_ ), .S(fanout_net_20 ), .Z(_01788_ ) );
OAI211_X1 _09505_ ( .A(fanout_net_24 ), .B(_01785_ ), .C1(_01788_ ), .C2(fanout_net_23 ), .ZN(_01789_ ) );
BUF_X16 _09506_ ( .A(_01726_ ), .Z(_01790_ ) );
OAI211_X4 _09507_ ( .A(_01780_ ), .B(_01789_ ), .C1(_01759_ ), .C2(_01790_ ), .ZN(_01791_ ) );
OR3_X2 _09508_ ( .A1(_01761_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01758_ ), .ZN(_01792_ ) );
NAND2_X4 _09509_ ( .A1(_01791_ ), .A2(_01792_ ), .ZN(_01793_ ) );
INV_X1 _09510_ ( .A(\ID_EX_imm [22] ), .ZN(_01794_ ) );
XNOR2_X1 _09511_ ( .A(_01793_ ), .B(_01794_ ), .ZN(_01795_ ) );
OR2_X1 _09512_ ( .A1(_01698_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01796_ ) );
OAI211_X1 _09513_ ( .A(_01796_ ), .B(_01777_ ), .C1(fanout_net_12 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01797_ ) );
OR2_X1 _09514_ ( .A1(fanout_net_12 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01798_ ) );
OAI211_X1 _09515_ ( .A(_01798_ ), .B(fanout_net_20 ), .C1(_01688_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01799_ ) );
NAND3_X1 _09516_ ( .A1(_01797_ ), .A2(_01720_ ), .A3(_01799_ ), .ZN(_01800_ ) );
MUX2_X1 _09517_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01801_ ) );
MUX2_X1 _09518_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01802_ ) );
MUX2_X1 _09519_ ( .A(_01801_ ), .B(_01802_ ), .S(_01737_ ), .Z(_01803_ ) );
OAI211_X1 _09520_ ( .A(_01712_ ), .B(_01800_ ), .C1(_01803_ ), .C2(_01771_ ), .ZN(_01804_ ) );
OR2_X1 _09521_ ( .A1(_01698_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01805_ ) );
OAI211_X1 _09522_ ( .A(_01805_ ), .B(fanout_net_20 ), .C1(fanout_net_12 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01806_ ) );
OR2_X1 _09523_ ( .A1(_01698_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01807_ ) );
OAI211_X1 _09524_ ( .A(_01807_ ), .B(_01777_ ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01808_ ) );
NAND3_X1 _09525_ ( .A1(_01806_ ), .A2(_01808_ ), .A3(fanout_net_23 ), .ZN(_01809_ ) );
MUX2_X1 _09526_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01810_ ) );
MUX2_X1 _09527_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01811_ ) );
MUX2_X1 _09528_ ( .A(_01810_ ), .B(_01811_ ), .S(fanout_net_20 ), .Z(_01812_ ) );
OAI211_X1 _09529_ ( .A(fanout_net_24 ), .B(_01809_ ), .C1(_01812_ ), .C2(fanout_net_23 ), .ZN(_01813_ ) );
OAI211_X1 _09530_ ( .A(_01804_ ), .B(_01813_ ), .C1(_01759_ ), .C2(_01761_ ), .ZN(_01814_ ) );
OR3_X4 _09531_ ( .A1(_01726_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01758_ ), .ZN(_01815_ ) );
NAND2_X2 _09532_ ( .A1(_01814_ ), .A2(_01815_ ), .ZN(_01816_ ) );
OR2_X1 _09533_ ( .A1(_01816_ ), .A2(\ID_EX_imm [23] ), .ZN(_01817_ ) );
NAND2_X1 _09534_ ( .A1(_01816_ ), .A2(\ID_EX_imm [23] ), .ZN(_01818_ ) );
AND3_X1 _09535_ ( .A1(_01795_ ), .A2(_01817_ ), .A3(_01818_ ), .ZN(_01819_ ) );
BUF_X4 _09536_ ( .A(_01687_ ), .Z(_01820_ ) );
OR2_X1 _09537_ ( .A1(_01820_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01821_ ) );
OAI211_X1 _09538_ ( .A(_01821_ ), .B(_01738_ ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01822_ ) );
BUF_X4 _09539_ ( .A(_01687_ ), .Z(_01823_ ) );
OR2_X1 _09540_ ( .A1(_01823_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01824_ ) );
OAI211_X1 _09541_ ( .A(_01824_ ), .B(fanout_net_20 ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01825_ ) );
NAND3_X1 _09542_ ( .A1(_01822_ ), .A2(_01825_ ), .A3(_01779_ ), .ZN(_01826_ ) );
MUX2_X1 _09543_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01827_ ) );
MUX2_X1 _09544_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01828_ ) );
MUX2_X1 _09545_ ( .A(_01827_ ), .B(_01828_ ), .S(_01696_ ), .Z(_01829_ ) );
OAI211_X1 _09546_ ( .A(_01713_ ), .B(_01826_ ), .C1(_01829_ ), .C2(_01721_ ), .ZN(_01830_ ) );
OR2_X1 _09547_ ( .A1(_01823_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01831_ ) );
OAI211_X1 _09548_ ( .A(_01831_ ), .B(fanout_net_20 ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01832_ ) );
OR2_X1 _09549_ ( .A1(_01823_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01833_ ) );
BUF_X4 _09550_ ( .A(_01737_ ), .Z(_01834_ ) );
OAI211_X1 _09551_ ( .A(_01833_ ), .B(_01834_ ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01835_ ) );
NAND3_X1 _09552_ ( .A1(_01832_ ), .A2(_01835_ ), .A3(fanout_net_23 ), .ZN(_01836_ ) );
MUX2_X1 _09553_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01837_ ) );
MUX2_X1 _09554_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01838_ ) );
MUX2_X1 _09555_ ( .A(_01837_ ), .B(_01838_ ), .S(fanout_net_20 ), .Z(_01839_ ) );
OAI211_X1 _09556_ ( .A(fanout_net_24 ), .B(_01836_ ), .C1(_01839_ ), .C2(fanout_net_23 ), .ZN(_01840_ ) );
OAI211_X1 _09557_ ( .A(_01830_ ), .B(_01840_ ), .C1(_01730_ ), .C2(_01727_ ), .ZN(_01841_ ) );
OR3_X4 _09558_ ( .A1(_01790_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01729_ ), .ZN(_01842_ ) );
NAND2_X4 _09559_ ( .A1(_01841_ ), .A2(_01842_ ), .ZN(_01843_ ) );
INV_X1 _09560_ ( .A(\ID_EX_imm [21] ), .ZN(_01844_ ) );
XNOR2_X1 _09561_ ( .A(_01843_ ), .B(_01844_ ), .ZN(_01845_ ) );
BUF_X4 _09562_ ( .A(_01767_ ), .Z(_01846_ ) );
OR2_X1 _09563_ ( .A1(_01846_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01847_ ) );
BUF_X4 _09564_ ( .A(_01696_ ), .Z(_01848_ ) );
OAI211_X1 _09565_ ( .A(_01847_ ), .B(_01848_ ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01849_ ) );
BUF_X4 _09566_ ( .A(_01771_ ), .Z(_01850_ ) );
OR2_X1 _09567_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01851_ ) );
OAI211_X1 _09568_ ( .A(_01851_ ), .B(fanout_net_20 ), .C1(_01700_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01852_ ) );
NAND3_X1 _09569_ ( .A1(_01849_ ), .A2(_01850_ ), .A3(_01852_ ), .ZN(_01853_ ) );
MUX2_X1 _09570_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01854_ ) );
MUX2_X1 _09571_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01855_ ) );
MUX2_X1 _09572_ ( .A(_01854_ ), .B(_01855_ ), .S(_01697_ ), .Z(_01856_ ) );
OAI211_X1 _09573_ ( .A(fanout_net_24 ), .B(_01853_ ), .C1(_01856_ ), .C2(_01722_ ), .ZN(_01857_ ) );
OR2_X1 _09574_ ( .A1(_01699_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01858_ ) );
OAI211_X1 _09575_ ( .A(_01858_ ), .B(_01848_ ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01859_ ) );
OR2_X1 _09576_ ( .A1(_01699_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01860_ ) );
OAI211_X1 _09577_ ( .A(_01860_ ), .B(fanout_net_20 ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01861_ ) );
NAND3_X1 _09578_ ( .A1(_01859_ ), .A2(_01861_ ), .A3(_01850_ ), .ZN(_01862_ ) );
MUX2_X1 _09579_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01863_ ) );
MUX2_X1 _09580_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01864_ ) );
MUX2_X1 _09581_ ( .A(_01863_ ), .B(_01864_ ), .S(_01697_ ), .Z(_01865_ ) );
OAI211_X1 _09582_ ( .A(_01714_ ), .B(_01862_ ), .C1(_01865_ ), .C2(_01722_ ), .ZN(_01866_ ) );
OAI211_X1 _09583_ ( .A(_01857_ ), .B(_01866_ ), .C1(_01760_ ), .C2(_01762_ ), .ZN(_01867_ ) );
OR3_X4 _09584_ ( .A1(_01727_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01730_ ), .ZN(_01868_ ) );
NAND2_X2 _09585_ ( .A1(_01867_ ), .A2(_01868_ ), .ZN(_01869_ ) );
INV_X1 _09586_ ( .A(\ID_EX_imm [20] ), .ZN(_01870_ ) );
XNOR2_X1 _09587_ ( .A(_01869_ ), .B(_01870_ ), .ZN(_01871_ ) );
AND2_X1 _09588_ ( .A1(_01845_ ), .A2(_01871_ ), .ZN(_01872_ ) );
AND2_X1 _09589_ ( .A1(_01819_ ), .A2(_01872_ ), .ZN(_01873_ ) );
INV_X1 _09590_ ( .A(_01873_ ), .ZN(_01874_ ) );
OR2_X1 _09591_ ( .A1(_01820_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01875_ ) );
OAI211_X1 _09592_ ( .A(_01875_ ), .B(_01738_ ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01876_ ) );
OR2_X1 _09593_ ( .A1(_01823_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01877_ ) );
OAI211_X1 _09594_ ( .A(_01877_ ), .B(fanout_net_20 ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01878_ ) );
NAND3_X1 _09595_ ( .A1(_01876_ ), .A2(_01878_ ), .A3(_01779_ ), .ZN(_01879_ ) );
MUX2_X1 _09596_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01880_ ) );
MUX2_X1 _09597_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01881_ ) );
MUX2_X1 _09598_ ( .A(_01880_ ), .B(_01881_ ), .S(_01834_ ), .Z(_01882_ ) );
OAI211_X1 _09599_ ( .A(_01713_ ), .B(_01879_ ), .C1(_01882_ ), .C2(_01721_ ), .ZN(_01883_ ) );
OR2_X1 _09600_ ( .A1(_01820_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01884_ ) );
OAI211_X1 _09601_ ( .A(_01884_ ), .B(fanout_net_20 ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01885_ ) );
OR2_X1 _09602_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01886_ ) );
OAI211_X1 _09603_ ( .A(_01886_ ), .B(_01834_ ), .C1(_01846_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01887_ ) );
NAND3_X1 _09604_ ( .A1(_01885_ ), .A2(fanout_net_23 ), .A3(_01887_ ), .ZN(_01888_ ) );
MUX2_X1 _09605_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01889_ ) );
MUX2_X1 _09606_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01890_ ) );
MUX2_X1 _09607_ ( .A(_01889_ ), .B(_01890_ ), .S(fanout_net_20 ), .Z(_01891_ ) );
OAI211_X1 _09608_ ( .A(fanout_net_24 ), .B(_01888_ ), .C1(_01891_ ), .C2(fanout_net_23 ), .ZN(_01892_ ) );
OAI211_X1 _09609_ ( .A(_01883_ ), .B(_01892_ ), .C1(_01730_ ), .C2(_01727_ ), .ZN(_01893_ ) );
OR3_X4 _09610_ ( .A1(_01790_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01729_ ), .ZN(_01894_ ) );
NAND2_X2 _09611_ ( .A1(_01893_ ), .A2(_01894_ ), .ZN(_01895_ ) );
INV_X1 _09612_ ( .A(\ID_EX_imm [18] ), .ZN(_01896_ ) );
XNOR2_X1 _09613_ ( .A(_01895_ ), .B(_01896_ ), .ZN(_01897_ ) );
OR2_X1 _09614_ ( .A1(_01820_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01898_ ) );
OAI211_X1 _09615_ ( .A(_01898_ ), .B(_01738_ ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01899_ ) );
OR2_X1 _09616_ ( .A1(_01820_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01900_ ) );
OAI211_X1 _09617_ ( .A(_01900_ ), .B(fanout_net_20 ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01901_ ) );
NAND3_X1 _09618_ ( .A1(_01899_ ), .A2(_01901_ ), .A3(_01779_ ), .ZN(_01902_ ) );
MUX2_X1 _09619_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01903_ ) );
MUX2_X1 _09620_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01904_ ) );
MUX2_X1 _09621_ ( .A(_01903_ ), .B(_01904_ ), .S(_01834_ ), .Z(_01905_ ) );
OAI211_X1 _09622_ ( .A(_01713_ ), .B(_01902_ ), .C1(_01905_ ), .C2(_01721_ ), .ZN(_01906_ ) );
OR2_X1 _09623_ ( .A1(_01820_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01907_ ) );
OAI211_X1 _09624_ ( .A(_01907_ ), .B(fanout_net_20 ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01908_ ) );
OR2_X1 _09625_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01909_ ) );
OAI211_X1 _09626_ ( .A(_01909_ ), .B(_01834_ ), .C1(_01846_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01910_ ) );
NAND3_X1 _09627_ ( .A1(_01908_ ), .A2(fanout_net_23 ), .A3(_01910_ ), .ZN(_01911_ ) );
MUX2_X1 _09628_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01912_ ) );
MUX2_X1 _09629_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01913_ ) );
MUX2_X1 _09630_ ( .A(_01912_ ), .B(_01913_ ), .S(fanout_net_20 ), .Z(_01914_ ) );
OAI211_X1 _09631_ ( .A(fanout_net_24 ), .B(_01911_ ), .C1(_01914_ ), .C2(fanout_net_23 ), .ZN(_01915_ ) );
OAI211_X1 _09632_ ( .A(_01906_ ), .B(_01915_ ), .C1(_01730_ ), .C2(_01727_ ), .ZN(_01916_ ) );
OR3_X1 _09633_ ( .A1(_01790_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01729_ ), .ZN(_01917_ ) );
NAND2_X2 _09634_ ( .A1(_01916_ ), .A2(_01917_ ), .ZN(_01918_ ) );
INV_X1 _09635_ ( .A(\ID_EX_imm [19] ), .ZN(_01919_ ) );
XNOR2_X1 _09636_ ( .A(_01918_ ), .B(_01919_ ), .ZN(_01920_ ) );
AND2_X1 _09637_ ( .A1(_01897_ ), .A2(_01920_ ), .ZN(_01921_ ) );
OR2_X1 _09638_ ( .A1(_01699_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01922_ ) );
OAI211_X1 _09639_ ( .A(_01922_ ), .B(fanout_net_20 ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01923_ ) );
OR2_X1 _09640_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01924_ ) );
OAI211_X1 _09641_ ( .A(_01924_ ), .B(_01697_ ), .C1(_01700_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01925_ ) );
NAND3_X1 _09642_ ( .A1(_01923_ ), .A2(_01721_ ), .A3(_01925_ ), .ZN(_01926_ ) );
MUX2_X1 _09643_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01927_ ) );
MUX2_X1 _09644_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01928_ ) );
MUX2_X1 _09645_ ( .A(_01927_ ), .B(_01928_ ), .S(_01697_ ), .Z(_01929_ ) );
OAI211_X1 _09646_ ( .A(fanout_net_24 ), .B(_01926_ ), .C1(_01929_ ), .C2(_01850_ ), .ZN(_01930_ ) );
NOR2_X1 _09647_ ( .A1(_01689_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01931_ ) );
OAI21_X1 _09648_ ( .A(fanout_net_20 ), .B1(fanout_net_14 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01932_ ) );
NOR2_X1 _09649_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01933_ ) );
OAI21_X1 _09650_ ( .A(_01738_ ), .B1(_01689_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01934_ ) );
OAI221_X1 _09651_ ( .A(_01721_ ), .B1(_01931_ ), .B2(_01932_ ), .C1(_01933_ ), .C2(_01934_ ), .ZN(_01935_ ) );
MUX2_X1 _09652_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01936_ ) );
MUX2_X1 _09653_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01937_ ) );
MUX2_X1 _09654_ ( .A(_01936_ ), .B(_01937_ ), .S(_01738_ ), .Z(_01938_ ) );
OAI211_X1 _09655_ ( .A(_01714_ ), .B(_01935_ ), .C1(_01938_ ), .C2(_01850_ ), .ZN(_01939_ ) );
OAI211_X1 _09656_ ( .A(_01930_ ), .B(_01939_ ), .C1(_01760_ ), .C2(_01762_ ), .ZN(_01940_ ) );
OR3_X4 _09657_ ( .A1(_01727_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01759_ ), .ZN(_01941_ ) );
NAND2_X2 _09658_ ( .A1(_01940_ ), .A2(_01941_ ), .ZN(_01942_ ) );
INV_X1 _09659_ ( .A(\ID_EX_imm [17] ), .ZN(_01943_ ) );
XNOR2_X1 _09660_ ( .A(_01942_ ), .B(_01943_ ), .ZN(_01944_ ) );
OR2_X1 _09661_ ( .A1(_01688_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01945_ ) );
OAI211_X1 _09662_ ( .A(_01945_ ), .B(_01738_ ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01946_ ) );
OR2_X1 _09663_ ( .A1(_01688_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01947_ ) );
OAI211_X1 _09664_ ( .A(_01947_ ), .B(fanout_net_20 ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01948_ ) );
NAND3_X1 _09665_ ( .A1(_01946_ ), .A2(_01948_ ), .A3(_01779_ ), .ZN(_01949_ ) );
MUX2_X1 _09666_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01950_ ) );
MUX2_X1 _09667_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01951_ ) );
MUX2_X1 _09668_ ( .A(_01950_ ), .B(_01951_ ), .S(_01834_ ), .Z(_01952_ ) );
OAI211_X1 _09669_ ( .A(_01713_ ), .B(_01949_ ), .C1(_01952_ ), .C2(_01850_ ), .ZN(_01953_ ) );
OR2_X1 _09670_ ( .A1(_01688_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01954_ ) );
OAI211_X1 _09671_ ( .A(_01954_ ), .B(fanout_net_20 ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01955_ ) );
OR2_X1 _09672_ ( .A1(_01688_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01956_ ) );
OAI211_X1 _09673_ ( .A(_01956_ ), .B(_01738_ ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01957_ ) );
NAND3_X1 _09674_ ( .A1(_01955_ ), .A2(_01957_ ), .A3(fanout_net_23 ), .ZN(_01958_ ) );
MUX2_X1 _09675_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01959_ ) );
MUX2_X1 _09676_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01960_ ) );
MUX2_X1 _09677_ ( .A(_01959_ ), .B(_01960_ ), .S(fanout_net_20 ), .Z(_01961_ ) );
OAI211_X1 _09678_ ( .A(fanout_net_24 ), .B(_01958_ ), .C1(_01961_ ), .C2(fanout_net_23 ), .ZN(_01962_ ) );
OAI211_X1 _09679_ ( .A(_01953_ ), .B(_01962_ ), .C1(_01730_ ), .C2(_01727_ ), .ZN(_01963_ ) );
OR3_X4 _09680_ ( .A1(_01790_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01759_ ), .ZN(_01964_ ) );
NAND2_X4 _09681_ ( .A1(_01963_ ), .A2(_01964_ ), .ZN(_01965_ ) );
INV_X1 _09682_ ( .A(\ID_EX_imm [16] ), .ZN(_01966_ ) );
XNOR2_X1 _09683_ ( .A(_01965_ ), .B(_01966_ ), .ZN(_01967_ ) );
NAND3_X1 _09684_ ( .A1(_01921_ ), .A2(_01944_ ), .A3(_01967_ ), .ZN(_01968_ ) );
INV_X1 _09685_ ( .A(\ID_EX_imm [2] ), .ZN(_01969_ ) );
OR2_X1 _09686_ ( .A1(_01686_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01970_ ) );
OAI211_X1 _09687_ ( .A(_01970_ ), .B(_01736_ ), .C1(fanout_net_14 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01971_ ) );
OR2_X1 _09688_ ( .A1(_01686_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01972_ ) );
OAI211_X1 _09689_ ( .A(_01972_ ), .B(fanout_net_20 ), .C1(fanout_net_14 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01973_ ) );
NAND3_X1 _09690_ ( .A1(_01971_ ), .A2(_01973_ ), .A3(_01719_ ), .ZN(_01974_ ) );
MUX2_X1 _09691_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01975_ ) );
MUX2_X1 _09692_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01976_ ) );
MUX2_X1 _09693_ ( .A(_01975_ ), .B(_01976_ ), .S(_01736_ ), .Z(_01977_ ) );
OAI211_X1 _09694_ ( .A(fanout_net_24 ), .B(_01974_ ), .C1(_01977_ ), .C2(_01770_ ), .ZN(_01978_ ) );
BUF_X2 _09695_ ( .A(_01685_ ), .Z(_01979_ ) );
NOR2_X1 _09696_ ( .A1(_01979_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01980_ ) );
OAI21_X1 _09697_ ( .A(fanout_net_20 ), .B1(fanout_net_14 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01981_ ) );
NOR2_X1 _09698_ ( .A1(fanout_net_14 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01982_ ) );
OAI21_X1 _09699_ ( .A(_01736_ ), .B1(_01979_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01983_ ) );
OAI221_X1 _09700_ ( .A(_01719_ ), .B1(_01980_ ), .B2(_01981_ ), .C1(_01982_ ), .C2(_01983_ ), .ZN(_01984_ ) );
MUX2_X1 _09701_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01985_ ) );
MUX2_X1 _09702_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01986_ ) );
MUX2_X1 _09703_ ( .A(_01985_ ), .B(_01986_ ), .S(_01736_ ), .Z(_01987_ ) );
OAI211_X1 _09704_ ( .A(_01712_ ), .B(_01984_ ), .C1(_01987_ ), .C2(_01770_ ), .ZN(_01988_ ) );
OAI211_X1 _09705_ ( .A(_01978_ ), .B(_01988_ ), .C1(_01728_ ), .C2(_01725_ ), .ZN(_01989_ ) );
OR3_X4 _09706_ ( .A1(_01725_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01728_ ), .ZN(_01990_ ) );
AOI21_X1 _09707_ ( .A(_01969_ ), .B1(_01989_ ), .B2(_01990_ ), .ZN(_01991_ ) );
OR2_X1 _09708_ ( .A1(_01685_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01992_ ) );
OAI211_X1 _09709_ ( .A(_01992_ ), .B(_01694_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(fanout_net_14 ), .ZN(_01993_ ) );
OR2_X1 _09710_ ( .A1(fanout_net_15 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01994_ ) );
OAI211_X1 _09711_ ( .A(_01994_ ), .B(fanout_net_21 ), .C1(_01685_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01995_ ) );
NAND3_X1 _09712_ ( .A1(_01993_ ), .A2(_01718_ ), .A3(_01995_ ), .ZN(_01996_ ) );
MUX2_X1 _09713_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01997_ ) );
MUX2_X1 _09714_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01998_ ) );
MUX2_X1 _09715_ ( .A(_01997_ ), .B(_01998_ ), .S(_01693_ ), .Z(_01999_ ) );
OAI211_X1 _09716_ ( .A(_01711_ ), .B(_01996_ ), .C1(_01999_ ), .C2(_01719_ ), .ZN(_02000_ ) );
OR2_X1 _09717_ ( .A1(_01685_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02001_ ) );
OAI211_X1 _09718_ ( .A(_02001_ ), .B(fanout_net_21 ), .C1(fanout_net_15 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02002_ ) );
OR2_X1 _09719_ ( .A1(_01684_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02003_ ) );
OAI211_X1 _09720_ ( .A(_02003_ ), .B(_01693_ ), .C1(fanout_net_15 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02004_ ) );
NAND3_X1 _09721_ ( .A1(_02002_ ), .A2(_02004_ ), .A3(fanout_net_23 ), .ZN(_02005_ ) );
MUX2_X1 _09722_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02006_ ) );
MUX2_X1 _09723_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02007_ ) );
MUX2_X1 _09724_ ( .A(_02006_ ), .B(_02007_ ), .S(fanout_net_21 ), .Z(_02008_ ) );
OAI211_X1 _09725_ ( .A(fanout_net_24 ), .B(_02005_ ), .C1(_02008_ ), .C2(fanout_net_23 ), .ZN(_02009_ ) );
NAND2_X1 _09726_ ( .A1(_02000_ ), .A2(_02009_ ), .ZN(_02010_ ) );
NAND2_X2 _09727_ ( .A1(_02010_ ), .A2(_01683_ ), .ZN(_02011_ ) );
INV_X8 _09728_ ( .A(_01681_ ), .ZN(_02012_ ) );
NAND4_X1 _09729_ ( .A1(_02012_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01671_ ), .A4(_01666_ ), .ZN(_02013_ ) );
AND2_X4 _09730_ ( .A1(_02011_ ), .A2(_02013_ ), .ZN(_02014_ ) );
INV_X1 _09731_ ( .A(\ID_EX_imm [1] ), .ZN(_02015_ ) );
XNOR2_X1 _09732_ ( .A(_02014_ ), .B(_02015_ ), .ZN(_02016_ ) );
OR2_X1 _09733_ ( .A1(_01685_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02017_ ) );
OAI211_X1 _09734_ ( .A(_02017_ ), .B(_01694_ ), .C1(fanout_net_15 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02018_ ) );
OR2_X1 _09735_ ( .A1(_01685_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02019_ ) );
OAI211_X1 _09736_ ( .A(_02019_ ), .B(fanout_net_21 ), .C1(fanout_net_15 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02020_ ) );
NAND3_X1 _09737_ ( .A1(_02018_ ), .A2(_02020_ ), .A3(_01719_ ), .ZN(_02021_ ) );
MUX2_X1 _09738_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02022_ ) );
MUX2_X1 _09739_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02023_ ) );
MUX2_X1 _09740_ ( .A(_02022_ ), .B(_02023_ ), .S(_01694_ ), .Z(_02024_ ) );
OAI211_X1 _09741_ ( .A(_01711_ ), .B(_02021_ ), .C1(_02024_ ), .C2(_01719_ ), .ZN(_02025_ ) );
OR2_X1 _09742_ ( .A1(_01685_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02026_ ) );
OAI211_X1 _09743_ ( .A(_02026_ ), .B(fanout_net_21 ), .C1(fanout_net_15 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02027_ ) );
OR2_X1 _09744_ ( .A1(fanout_net_15 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02028_ ) );
OAI211_X1 _09745_ ( .A(_02028_ ), .B(_01694_ ), .C1(_01686_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02029_ ) );
NAND3_X1 _09746_ ( .A1(_02027_ ), .A2(fanout_net_23 ), .A3(_02029_ ), .ZN(_02030_ ) );
MUX2_X1 _09747_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02031_ ) );
MUX2_X1 _09748_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02032_ ) );
MUX2_X1 _09749_ ( .A(_02031_ ), .B(_02032_ ), .S(fanout_net_21 ), .Z(_02033_ ) );
OAI211_X1 _09750_ ( .A(fanout_net_24 ), .B(_02030_ ), .C1(_02033_ ), .C2(fanout_net_23 ), .ZN(_02034_ ) );
NAND2_X1 _09751_ ( .A1(_02025_ ), .A2(_02034_ ), .ZN(_02035_ ) );
NAND2_X1 _09752_ ( .A1(_02035_ ), .A2(_01683_ ), .ZN(_02036_ ) );
BUF_X4 _09753_ ( .A(_02012_ ), .Z(_02037_ ) );
NAND4_X1 _09754_ ( .A1(_02037_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_01671_ ), .A4(_01666_ ), .ZN(_02038_ ) );
AND3_X1 _09755_ ( .A1(_02036_ ), .A2(\ID_EX_imm [0] ), .A3(_02038_ ), .ZN(_02039_ ) );
NAND2_X1 _09756_ ( .A1(_02016_ ), .A2(_02039_ ), .ZN(_02040_ ) );
INV_X4 _09757_ ( .A(_02014_ ), .ZN(_02041_ ) );
OR2_X4 _09758_ ( .A1(_02041_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02042_ ) );
AND2_X2 _09759_ ( .A1(_02040_ ), .A2(_02042_ ), .ZN(_02043_ ) );
INV_X2 _09760_ ( .A(_02043_ ), .ZN(_02044_ ) );
NAND2_X1 _09761_ ( .A1(_01989_ ), .A2(_01990_ ), .ZN(_02045_ ) );
XNOR2_X1 _09762_ ( .A(_02045_ ), .B(_01969_ ), .ZN(_02046_ ) );
AOI21_X2 _09763_ ( .A(_01991_ ), .B1(_02044_ ), .B2(_02046_ ), .ZN(_02047_ ) );
OR2_X1 _09764_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02048_ ) );
OAI211_X1 _09765_ ( .A(_02048_ ), .B(fanout_net_21 ), .C1(_01698_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02049_ ) );
INV_X1 _09766_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02050_ ) );
INV_X1 _09767_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02051_ ) );
MUX2_X1 _09768_ ( .A(_02050_ ), .B(_02051_ ), .S(fanout_net_15 ), .Z(_02052_ ) );
OAI211_X1 _09769_ ( .A(_02049_ ), .B(_01770_ ), .C1(_02052_ ), .C2(fanout_net_21 ), .ZN(_02053_ ) );
MUX2_X1 _09770_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02054_ ) );
MUX2_X1 _09771_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02055_ ) );
MUX2_X1 _09772_ ( .A(_02054_ ), .B(_02055_ ), .S(_01736_ ), .Z(_02056_ ) );
OAI211_X1 _09773_ ( .A(fanout_net_24 ), .B(_02053_ ), .C1(_02056_ ), .C2(_01770_ ), .ZN(_02057_ ) );
OR2_X1 _09774_ ( .A1(_01686_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02058_ ) );
OAI211_X1 _09775_ ( .A(_02058_ ), .B(fanout_net_21 ), .C1(fanout_net_15 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02059_ ) );
OR2_X1 _09776_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02060_ ) );
OAI211_X1 _09777_ ( .A(_02060_ ), .B(_01736_ ), .C1(_01698_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02061_ ) );
NAND3_X1 _09778_ ( .A1(_02059_ ), .A2(_01770_ ), .A3(_02061_ ), .ZN(_02062_ ) );
MUX2_X1 _09779_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02063_ ) );
MUX2_X1 _09780_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02064_ ) );
MUX2_X1 _09781_ ( .A(_02063_ ), .B(_02064_ ), .S(_01736_ ), .Z(_02065_ ) );
OAI211_X1 _09782_ ( .A(_01712_ ), .B(_02062_ ), .C1(_02065_ ), .C2(_01770_ ), .ZN(_02066_ ) );
OAI211_X1 _09783_ ( .A(_02057_ ), .B(_02066_ ), .C1(_01758_ ), .C2(_01725_ ), .ZN(_02067_ ) );
OR3_X1 _09784_ ( .A1(_01725_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01728_ ), .ZN(_02068_ ) );
NAND2_X2 _09785_ ( .A1(_02067_ ), .A2(_02068_ ), .ZN(_02069_ ) );
XNOR2_X1 _09786_ ( .A(_02069_ ), .B(\ID_EX_imm [3] ), .ZN(_02070_ ) );
NOR2_X2 _09787_ ( .A1(_02047_ ), .A2(_02070_ ), .ZN(_02071_ ) );
AOI21_X1 _09788_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B1(_02067_ ), .B2(_02068_ ), .ZN(_02072_ ) );
NOR2_X2 _09789_ ( .A1(_02071_ ), .A2(_02072_ ), .ZN(_02073_ ) );
OR2_X1 _09790_ ( .A1(_01685_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02074_ ) );
OAI211_X1 _09791_ ( .A(_02074_ ), .B(_01694_ ), .C1(fanout_net_15 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02075_ ) );
NOR2_X1 _09792_ ( .A1(_01686_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02076_ ) );
OAI21_X1 _09793_ ( .A(fanout_net_21 ), .B1(fanout_net_15 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02077_ ) );
OAI211_X1 _09794_ ( .A(_02075_ ), .B(fanout_net_23 ), .C1(_02076_ ), .C2(_02077_ ), .ZN(_02078_ ) );
MUX2_X1 _09795_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02079_ ) );
MUX2_X1 _09796_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02080_ ) );
MUX2_X1 _09797_ ( .A(_02079_ ), .B(_02080_ ), .S(fanout_net_21 ), .Z(_02081_ ) );
OAI211_X1 _09798_ ( .A(_02078_ ), .B(fanout_net_24 ), .C1(_02081_ ), .C2(fanout_net_23 ), .ZN(_02082_ ) );
OR2_X1 _09799_ ( .A1(_01685_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02083_ ) );
OAI211_X1 _09800_ ( .A(_02083_ ), .B(_01694_ ), .C1(fanout_net_15 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02084_ ) );
OR2_X1 _09801_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02085_ ) );
OAI211_X1 _09802_ ( .A(_02085_ ), .B(fanout_net_21 ), .C1(_01686_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02086_ ) );
NAND3_X1 _09803_ ( .A1(_02084_ ), .A2(_01719_ ), .A3(_02086_ ), .ZN(_02087_ ) );
MUX2_X1 _09804_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02088_ ) );
MUX2_X1 _09805_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02089_ ) );
MUX2_X1 _09806_ ( .A(_02088_ ), .B(_02089_ ), .S(_01694_ ), .Z(_02090_ ) );
OAI211_X1 _09807_ ( .A(_01711_ ), .B(_02087_ ), .C1(_02090_ ), .C2(_01719_ ), .ZN(_02091_ ) );
NAND2_X1 _09808_ ( .A1(_02082_ ), .A2(_02091_ ), .ZN(_02092_ ) );
NAND2_X1 _09809_ ( .A1(_02092_ ), .A2(_01683_ ), .ZN(_02093_ ) );
NAND4_X1 _09810_ ( .A1(_02012_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01671_ ), .A4(_01666_ ), .ZN(_02094_ ) );
AND2_X1 _09811_ ( .A1(_02093_ ), .A2(_02094_ ), .ZN(_02095_ ) );
BUF_X2 _09812_ ( .A(_02095_ ), .Z(_02096_ ) );
XNOR2_X1 _09813_ ( .A(_02096_ ), .B(\ID_EX_imm [5] ), .ZN(_02097_ ) );
OR2_X1 _09814_ ( .A1(fanout_net_16 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02098_ ) );
OAI211_X1 _09815_ ( .A(_02098_ ), .B(_01737_ ), .C1(_01688_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02099_ ) );
OR2_X1 _09816_ ( .A1(fanout_net_16 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02100_ ) );
OAI211_X1 _09817_ ( .A(_02100_ ), .B(fanout_net_21 ), .C1(_01820_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02101_ ) );
NAND3_X1 _09818_ ( .A1(_02099_ ), .A2(_02101_ ), .A3(_01720_ ), .ZN(_02102_ ) );
MUX2_X1 _09819_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02103_ ) );
MUX2_X1 _09820_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02104_ ) );
MUX2_X1 _09821_ ( .A(_02103_ ), .B(_02104_ ), .S(_01695_ ), .Z(_02105_ ) );
OAI211_X1 _09822_ ( .A(_01712_ ), .B(_02102_ ), .C1(_02105_ ), .C2(_01771_ ), .ZN(_02106_ ) );
OR2_X1 _09823_ ( .A1(_01687_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02107_ ) );
OAI211_X1 _09824_ ( .A(_02107_ ), .B(fanout_net_21 ), .C1(fanout_net_16 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02108_ ) );
OR2_X1 _09825_ ( .A1(fanout_net_16 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02109_ ) );
OAI211_X1 _09826_ ( .A(_02109_ ), .B(_01737_ ), .C1(_01820_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02110_ ) );
NAND3_X1 _09827_ ( .A1(_02108_ ), .A2(fanout_net_23 ), .A3(_02110_ ), .ZN(_02111_ ) );
MUX2_X1 _09828_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02112_ ) );
MUX2_X1 _09829_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02113_ ) );
MUX2_X1 _09830_ ( .A(_02112_ ), .B(_02113_ ), .S(fanout_net_21 ), .Z(_02114_ ) );
OAI211_X1 _09831_ ( .A(fanout_net_24 ), .B(_02111_ ), .C1(_02114_ ), .C2(fanout_net_23 ), .ZN(_02115_ ) );
OAI211_X1 _09832_ ( .A(_02106_ ), .B(_02115_ ), .C1(_01729_ ), .C2(_01761_ ), .ZN(_02116_ ) );
OR3_X4 _09833_ ( .A1(_01726_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01758_ ), .ZN(_02117_ ) );
NAND2_X2 _09834_ ( .A1(_02116_ ), .A2(_02117_ ), .ZN(_02118_ ) );
INV_X1 _09835_ ( .A(\ID_EX_imm [4] ), .ZN(_02119_ ) );
XNOR2_X1 _09836_ ( .A(_02118_ ), .B(_02119_ ), .ZN(_02120_ ) );
INV_X1 _09837_ ( .A(_02120_ ), .ZN(_02121_ ) );
NOR3_X2 _09838_ ( .A1(_02073_ ), .A2(_02097_ ), .A3(_02121_ ), .ZN(_02122_ ) );
INV_X4 _09839_ ( .A(_02118_ ), .ZN(_02123_ ) );
NOR3_X1 _09840_ ( .A1(_02097_ ), .A2(_02119_ ), .A3(_02123_ ), .ZN(_02124_ ) );
INV_X1 _09841_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02125_ ) );
AOI21_X1 _09842_ ( .A(_02124_ ), .B1(_02125_ ), .B2(_02096_ ), .ZN(_02126_ ) );
INV_X1 _09843_ ( .A(_02126_ ), .ZN(_02127_ ) );
NOR2_X2 _09844_ ( .A1(_02122_ ), .A2(_02127_ ), .ZN(_02128_ ) );
NOR2_X1 _09845_ ( .A1(_01979_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02129_ ) );
OAI21_X1 _09846_ ( .A(fanout_net_21 ), .B1(fanout_net_16 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02130_ ) );
NOR2_X1 _09847_ ( .A1(fanout_net_16 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02131_ ) );
OAI21_X1 _09848_ ( .A(_01736_ ), .B1(_01979_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02132_ ) );
OAI221_X1 _09849_ ( .A(_01719_ ), .B1(_02129_ ), .B2(_02130_ ), .C1(_02131_ ), .C2(_02132_ ), .ZN(_02133_ ) );
MUX2_X1 _09850_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02134_ ) );
MUX2_X1 _09851_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02135_ ) );
MUX2_X1 _09852_ ( .A(_02134_ ), .B(_02135_ ), .S(fanout_net_21 ), .Z(_02136_ ) );
OAI211_X1 _09853_ ( .A(fanout_net_24 ), .B(_02133_ ), .C1(_02136_ ), .C2(_01770_ ), .ZN(_02137_ ) );
OR2_X1 _09854_ ( .A1(_01686_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02138_ ) );
OAI211_X1 _09855_ ( .A(_02138_ ), .B(_01736_ ), .C1(fanout_net_16 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02139_ ) );
OR2_X1 _09856_ ( .A1(fanout_net_16 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02140_ ) );
OAI211_X1 _09857_ ( .A(_02140_ ), .B(fanout_net_21 ), .C1(_01979_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02141_ ) );
NAND3_X1 _09858_ ( .A1(_02139_ ), .A2(fanout_net_23 ), .A3(_02141_ ), .ZN(_02142_ ) );
MUX2_X1 _09859_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02143_ ) );
MUX2_X1 _09860_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02144_ ) );
MUX2_X1 _09861_ ( .A(_02143_ ), .B(_02144_ ), .S(_01694_ ), .Z(_02145_ ) );
OAI211_X1 _09862_ ( .A(_01711_ ), .B(_02142_ ), .C1(_02145_ ), .C2(fanout_net_23 ), .ZN(_02146_ ) );
OAI211_X2 _09863_ ( .A(_02137_ ), .B(_02146_ ), .C1(_01728_ ), .C2(_01725_ ), .ZN(_02147_ ) );
OR3_X1 _09864_ ( .A1(_01725_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01728_ ), .ZN(_02148_ ) );
NAND2_X2 _09865_ ( .A1(_02147_ ), .A2(_02148_ ), .ZN(_02149_ ) );
XNOR2_X1 _09866_ ( .A(_02149_ ), .B(\ID_EX_imm [7] ), .ZN(_02150_ ) );
OR2_X1 _09867_ ( .A1(_01979_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02151_ ) );
OAI211_X1 _09868_ ( .A(_02151_ ), .B(_01695_ ), .C1(fanout_net_16 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02152_ ) );
OR2_X1 _09869_ ( .A1(_01979_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02153_ ) );
OAI211_X1 _09870_ ( .A(_02153_ ), .B(fanout_net_21 ), .C1(fanout_net_16 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02154_ ) );
NAND3_X1 _09871_ ( .A1(_02152_ ), .A2(_02154_ ), .A3(_01770_ ), .ZN(_02155_ ) );
MUX2_X1 _09872_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02156_ ) );
MUX2_X1 _09873_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02157_ ) );
MUX2_X1 _09874_ ( .A(_02156_ ), .B(_02157_ ), .S(_01695_ ), .Z(_02158_ ) );
OAI211_X1 _09875_ ( .A(_01712_ ), .B(_02155_ ), .C1(_02158_ ), .C2(_01720_ ), .ZN(_02159_ ) );
OR2_X1 _09876_ ( .A1(_01979_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02160_ ) );
OAI211_X1 _09877_ ( .A(_02160_ ), .B(_01695_ ), .C1(fanout_net_16 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02161_ ) );
OR2_X1 _09878_ ( .A1(fanout_net_16 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02162_ ) );
OAI211_X1 _09879_ ( .A(_02162_ ), .B(fanout_net_21 ), .C1(_01698_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02163_ ) );
NAND3_X1 _09880_ ( .A1(_02161_ ), .A2(fanout_net_23 ), .A3(_02163_ ), .ZN(_02164_ ) );
MUX2_X1 _09881_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02165_ ) );
MUX2_X1 _09882_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02166_ ) );
MUX2_X1 _09883_ ( .A(_02165_ ), .B(_02166_ ), .S(fanout_net_21 ), .Z(_02167_ ) );
OAI211_X1 _09884_ ( .A(fanout_net_24 ), .B(_02164_ ), .C1(_02167_ ), .C2(fanout_net_23 ), .ZN(_02168_ ) );
OAI211_X1 _09885_ ( .A(_02159_ ), .B(_02168_ ), .C1(_01758_ ), .C2(_01726_ ), .ZN(_02169_ ) );
OR3_X1 _09886_ ( .A1(_01725_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01728_ ), .ZN(_02170_ ) );
NAND2_X2 _09887_ ( .A1(_02169_ ), .A2(_02170_ ), .ZN(_02171_ ) );
XOR2_X1 _09888_ ( .A(_02171_ ), .B(\ID_EX_imm [6] ), .Z(_02172_ ) );
INV_X1 _09889_ ( .A(_02172_ ), .ZN(_02173_ ) );
NOR3_X2 _09890_ ( .A1(_02128_ ), .A2(_02150_ ), .A3(_02173_ ), .ZN(_02174_ ) );
AND2_X1 _09891_ ( .A1(_02171_ ), .A2(\ID_EX_imm [6] ), .ZN(_02175_ ) );
INV_X1 _09892_ ( .A(_02175_ ), .ZN(_02176_ ) );
NOR2_X1 _09893_ ( .A1(_02150_ ), .A2(_02176_ ), .ZN(_02177_ ) );
AOI21_X1 _09894_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B1(_02147_ ), .B2(_02148_ ), .ZN(_02178_ ) );
NOR2_X1 _09895_ ( .A1(_02177_ ), .A2(_02178_ ), .ZN(_02179_ ) );
INV_X1 _09896_ ( .A(_02179_ ), .ZN(_02180_ ) );
NOR2_X2 _09897_ ( .A1(_02174_ ), .A2(_02180_ ), .ZN(_02181_ ) );
OR2_X1 _09898_ ( .A1(_01846_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02182_ ) );
OAI211_X1 _09899_ ( .A(_02182_ ), .B(_01848_ ), .C1(fanout_net_16 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02183_ ) );
OR2_X1 _09900_ ( .A1(_01846_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02184_ ) );
OAI211_X1 _09901_ ( .A(_02184_ ), .B(fanout_net_21 ), .C1(fanout_net_16 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02185_ ) );
NAND3_X1 _09902_ ( .A1(_02183_ ), .A2(_02185_ ), .A3(_01850_ ), .ZN(_02186_ ) );
MUX2_X1 _09903_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02187_ ) );
MUX2_X1 _09904_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02188_ ) );
MUX2_X1 _09905_ ( .A(_02187_ ), .B(_02188_ ), .S(_01848_ ), .Z(_02189_ ) );
OAI211_X1 _09906_ ( .A(fanout_net_24 ), .B(_02186_ ), .C1(_02189_ ), .C2(_01722_ ), .ZN(_02190_ ) );
NOR2_X1 _09907_ ( .A1(_01700_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02191_ ) );
OAI21_X1 _09908_ ( .A(fanout_net_21 ), .B1(fanout_net_16 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02192_ ) );
NOR2_X1 _09909_ ( .A1(fanout_net_17 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02193_ ) );
OAI21_X1 _09910_ ( .A(_01848_ ), .B1(_01700_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02194_ ) );
OAI221_X1 _09911_ ( .A(_01850_ ), .B1(_02191_ ), .B2(_02192_ ), .C1(_02193_ ), .C2(_02194_ ), .ZN(_02195_ ) );
MUX2_X1 _09912_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02196_ ) );
MUX2_X1 _09913_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02197_ ) );
MUX2_X1 _09914_ ( .A(_02196_ ), .B(_02197_ ), .S(_01848_ ), .Z(_02198_ ) );
OAI211_X1 _09915_ ( .A(_01714_ ), .B(_02195_ ), .C1(_02198_ ), .C2(_01722_ ), .ZN(_02199_ ) );
OAI211_X1 _09916_ ( .A(_02190_ ), .B(_02199_ ), .C1(_01760_ ), .C2(_01762_ ), .ZN(_02200_ ) );
OR3_X1 _09917_ ( .A1(_01727_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01730_ ), .ZN(_02201_ ) );
NAND2_X4 _09918_ ( .A1(_02200_ ), .A2(_02201_ ), .ZN(_02202_ ) );
INV_X1 _09919_ ( .A(\ID_EX_imm [8] ), .ZN(_02203_ ) );
XNOR2_X1 _09920_ ( .A(_02202_ ), .B(_02203_ ), .ZN(_02204_ ) );
OR2_X1 _09921_ ( .A1(_01979_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02205_ ) );
OAI211_X1 _09922_ ( .A(_02205_ ), .B(fanout_net_21 ), .C1(fanout_net_17 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02206_ ) );
OR2_X1 _09923_ ( .A1(fanout_net_17 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02207_ ) );
OAI211_X1 _09924_ ( .A(_02207_ ), .B(_01695_ ), .C1(_01767_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02208_ ) );
NAND3_X1 _09925_ ( .A1(_02206_ ), .A2(_01770_ ), .A3(_02208_ ), .ZN(_02209_ ) );
MUX2_X1 _09926_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02210_ ) );
MUX2_X1 _09927_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02211_ ) );
MUX2_X1 _09928_ ( .A(_02210_ ), .B(_02211_ ), .S(_01695_ ), .Z(_02212_ ) );
OAI211_X1 _09929_ ( .A(_01712_ ), .B(_02209_ ), .C1(_02212_ ), .C2(_01720_ ), .ZN(_02213_ ) );
OR2_X1 _09930_ ( .A1(_01979_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02214_ ) );
OAI211_X1 _09931_ ( .A(_02214_ ), .B(_01695_ ), .C1(fanout_net_17 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02215_ ) );
OR2_X1 _09932_ ( .A1(fanout_net_17 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02216_ ) );
OAI211_X1 _09933_ ( .A(_02216_ ), .B(fanout_net_21 ), .C1(_01767_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02217_ ) );
NAND3_X1 _09934_ ( .A1(_02215_ ), .A2(fanout_net_23 ), .A3(_02217_ ), .ZN(_02218_ ) );
MUX2_X1 _09935_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02219_ ) );
MUX2_X1 _09936_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02220_ ) );
MUX2_X1 _09937_ ( .A(_02219_ ), .B(_02220_ ), .S(fanout_net_21 ), .Z(_02221_ ) );
OAI211_X1 _09938_ ( .A(fanout_net_24 ), .B(_02218_ ), .C1(_02221_ ), .C2(fanout_net_23 ), .ZN(_02222_ ) );
OAI211_X1 _09939_ ( .A(_02213_ ), .B(_02222_ ), .C1(_01758_ ), .C2(_01726_ ), .ZN(_02223_ ) );
OR3_X1 _09940_ ( .A1(_01725_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01728_ ), .ZN(_02224_ ) );
NAND2_X2 _09941_ ( .A1(_02223_ ), .A2(_02224_ ), .ZN(_02225_ ) );
INV_X1 _09942_ ( .A(\ID_EX_imm [9] ), .ZN(_02226_ ) );
XNOR2_X1 _09943_ ( .A(_02225_ ), .B(_02226_ ), .ZN(_02227_ ) );
AND2_X1 _09944_ ( .A1(_02204_ ), .A2(_02227_ ), .ZN(_02228_ ) );
OR2_X1 _09945_ ( .A1(_01687_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02229_ ) );
OAI211_X1 _09946_ ( .A(_02229_ ), .B(fanout_net_21 ), .C1(fanout_net_17 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02230_ ) );
OR2_X1 _09947_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02231_ ) );
OAI211_X1 _09948_ ( .A(_02231_ ), .B(_01737_ ), .C1(_01820_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02232_ ) );
NAND3_X1 _09949_ ( .A1(_02230_ ), .A2(_01720_ ), .A3(_02232_ ), .ZN(_02233_ ) );
MUX2_X1 _09950_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02234_ ) );
MUX2_X1 _09951_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02235_ ) );
MUX2_X1 _09952_ ( .A(_02234_ ), .B(_02235_ ), .S(_01737_ ), .Z(_02236_ ) );
OAI211_X1 _09953_ ( .A(_01712_ ), .B(_02233_ ), .C1(_02236_ ), .C2(_01771_ ), .ZN(_02237_ ) );
OR2_X1 _09954_ ( .A1(_01687_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02238_ ) );
OAI211_X1 _09955_ ( .A(_02238_ ), .B(_01737_ ), .C1(fanout_net_17 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02239_ ) );
OR2_X1 _09956_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02240_ ) );
OAI211_X1 _09957_ ( .A(_02240_ ), .B(fanout_net_21 ), .C1(_01820_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02241_ ) );
NAND3_X1 _09958_ ( .A1(_02239_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02241_ ), .ZN(_02242_ ) );
MUX2_X1 _09959_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02243_ ) );
MUX2_X1 _09960_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02244_ ) );
MUX2_X1 _09961_ ( .A(_02243_ ), .B(_02244_ ), .S(fanout_net_21 ), .Z(_02245_ ) );
OAI211_X1 _09962_ ( .A(fanout_net_24 ), .B(_02242_ ), .C1(_02245_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02246_ ) );
OAI211_X1 _09963_ ( .A(_02237_ ), .B(_02246_ ), .C1(_01729_ ), .C2(_01726_ ), .ZN(_02247_ ) );
OR3_X1 _09964_ ( .A1(_01726_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01758_ ), .ZN(_02248_ ) );
NAND2_X2 _09965_ ( .A1(_02247_ ), .A2(_02248_ ), .ZN(_02249_ ) );
INV_X1 _09966_ ( .A(\ID_EX_imm [10] ), .ZN(_02250_ ) );
XNOR2_X1 _09967_ ( .A(_02249_ ), .B(_02250_ ), .ZN(_02251_ ) );
OR2_X1 _09968_ ( .A1(_01687_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02252_ ) );
OAI211_X1 _09969_ ( .A(_02252_ ), .B(_01737_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02253_ ) );
OR2_X1 _09970_ ( .A1(_01687_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02254_ ) );
OAI211_X1 _09971_ ( .A(_02254_ ), .B(fanout_net_21 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02255_ ) );
NAND3_X1 _09972_ ( .A1(_02253_ ), .A2(_02255_ ), .A3(_01720_ ), .ZN(_02256_ ) );
MUX2_X1 _09973_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02257_ ) );
MUX2_X1 _09974_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02258_ ) );
MUX2_X1 _09975_ ( .A(_02257_ ), .B(_02258_ ), .S(_01695_ ), .Z(_02259_ ) );
OAI211_X1 _09976_ ( .A(_01712_ ), .B(_02256_ ), .C1(_02259_ ), .C2(_01771_ ), .ZN(_02260_ ) );
OR2_X1 _09977_ ( .A1(_01687_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02261_ ) );
OAI211_X1 _09978_ ( .A(_02261_ ), .B(fanout_net_22 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02262_ ) );
OR2_X1 _09979_ ( .A1(_01687_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02263_ ) );
OAI211_X1 _09980_ ( .A(_02263_ ), .B(_01737_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02264_ ) );
NAND3_X1 _09981_ ( .A1(_02262_ ), .A2(_02264_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02265_ ) );
MUX2_X1 _09982_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02266_ ) );
MUX2_X1 _09983_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02267_ ) );
MUX2_X1 _09984_ ( .A(_02266_ ), .B(_02267_ ), .S(fanout_net_22 ), .Z(_02268_ ) );
OAI211_X1 _09985_ ( .A(fanout_net_24 ), .B(_02265_ ), .C1(_02268_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02269_ ) );
OAI211_X1 _09986_ ( .A(_02260_ ), .B(_02269_ ), .C1(_01729_ ), .C2(_01761_ ), .ZN(_02270_ ) );
OR3_X1 _09987_ ( .A1(_01726_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_01728_ ), .ZN(_02271_ ) );
NAND2_X2 _09988_ ( .A1(_02270_ ), .A2(_02271_ ), .ZN(_02272_ ) );
INV_X1 _09989_ ( .A(\ID_EX_imm [11] ), .ZN(_02273_ ) );
XNOR2_X1 _09990_ ( .A(_02272_ ), .B(_02273_ ), .ZN(_02274_ ) );
AND2_X1 _09991_ ( .A1(_02251_ ), .A2(_02274_ ), .ZN(_02275_ ) );
AND2_X1 _09992_ ( .A1(_02228_ ), .A2(_02275_ ), .ZN(_02276_ ) );
INV_X1 _09993_ ( .A(_02276_ ), .ZN(_02277_ ) );
NOR2_X2 _09994_ ( .A1(_02181_ ), .A2(_02277_ ), .ZN(_02278_ ) );
AND2_X1 _09995_ ( .A1(_02249_ ), .A2(\ID_EX_imm [10] ), .ZN(_02279_ ) );
AND2_X1 _09996_ ( .A1(_02274_ ), .A2(_02279_ ), .ZN(_02280_ ) );
AOI21_X1 _09997_ ( .A(_02280_ ), .B1(\ID_EX_imm [11] ), .B2(_02272_ ), .ZN(_02281_ ) );
AOI21_X1 _09998_ ( .A(_02226_ ), .B1(_02223_ ), .B2(_02224_ ), .ZN(_02282_ ) );
AND2_X1 _09999_ ( .A1(_02202_ ), .A2(\ID_EX_imm [8] ), .ZN(_02283_ ) );
AND2_X1 _10000_ ( .A1(_02227_ ), .A2(_02283_ ), .ZN(_02284_ ) );
OAI21_X1 _10001_ ( .A(_02275_ ), .B1(_02282_ ), .B2(_02284_ ), .ZN(_02285_ ) );
AND2_X1 _10002_ ( .A1(_02281_ ), .A2(_02285_ ), .ZN(_02286_ ) );
INV_X1 _10003_ ( .A(_02286_ ), .ZN(_02287_ ) );
NOR2_X2 _10004_ ( .A1(_02278_ ), .A2(_02287_ ), .ZN(_02288_ ) );
OR2_X1 _10005_ ( .A1(_01767_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02289_ ) );
OAI211_X1 _10006_ ( .A(_02289_ ), .B(_01696_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02290_ ) );
OR2_X1 _10007_ ( .A1(_01767_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02291_ ) );
OAI211_X1 _10008_ ( .A(_02291_ ), .B(fanout_net_22 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02292_ ) );
NAND3_X1 _10009_ ( .A1(_02290_ ), .A2(_02292_ ), .A3(_01771_ ), .ZN(_02293_ ) );
MUX2_X1 _10010_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02294_ ) );
MUX2_X1 _10011_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02295_ ) );
MUX2_X1 _10012_ ( .A(_02294_ ), .B(_02295_ ), .S(_01777_ ), .Z(_02296_ ) );
OAI211_X1 _10013_ ( .A(fanout_net_24 ), .B(_02293_ ), .C1(_02296_ ), .C2(_01779_ ), .ZN(_02297_ ) );
OR2_X1 _10014_ ( .A1(_01767_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02298_ ) );
OAI211_X1 _10015_ ( .A(_02298_ ), .B(_01696_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02299_ ) );
OR2_X1 _10016_ ( .A1(_01767_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02300_ ) );
OAI211_X1 _10017_ ( .A(_02300_ ), .B(fanout_net_22 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02301_ ) );
NAND3_X1 _10018_ ( .A1(_02299_ ), .A2(_02301_ ), .A3(_01771_ ), .ZN(_02302_ ) );
MUX2_X1 _10019_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02303_ ) );
MUX2_X1 _10020_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02304_ ) );
MUX2_X1 _10021_ ( .A(_02303_ ), .B(_02304_ ), .S(_01777_ ), .Z(_02305_ ) );
OAI211_X1 _10022_ ( .A(_01713_ ), .B(_02302_ ), .C1(_02305_ ), .C2(_01779_ ), .ZN(_02306_ ) );
OAI211_X1 _10023_ ( .A(_02297_ ), .B(_02306_ ), .C1(_01759_ ), .C2(_01790_ ), .ZN(_02307_ ) );
OR3_X2 _10024_ ( .A1(_01761_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01758_ ), .ZN(_02308_ ) );
NAND2_X2 _10025_ ( .A1(_02307_ ), .A2(_02308_ ), .ZN(_02309_ ) );
INV_X1 _10026_ ( .A(\ID_EX_imm [15] ), .ZN(_02310_ ) );
XNOR2_X1 _10027_ ( .A(_02309_ ), .B(_02310_ ), .ZN(_02311_ ) );
OR2_X1 _10028_ ( .A1(_01823_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02312_ ) );
OAI211_X1 _10029_ ( .A(_02312_ ), .B(_01834_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02313_ ) );
OR2_X1 _10030_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02314_ ) );
OAI211_X1 _10031_ ( .A(_02314_ ), .B(fanout_net_22 ), .C1(_01846_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02315_ ) );
NAND3_X1 _10032_ ( .A1(_02313_ ), .A2(_01771_ ), .A3(_02315_ ), .ZN(_02316_ ) );
MUX2_X1 _10033_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02317_ ) );
MUX2_X1 _10034_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02318_ ) );
MUX2_X1 _10035_ ( .A(_02317_ ), .B(_02318_ ), .S(_01696_ ), .Z(_02319_ ) );
OAI211_X1 _10036_ ( .A(_01713_ ), .B(_02316_ ), .C1(_02319_ ), .C2(_01721_ ), .ZN(_02320_ ) );
OR2_X1 _10037_ ( .A1(_01823_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02321_ ) );
OAI211_X1 _10038_ ( .A(_02321_ ), .B(fanout_net_22 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02322_ ) );
OR2_X1 _10039_ ( .A1(_01823_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02323_ ) );
OAI211_X1 _10040_ ( .A(_02323_ ), .B(_01834_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02324_ ) );
NAND3_X1 _10041_ ( .A1(_02322_ ), .A2(_02324_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02325_ ) );
MUX2_X1 _10042_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02326_ ) );
MUX2_X1 _10043_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02327_ ) );
MUX2_X1 _10044_ ( .A(_02326_ ), .B(_02327_ ), .S(fanout_net_22 ), .Z(_02328_ ) );
OAI211_X1 _10045_ ( .A(fanout_net_24 ), .B(_02325_ ), .C1(_02328_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02329_ ) );
OAI211_X1 _10046_ ( .A(_02320_ ), .B(_02329_ ), .C1(_01730_ ), .C2(_01790_ ), .ZN(_02330_ ) );
OR3_X4 _10047_ ( .A1(_01761_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01729_ ), .ZN(_02331_ ) );
NAND2_X2 _10048_ ( .A1(_02330_ ), .A2(_02331_ ), .ZN(_02332_ ) );
INV_X1 _10049_ ( .A(\ID_EX_imm [14] ), .ZN(_02333_ ) );
XNOR2_X1 _10050_ ( .A(_02332_ ), .B(_02333_ ), .ZN(_02334_ ) );
AND2_X1 _10051_ ( .A1(_02311_ ), .A2(_02334_ ), .ZN(_02335_ ) );
OR2_X1 _10052_ ( .A1(_01698_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02336_ ) );
OAI211_X1 _10053_ ( .A(_02336_ ), .B(_01777_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02337_ ) );
OR2_X1 _10054_ ( .A1(_01698_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02338_ ) );
OAI211_X1 _10055_ ( .A(_02338_ ), .B(fanout_net_22 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02339_ ) );
NAND3_X1 _10056_ ( .A1(_02337_ ), .A2(_02339_ ), .A3(_01720_ ), .ZN(_02340_ ) );
MUX2_X1 _10057_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02341_ ) );
MUX2_X1 _10058_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02342_ ) );
MUX2_X1 _10059_ ( .A(_02341_ ), .B(_02342_ ), .S(_01777_ ), .Z(_02343_ ) );
OAI211_X1 _10060_ ( .A(_01712_ ), .B(_02340_ ), .C1(_02343_ ), .C2(_01771_ ), .ZN(_02344_ ) );
OR2_X1 _10061_ ( .A1(_01698_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02345_ ) );
OAI211_X1 _10062_ ( .A(_02345_ ), .B(fanout_net_22 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02346_ ) );
OR2_X1 _10063_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02347_ ) );
OAI211_X1 _10064_ ( .A(_02347_ ), .B(_01777_ ), .C1(_01688_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02348_ ) );
NAND3_X1 _10065_ ( .A1(_02346_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02348_ ), .ZN(_02349_ ) );
MUX2_X1 _10066_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02350_ ) );
MUX2_X1 _10067_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02351_ ) );
MUX2_X1 _10068_ ( .A(_02350_ ), .B(_02351_ ), .S(fanout_net_22 ), .Z(_02352_ ) );
OAI211_X1 _10069_ ( .A(fanout_net_24 ), .B(_02349_ ), .C1(_02352_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02353_ ) );
OAI211_X1 _10070_ ( .A(_02344_ ), .B(_02353_ ), .C1(_01759_ ), .C2(_01761_ ), .ZN(_02354_ ) );
INV_X1 _10071_ ( .A(\ID_EX_imm [13] ), .ZN(_02355_ ) );
OR3_X1 _10072_ ( .A1(_01726_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01758_ ), .ZN(_02356_ ) );
AND3_X1 _10073_ ( .A1(_02354_ ), .A2(_02355_ ), .A3(_02356_ ), .ZN(_02357_ ) );
AOI21_X1 _10074_ ( .A(_02355_ ), .B1(_02354_ ), .B2(_02356_ ), .ZN(_02358_ ) );
NOR2_X1 _10075_ ( .A1(_02357_ ), .A2(_02358_ ), .ZN(_02359_ ) );
NOR2_X1 _10076_ ( .A1(_01688_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02360_ ) );
OAI21_X1 _10077_ ( .A(fanout_net_22 ), .B1(fanout_net_18 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02361_ ) );
NOR2_X1 _10078_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02362_ ) );
OAI21_X1 _10079_ ( .A(_01777_ ), .B1(_01699_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02363_ ) );
OAI221_X1 _10080_ ( .A(_01720_ ), .B1(_02360_ ), .B2(_02361_ ), .C1(_02362_ ), .C2(_02363_ ), .ZN(_02364_ ) );
MUX2_X1 _10081_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02365_ ) );
MUX2_X1 _10082_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02366_ ) );
MUX2_X1 _10083_ ( .A(_02365_ ), .B(_02366_ ), .S(fanout_net_22 ), .Z(_02367_ ) );
OAI211_X1 _10084_ ( .A(fanout_net_24 ), .B(_02364_ ), .C1(_02367_ ), .C2(_01779_ ), .ZN(_02368_ ) );
OR2_X1 _10085_ ( .A1(_01767_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02369_ ) );
OAI211_X1 _10086_ ( .A(_02369_ ), .B(fanout_net_22 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02370_ ) );
OR2_X1 _10087_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02371_ ) );
OAI211_X1 _10088_ ( .A(_02371_ ), .B(_01696_ ), .C1(_01699_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02372_ ) );
NAND3_X1 _10089_ ( .A1(_02370_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02372_ ), .ZN(_02373_ ) );
MUX2_X1 _10090_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02374_ ) );
MUX2_X1 _10091_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02375_ ) );
MUX2_X1 _10092_ ( .A(_02374_ ), .B(_02375_ ), .S(_01777_ ), .Z(_02376_ ) );
OAI211_X1 _10093_ ( .A(_01713_ ), .B(_02373_ ), .C1(_02376_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02377_ ) );
OAI211_X1 _10094_ ( .A(_02368_ ), .B(_02377_ ), .C1(_01759_ ), .C2(_01790_ ), .ZN(_02378_ ) );
OR3_X1 _10095_ ( .A1(_01761_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01729_ ), .ZN(_02379_ ) );
NAND2_X2 _10096_ ( .A1(_02378_ ), .A2(_02379_ ), .ZN(_02380_ ) );
INV_X1 _10097_ ( .A(\ID_EX_imm [12] ), .ZN(_02381_ ) );
XNOR2_X1 _10098_ ( .A(_02380_ ), .B(_02381_ ), .ZN(_02382_ ) );
NAND3_X1 _10099_ ( .A1(_02335_ ), .A2(_02359_ ), .A3(_02382_ ), .ZN(_02383_ ) );
OR2_X4 _10100_ ( .A1(_02288_ ), .A2(_02383_ ), .ZN(_02384_ ) );
NAND2_X1 _10101_ ( .A1(_02380_ ), .A2(\ID_EX_imm [12] ), .ZN(_02385_ ) );
NOR3_X1 _10102_ ( .A1(_02385_ ), .A2(_02357_ ), .A3(_02358_ ), .ZN(_02386_ ) );
OAI211_X1 _10103_ ( .A(_02311_ ), .B(_02334_ ), .C1(_02386_ ), .C2(_02358_ ), .ZN(_02387_ ) );
NAND2_X1 _10104_ ( .A1(_02309_ ), .A2(\ID_EX_imm [15] ), .ZN(_02388_ ) );
NAND3_X1 _10105_ ( .A1(_02311_ ), .A2(\ID_EX_imm [14] ), .A3(_02332_ ), .ZN(_02389_ ) );
AND3_X1 _10106_ ( .A1(_02387_ ), .A2(_02388_ ), .A3(_02389_ ), .ZN(_02390_ ) );
AOI211_X2 _10107_ ( .A(_01874_ ), .B(_01968_ ), .C1(_02384_ ), .C2(_02390_ ), .ZN(_02391_ ) );
AND2_X1 _10108_ ( .A1(_01965_ ), .A2(\ID_EX_imm [16] ), .ZN(_02392_ ) );
AND2_X1 _10109_ ( .A1(_01944_ ), .A2(_02392_ ), .ZN(_02393_ ) );
AOI21_X1 _10110_ ( .A(_02393_ ), .B1(\ID_EX_imm [17] ), .B2(_01942_ ), .ZN(_02394_ ) );
INV_X1 _10111_ ( .A(_02394_ ), .ZN(_02395_ ) );
NAND2_X1 _10112_ ( .A1(_02395_ ), .A2(_01921_ ), .ZN(_02396_ ) );
AND2_X1 _10113_ ( .A1(_01895_ ), .A2(\ID_EX_imm [18] ), .ZN(_02397_ ) );
AND2_X1 _10114_ ( .A1(_01920_ ), .A2(_02397_ ), .ZN(_02398_ ) );
AOI21_X1 _10115_ ( .A(_02398_ ), .B1(\ID_EX_imm [19] ), .B2(_01918_ ), .ZN(_02399_ ) );
AND2_X1 _10116_ ( .A1(_02396_ ), .A2(_02399_ ), .ZN(_02400_ ) );
OR2_X1 _10117_ ( .A1(_02400_ ), .A2(_01874_ ), .ZN(_02401_ ) );
OAI211_X1 _10118_ ( .A(\ID_EX_imm [20] ), .B(_01869_ ), .C1(_01843_ ), .C2(\ID_EX_imm [21] ), .ZN(_02402_ ) );
INV_X2 _10119_ ( .A(_01843_ ), .ZN(_02403_ ) );
OAI21_X1 _10120_ ( .A(_02402_ ), .B1(_01844_ ), .B2(_02403_ ), .ZN(_02404_ ) );
NAND2_X1 _10121_ ( .A1(_01819_ ), .A2(_02404_ ), .ZN(_02405_ ) );
AND2_X1 _10122_ ( .A1(_01793_ ), .A2(\ID_EX_imm [22] ), .ZN(_02406_ ) );
NAND3_X1 _10123_ ( .A1(_02406_ ), .A2(_01817_ ), .A3(_01818_ ), .ZN(_02407_ ) );
NAND4_X1 _10124_ ( .A1(_02401_ ), .A2(_01818_ ), .A3(_02405_ ), .A4(_02407_ ), .ZN(_02408_ ) );
OR2_X2 _10125_ ( .A1(_02391_ ), .A2(_02408_ ), .ZN(_02409_ ) );
OR2_X1 _10126_ ( .A1(_01689_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02410_ ) );
OAI211_X1 _10127_ ( .A(_02410_ ), .B(_01739_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02411_ ) );
INV_X1 _10128_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02412_ ) );
NAND2_X1 _10129_ ( .A1(_02412_ ), .A2(fanout_net_19 ), .ZN(_02413_ ) );
OAI211_X1 _10130_ ( .A(_02413_ ), .B(fanout_net_22 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02414_ ) );
NAND3_X1 _10131_ ( .A1(_02411_ ), .A2(_02414_ ), .A3(_01722_ ), .ZN(_02415_ ) );
MUX2_X1 _10132_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02416_ ) );
MUX2_X1 _10133_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02417_ ) );
MUX2_X1 _10134_ ( .A(_02416_ ), .B(_02417_ ), .S(_01739_ ), .Z(_02418_ ) );
OAI211_X1 _10135_ ( .A(fanout_net_24 ), .B(_02415_ ), .C1(_02418_ ), .C2(_01747_ ), .ZN(_02419_ ) );
OR2_X1 _10136_ ( .A1(_01689_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02420_ ) );
OAI211_X1 _10137_ ( .A(_02420_ ), .B(_01739_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02421_ ) );
INV_X1 _10138_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02422_ ) );
NAND2_X1 _10139_ ( .A1(_02422_ ), .A2(fanout_net_19 ), .ZN(_02423_ ) );
OAI211_X1 _10140_ ( .A(_02423_ ), .B(fanout_net_22 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02424_ ) );
NAND3_X1 _10141_ ( .A1(_02421_ ), .A2(_02424_ ), .A3(_01722_ ), .ZN(_02425_ ) );
MUX2_X1 _10142_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02426_ ) );
MUX2_X1 _10143_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02427_ ) );
MUX2_X1 _10144_ ( .A(_02426_ ), .B(_02427_ ), .S(_01848_ ), .Z(_02428_ ) );
OAI211_X1 _10145_ ( .A(_01714_ ), .B(_02425_ ), .C1(_02428_ ), .C2(_01747_ ), .ZN(_02429_ ) );
OAI211_X1 _10146_ ( .A(_02419_ ), .B(_02429_ ), .C1(_01760_ ), .C2(_01762_ ), .ZN(_02430_ ) );
OR3_X1 _10147_ ( .A1(_01762_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01730_ ), .ZN(_02431_ ) );
NAND2_X2 _10148_ ( .A1(_02430_ ), .A2(_02431_ ), .ZN(_02432_ ) );
INV_X1 _10149_ ( .A(\ID_EX_imm [24] ), .ZN(_02433_ ) );
XNOR2_X1 _10150_ ( .A(_02432_ ), .B(_02433_ ), .ZN(_02434_ ) );
OR2_X1 _10151_ ( .A1(_01823_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02435_ ) );
OAI211_X1 _10152_ ( .A(_02435_ ), .B(_01834_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02436_ ) );
INV_X1 _10153_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02437_ ) );
NAND2_X1 _10154_ ( .A1(_02437_ ), .A2(fanout_net_19 ), .ZN(_02438_ ) );
OAI211_X1 _10155_ ( .A(_02438_ ), .B(fanout_net_22 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02439_ ) );
NAND3_X1 _10156_ ( .A1(_02436_ ), .A2(_02439_ ), .A3(_01779_ ), .ZN(_02440_ ) );
MUX2_X1 _10157_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02441_ ) );
MUX2_X1 _10158_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02442_ ) );
MUX2_X1 _10159_ ( .A(_02441_ ), .B(_02442_ ), .S(_01696_ ), .Z(_02443_ ) );
OAI211_X1 _10160_ ( .A(_01713_ ), .B(_02440_ ), .C1(_02443_ ), .C2(_01721_ ), .ZN(_02444_ ) );
OR2_X1 _10161_ ( .A1(_01823_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02445_ ) );
OAI211_X1 _10162_ ( .A(_02445_ ), .B(fanout_net_22 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02446_ ) );
OR2_X1 _10163_ ( .A1(_01823_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02447_ ) );
OAI211_X1 _10164_ ( .A(_02447_ ), .B(_01834_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02448_ ) );
NAND3_X1 _10165_ ( .A1(_02446_ ), .A2(_02448_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02449_ ) );
MUX2_X1 _10166_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02450_ ) );
MUX2_X1 _10167_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02451_ ) );
MUX2_X1 _10168_ ( .A(_02450_ ), .B(_02451_ ), .S(fanout_net_22 ), .Z(_02452_ ) );
OAI211_X1 _10169_ ( .A(fanout_net_24 ), .B(_02449_ ), .C1(_02452_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02453_ ) );
OAI211_X1 _10170_ ( .A(_02444_ ), .B(_02453_ ), .C1(_01730_ ), .C2(_01790_ ), .ZN(_02454_ ) );
OR3_X1 _10171_ ( .A1(_01761_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01729_ ), .ZN(_02455_ ) );
NAND2_X2 _10172_ ( .A1(_02454_ ), .A2(_02455_ ), .ZN(_02456_ ) );
INV_X1 _10173_ ( .A(\ID_EX_imm [25] ), .ZN(_02457_ ) );
XNOR2_X1 _10174_ ( .A(_02456_ ), .B(_02457_ ), .ZN(_02458_ ) );
AND3_X4 _10175_ ( .A1(_02409_ ), .A2(_02434_ ), .A3(_02458_ ), .ZN(_02459_ ) );
INV_X2 _10176_ ( .A(_02459_ ), .ZN(_02460_ ) );
AND2_X1 _10177_ ( .A1(_02432_ ), .A2(\ID_EX_imm [24] ), .ZN(_02461_ ) );
AND2_X1 _10178_ ( .A1(_02458_ ), .A2(_02461_ ), .ZN(_02462_ ) );
AOI21_X1 _10179_ ( .A(_02462_ ), .B1(\ID_EX_imm [25] ), .B2(_02456_ ), .ZN(_02463_ ) );
NAND2_X2 _10180_ ( .A1(_02460_ ), .A2(_02463_ ), .ZN(_02464_ ) );
OR2_X1 _10181_ ( .A1(_01699_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02465_ ) );
OAI211_X1 _10182_ ( .A(_02465_ ), .B(fanout_net_22 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02466_ ) );
OR2_X1 _10183_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02467_ ) );
OAI211_X1 _10184_ ( .A(_02467_ ), .B(_01697_ ), .C1(_01700_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02468_ ) );
NAND3_X1 _10185_ ( .A1(_02466_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02468_ ), .ZN(_02469_ ) );
MUX2_X1 _10186_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02470_ ) );
MUX2_X1 _10187_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02471_ ) );
MUX2_X1 _10188_ ( .A(_02470_ ), .B(_02471_ ), .S(_01697_ ), .Z(_02472_ ) );
OAI211_X1 _10189_ ( .A(_01714_ ), .B(_02469_ ), .C1(_02472_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02473_ ) );
NOR2_X1 _10190_ ( .A1(_01689_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02474_ ) );
OAI21_X1 _10191_ ( .A(fanout_net_22 ), .B1(fanout_net_19 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02475_ ) );
INV_X1 _10192_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02476_ ) );
INV_X1 _10193_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02477_ ) );
MUX2_X1 _10194_ ( .A(_02476_ ), .B(_02477_ ), .S(fanout_net_19 ), .Z(_02478_ ) );
OAI221_X1 _10195_ ( .A(_01721_ ), .B1(_02474_ ), .B2(_02475_ ), .C1(_02478_ ), .C2(fanout_net_22 ), .ZN(_02479_ ) );
MUX2_X1 _10196_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02480_ ) );
MUX2_X1 _10197_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02481_ ) );
MUX2_X1 _10198_ ( .A(_02480_ ), .B(_02481_ ), .S(fanout_net_22 ), .Z(_02482_ ) );
OAI211_X1 _10199_ ( .A(fanout_net_24 ), .B(_02479_ ), .C1(_02482_ ), .C2(_01722_ ), .ZN(_02483_ ) );
OAI211_X1 _10200_ ( .A(_02473_ ), .B(_02483_ ), .C1(_01760_ ), .C2(_01762_ ), .ZN(_02484_ ) );
INV_X1 _10201_ ( .A(\ID_EX_imm [27] ), .ZN(_02485_ ) );
OR3_X1 _10202_ ( .A1(_01727_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01759_ ), .ZN(_02486_ ) );
AND3_X1 _10203_ ( .A1(_02484_ ), .A2(_02485_ ), .A3(_02486_ ), .ZN(_02487_ ) );
AOI21_X1 _10204_ ( .A(_02485_ ), .B1(_02484_ ), .B2(_02486_ ), .ZN(_02488_ ) );
NOR2_X1 _10205_ ( .A1(_02487_ ), .A2(_02488_ ), .ZN(_02489_ ) );
OR2_X1 _10206_ ( .A1(_01699_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02490_ ) );
OAI211_X1 _10207_ ( .A(_02490_ ), .B(_01697_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02491_ ) );
OR2_X1 _10208_ ( .A1(_01688_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02492_ ) );
OAI211_X1 _10209_ ( .A(_02492_ ), .B(fanout_net_22 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02493_ ) );
NAND3_X1 _10210_ ( .A1(_02491_ ), .A2(_02493_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02494_ ) );
MUX2_X1 _10211_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02495_ ) );
MUX2_X1 _10212_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02496_ ) );
MUX2_X1 _10213_ ( .A(_02495_ ), .B(_02496_ ), .S(_01738_ ), .Z(_02497_ ) );
OAI211_X1 _10214_ ( .A(_01714_ ), .B(_02494_ ), .C1(_02497_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02498_ ) );
NOR2_X1 _10215_ ( .A1(_01846_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02499_ ) );
OAI21_X1 _10216_ ( .A(fanout_net_22 ), .B1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02500_ ) );
NOR2_X1 _10217_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02501_ ) );
OAI21_X1 _10218_ ( .A(_01738_ ), .B1(_01689_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02502_ ) );
OAI221_X1 _10219_ ( .A(_01779_ ), .B1(_02499_ ), .B2(_02500_ ), .C1(_02501_ ), .C2(_02502_ ), .ZN(_02503_ ) );
MUX2_X1 _10220_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02504_ ) );
MUX2_X1 _10221_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02505_ ) );
MUX2_X1 _10222_ ( .A(_02504_ ), .B(_02505_ ), .S(fanout_net_22 ), .Z(_02506_ ) );
OAI211_X1 _10223_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02503_ ), .C1(_02506_ ), .C2(_01850_ ), .ZN(_02507_ ) );
OAI211_X1 _10224_ ( .A(_02498_ ), .B(_02507_ ), .C1(_01760_ ), .C2(_01727_ ), .ZN(_02508_ ) );
OR3_X1 _10225_ ( .A1(_01790_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01759_ ), .ZN(_02509_ ) );
NAND2_X2 _10226_ ( .A1(_02508_ ), .A2(_02509_ ), .ZN(_02510_ ) );
INV_X1 _10227_ ( .A(\ID_EX_imm [26] ), .ZN(_02511_ ) );
XNOR2_X1 _10228_ ( .A(_02510_ ), .B(_02511_ ), .ZN(_02512_ ) );
NAND3_X2 _10229_ ( .A1(_02464_ ), .A2(_02489_ ), .A3(_02512_ ), .ZN(_02513_ ) );
INV_X1 _10230_ ( .A(_02510_ ), .ZN(_02514_ ) );
NOR4_X1 _10231_ ( .A1(_02487_ ), .A2(_02514_ ), .A3(_02488_ ), .A4(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02515_ ) );
NOR2_X1 _10232_ ( .A1(_02515_ ), .A2(_02488_ ), .ZN(_02516_ ) );
AOI21_X2 _10233_ ( .A(_01766_ ), .B1(_02513_ ), .B2(_02516_ ), .ZN(_02517_ ) );
OR2_X1 _10234_ ( .A1(_01700_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02518_ ) );
OAI211_X1 _10235_ ( .A(_02518_ ), .B(fanout_net_22 ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02519_ ) );
INV_X1 _10236_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02520_ ) );
INV_X1 _10237_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02521_ ) );
MUX2_X1 _10238_ ( .A(_02520_ ), .B(_02521_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02522_ ) );
OAI211_X1 _10239_ ( .A(_02519_ ), .B(_01747_ ), .C1(_02522_ ), .C2(fanout_net_22 ), .ZN(_02523_ ) );
MUX2_X1 _10240_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02524_ ) );
MUX2_X1 _10241_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02525_ ) );
MUX2_X1 _10242_ ( .A(_02524_ ), .B(_02525_ ), .S(_01739_ ), .Z(_02526_ ) );
OAI211_X1 _10243_ ( .A(_02523_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .C1(_02526_ ), .C2(_01747_ ), .ZN(_02527_ ) );
OR2_X1 _10244_ ( .A1(_01700_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02528_ ) );
OAI211_X1 _10245_ ( .A(_02528_ ), .B(_01739_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02529_ ) );
OR2_X1 _10246_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02530_ ) );
OAI211_X1 _10247_ ( .A(_02530_ ), .B(fanout_net_22 ), .C1(_01700_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02531_ ) );
NAND3_X1 _10248_ ( .A1(_02529_ ), .A2(_02531_ ), .A3(_01747_ ), .ZN(_02532_ ) );
MUX2_X1 _10249_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02533_ ) );
MUX2_X1 _10250_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02534_ ) );
MUX2_X1 _10251_ ( .A(_02533_ ), .B(_02534_ ), .S(_01739_ ), .Z(_02535_ ) );
OAI211_X1 _10252_ ( .A(_01714_ ), .B(_02532_ ), .C1(_02535_ ), .C2(_01747_ ), .ZN(_02536_ ) );
OAI211_X1 _10253_ ( .A(_02527_ ), .B(_02536_ ), .C1(_01760_ ), .C2(_01762_ ), .ZN(_02537_ ) );
OR3_X1 _10254_ ( .A1(_01762_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01760_ ), .ZN(_02538_ ) );
NAND2_X2 _10255_ ( .A1(_02537_ ), .A2(_02538_ ), .ZN(_02539_ ) );
INV_X1 _10256_ ( .A(\ID_EX_imm [29] ), .ZN(_02540_ ) );
XNOR2_X1 _10257_ ( .A(_02539_ ), .B(_02540_ ), .ZN(_02541_ ) );
NAND2_X2 _10258_ ( .A1(_02517_ ), .A2(_02541_ ), .ZN(_02542_ ) );
AOI21_X1 _10259_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_01763_ ), .B2(_01764_ ), .ZN(_02543_ ) );
INV_X1 _10260_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02544_ ) );
AOI22_X1 _10261_ ( .A1(_02541_ ), .A2(_02543_ ), .B1(_02544_ ), .B2(_02539_ ), .ZN(_02545_ ) );
AOI21_X1 _10262_ ( .A(_01734_ ), .B1(_02542_ ), .B2(_02545_ ), .ZN(_02546_ ) );
AOI21_X1 _10263_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_01724_ ), .B2(_01731_ ), .ZN(_02547_ ) );
NOR2_X1 _10264_ ( .A1(_02546_ ), .A2(_02547_ ), .ZN(_02548_ ) );
OR2_X1 _10265_ ( .A1(_01846_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02549_ ) );
OAI211_X1 _10266_ ( .A(_02549_ ), .B(fanout_net_22 ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02550_ ) );
INV_X1 _10267_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02551_ ) );
INV_X1 _10268_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02552_ ) );
MUX2_X1 _10269_ ( .A(_02551_ ), .B(_02552_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02553_ ) );
OAI211_X1 _10270_ ( .A(_02550_ ), .B(_01850_ ), .C1(_02553_ ), .C2(fanout_net_22 ), .ZN(_02554_ ) );
MUX2_X1 _10271_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02555_ ) );
MUX2_X1 _10272_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02556_ ) );
MUX2_X1 _10273_ ( .A(_02555_ ), .B(_02556_ ), .S(_01848_ ), .Z(_02557_ ) );
OAI211_X1 _10274_ ( .A(_02554_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .C1(_02557_ ), .C2(_01747_ ), .ZN(_02558_ ) );
OR2_X1 _10275_ ( .A1(_01846_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02559_ ) );
OAI211_X1 _10276_ ( .A(_02559_ ), .B(_01848_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02560_ ) );
OR2_X1 _10277_ ( .A1(_01846_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02561_ ) );
OAI211_X1 _10278_ ( .A(_02561_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02562_ ) );
NAND3_X1 _10279_ ( .A1(_02560_ ), .A2(_02562_ ), .A3(_01850_ ), .ZN(_02563_ ) );
MUX2_X1 _10280_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02564_ ) );
MUX2_X1 _10281_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02565_ ) );
MUX2_X1 _10282_ ( .A(_02564_ ), .B(_02565_ ), .S(_01848_ ), .Z(_02566_ ) );
OAI211_X1 _10283_ ( .A(_01714_ ), .B(_02563_ ), .C1(_02566_ ), .C2(_01747_ ), .ZN(_02567_ ) );
NAND2_X1 _10284_ ( .A1(_02558_ ), .A2(_02567_ ), .ZN(_02568_ ) );
NAND2_X1 _10285_ ( .A1(_02568_ ), .A2(_01683_ ), .ZN(_02569_ ) );
NAND4_X1 _10286_ ( .A1(_02037_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01671_ ), .A4(_01666_ ), .ZN(_02570_ ) );
AND2_X2 _10287_ ( .A1(_02569_ ), .A2(_02570_ ), .ZN(_02571_ ) );
XNOR2_X1 _10288_ ( .A(_02571_ ), .B(\ID_EX_imm [31] ), .ZN(_02572_ ) );
XNOR2_X1 _10289_ ( .A(_02548_ ), .B(_02572_ ), .ZN(_02573_ ) );
NOR2_X1 _10290_ ( .A1(_01659_ ), .A2(\ID_EX_typ [5] ), .ZN(_02574_ ) );
AND2_X1 _10291_ ( .A1(_02574_ ), .A2(\ID_EX_typ [7] ), .ZN(_02575_ ) );
BUF_X4 _10292_ ( .A(_02575_ ), .Z(_02576_ ) );
AND2_X1 _10293_ ( .A1(_01646_ ), .A2(\ID_EX_typ [7] ), .ZN(_02577_ ) );
BUF_X4 _10294_ ( .A(_02577_ ), .Z(_02578_ ) );
NOR2_X1 _10295_ ( .A1(_02576_ ), .A2(_02578_ ), .ZN(_02579_ ) );
INV_X1 _10296_ ( .A(_02579_ ), .ZN(_02580_ ) );
BUF_X4 _10297_ ( .A(_02580_ ), .Z(_02581_ ) );
NOR2_X1 _10298_ ( .A1(_02573_ ), .A2(_02581_ ), .ZN(_00095_ ) );
NAND2_X1 _10299_ ( .A1(_02542_ ), .A2(_02545_ ), .ZN(_02582_ ) );
XNOR2_X1 _10300_ ( .A(_02582_ ), .B(_01734_ ), .ZN(_02583_ ) );
CLKBUF_X2 _10301_ ( .A(_02579_ ), .Z(_02584_ ) );
AND2_X1 _10302_ ( .A1(_02583_ ), .A2(_02584_ ), .ZN(_00096_ ) );
AOI21_X1 _10303_ ( .A(_01968_ ), .B1(_02384_ ), .B2(_02390_ ), .ZN(_02585_ ) );
INV_X1 _10304_ ( .A(_02400_ ), .ZN(_02586_ ) );
OAI21_X1 _10305_ ( .A(_01871_ ), .B1(_02585_ ), .B2(_02586_ ), .ZN(_02587_ ) );
NAND2_X1 _10306_ ( .A1(_01869_ ), .A2(\ID_EX_imm [20] ), .ZN(_02588_ ) );
AND2_X1 _10307_ ( .A1(_02587_ ), .A2(_02588_ ), .ZN(_02589_ ) );
XNOR2_X1 _10308_ ( .A(_02589_ ), .B(_01845_ ), .ZN(_02590_ ) );
AND2_X1 _10309_ ( .A1(_02590_ ), .A2(_02584_ ), .ZN(_00097_ ) );
NOR2_X1 _10310_ ( .A1(_02585_ ), .A2(_02586_ ), .ZN(_02591_ ) );
XNOR2_X1 _10311_ ( .A(_02591_ ), .B(_01871_ ), .ZN(_02592_ ) );
AND2_X1 _10312_ ( .A1(_02592_ ), .A2(_02584_ ), .ZN(_00098_ ) );
INV_X1 _10313_ ( .A(_01967_ ), .ZN(_02593_ ) );
AOI21_X1 _10314_ ( .A(_02593_ ), .B1(_02384_ ), .B2(_02390_ ), .ZN(_02594_ ) );
AND2_X1 _10315_ ( .A1(_02594_ ), .A2(_01944_ ), .ZN(_02595_ ) );
OAI21_X1 _10316_ ( .A(_01897_ ), .B1(_02595_ ), .B2(_02395_ ), .ZN(_02596_ ) );
INV_X1 _10317_ ( .A(_02397_ ), .ZN(_02597_ ) );
NAND2_X1 _10318_ ( .A1(_02596_ ), .A2(_02597_ ), .ZN(_02598_ ) );
XNOR2_X1 _10319_ ( .A(_02598_ ), .B(_01920_ ), .ZN(_02599_ ) );
NOR2_X1 _10320_ ( .A1(_02599_ ), .A2(_02581_ ), .ZN(_00099_ ) );
NOR2_X1 _10321_ ( .A1(_02595_ ), .A2(_02395_ ), .ZN(_02600_ ) );
XNOR2_X1 _10322_ ( .A(_02600_ ), .B(_01897_ ), .ZN(_02601_ ) );
AND2_X1 _10323_ ( .A1(_02601_ ), .A2(_02584_ ), .ZN(_00100_ ) );
OR2_X1 _10324_ ( .A1(_02594_ ), .A2(_02392_ ), .ZN(_02602_ ) );
XNOR2_X1 _10325_ ( .A(_02602_ ), .B(_01944_ ), .ZN(_02603_ ) );
NOR2_X1 _10326_ ( .A1(_02603_ ), .A2(_02581_ ), .ZN(_00101_ ) );
AND3_X1 _10327_ ( .A1(_02384_ ), .A2(_02390_ ), .A3(_02593_ ), .ZN(_02604_ ) );
NOR3_X1 _10328_ ( .A1(_02604_ ), .A2(_02594_ ), .A3(_02580_ ), .ZN(_00102_ ) );
INV_X1 _10329_ ( .A(_02382_ ), .ZN(_02605_ ) );
NOR4_X1 _10330_ ( .A1(_02288_ ), .A2(_02357_ ), .A3(_02358_ ), .A4(_02605_ ), .ZN(_02606_ ) );
OR2_X1 _10331_ ( .A1(_02386_ ), .A2(_02358_ ), .ZN(_02607_ ) );
OAI21_X1 _10332_ ( .A(_02334_ ), .B1(_02606_ ), .B2(_02607_ ), .ZN(_02608_ ) );
NAND2_X1 _10333_ ( .A1(_02332_ ), .A2(\ID_EX_imm [14] ), .ZN(_02609_ ) );
NAND2_X1 _10334_ ( .A1(_02608_ ), .A2(_02609_ ), .ZN(_02610_ ) );
XNOR2_X1 _10335_ ( .A(_02610_ ), .B(_02311_ ), .ZN(_02611_ ) );
NOR2_X1 _10336_ ( .A1(_02611_ ), .A2(_02581_ ), .ZN(_00103_ ) );
OR3_X1 _10337_ ( .A1(_02606_ ), .A2(_02334_ ), .A3(_02607_ ), .ZN(_02612_ ) );
AND3_X1 _10338_ ( .A1(_02612_ ), .A2(_02579_ ), .A3(_02608_ ), .ZN(_00104_ ) );
OAI21_X1 _10339_ ( .A(_02382_ ), .B1(_02278_ ), .B2(_02287_ ), .ZN(_02613_ ) );
NAND2_X1 _10340_ ( .A1(_02613_ ), .A2(_02385_ ), .ZN(_02614_ ) );
XNOR2_X1 _10341_ ( .A(_02614_ ), .B(_02359_ ), .ZN(_02615_ ) );
NOR2_X1 _10342_ ( .A1(_02615_ ), .A2(_02581_ ), .ZN(_00105_ ) );
XNOR2_X1 _10343_ ( .A(_02288_ ), .B(_02382_ ), .ZN(_02616_ ) );
AND2_X1 _10344_ ( .A1(_02616_ ), .A2(_02584_ ), .ZN(_00106_ ) );
OR2_X1 _10345_ ( .A1(_02517_ ), .A2(_02543_ ), .ZN(_02617_ ) );
XNOR2_X1 _10346_ ( .A(_02617_ ), .B(_02541_ ), .ZN(_02618_ ) );
NOR2_X1 _10347_ ( .A1(_02618_ ), .A2(_02581_ ), .ZN(_00107_ ) );
AND3_X1 _10348_ ( .A1(_02513_ ), .A2(_02516_ ), .A3(_01766_ ), .ZN(_02619_ ) );
NOR3_X1 _10349_ ( .A1(_02619_ ), .A2(_02517_ ), .A3(_02580_ ), .ZN(_00108_ ) );
NAND2_X1 _10350_ ( .A1(_02464_ ), .A2(_02512_ ), .ZN(_02620_ ) );
OR2_X1 _10351_ ( .A1(_02514_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02621_ ) );
NAND2_X1 _10352_ ( .A1(_02620_ ), .A2(_02621_ ), .ZN(_02622_ ) );
XNOR2_X1 _10353_ ( .A(_02622_ ), .B(_02489_ ), .ZN(_02623_ ) );
NOR2_X1 _10354_ ( .A1(_02623_ ), .A2(_02581_ ), .ZN(_00109_ ) );
XOR2_X1 _10355_ ( .A(_02464_ ), .B(_02512_ ), .Z(_02624_ ) );
AND2_X1 _10356_ ( .A1(_02624_ ), .A2(_02584_ ), .ZN(_00110_ ) );
AND2_X1 _10357_ ( .A1(_02409_ ), .A2(_02434_ ), .ZN(_02625_ ) );
NOR2_X1 _10358_ ( .A1(_02625_ ), .A2(_02461_ ), .ZN(_02626_ ) );
XNOR2_X1 _10359_ ( .A(_02626_ ), .B(_02458_ ), .ZN(_02627_ ) );
AND2_X1 _10360_ ( .A1(_02627_ ), .A2(_02584_ ), .ZN(_00111_ ) );
XOR2_X1 _10361_ ( .A(_02409_ ), .B(_02434_ ), .Z(_02628_ ) );
AND2_X1 _10362_ ( .A1(_02628_ ), .A2(_02584_ ), .ZN(_00112_ ) );
INV_X1 _10363_ ( .A(_01872_ ), .ZN(_02629_ ) );
NOR2_X1 _10364_ ( .A1(_02591_ ), .A2(_02629_ ), .ZN(_02630_ ) );
OAI21_X1 _10365_ ( .A(_01795_ ), .B1(_02630_ ), .B2(_02404_ ), .ZN(_02631_ ) );
INV_X1 _10366_ ( .A(_02406_ ), .ZN(_02632_ ) );
AND4_X1 _10367_ ( .A1(_01817_ ), .A2(_02631_ ), .A3(_01818_ ), .A4(_02632_ ), .ZN(_02633_ ) );
AOI22_X1 _10368_ ( .A1(_02631_ ), .A2(_02632_ ), .B1(_01817_ ), .B2(_01818_ ), .ZN(_02634_ ) );
NOR2_X1 _10369_ ( .A1(_02633_ ), .A2(_02634_ ), .ZN(_02635_ ) );
NOR2_X1 _10370_ ( .A1(_02635_ ), .A2(_02581_ ), .ZN(_00113_ ) );
OR3_X1 _10371_ ( .A1(_02630_ ), .A2(_01795_ ), .A3(_02404_ ), .ZN(_02636_ ) );
AND3_X1 _10372_ ( .A1(_02636_ ), .A2(_02579_ ), .A3(_02631_ ), .ZN(_00114_ ) );
AND2_X1 _10373_ ( .A1(_01329_ ), .A2(\ID_EX_rd [4] ), .ZN(_00115_ ) );
AND2_X1 _10374_ ( .A1(_01329_ ), .A2(\ID_EX_rd [3] ), .ZN(_00116_ ) );
AND2_X1 _10375_ ( .A1(_01329_ ), .A2(\ID_EX_rd [2] ), .ZN(_00117_ ) );
INV_X1 _10376_ ( .A(\ID_EX_rd [1] ), .ZN(_02637_ ) );
NOR2_X1 _10377_ ( .A1(_02637_ ), .A2(fanout_net_2 ), .ZN(_00118_ ) );
AND2_X1 _10378_ ( .A1(_01329_ ), .A2(\ID_EX_rd [0] ), .ZN(_00119_ ) );
BUF_X4 _10379_ ( .A(_02578_ ), .Z(_02638_ ) );
INV_X1 _10380_ ( .A(\EX_LS_dest_csreg_mem [4] ), .ZN(_02639_ ) );
INV_X1 _10381_ ( .A(\ID_EX_csr [8] ), .ZN(_02640_ ) );
AOI22_X1 _10382_ ( .A1(_02639_ ), .A2(\ID_EX_csr [4] ), .B1(_02640_ ), .B2(\EX_LS_dest_csreg_mem [8] ), .ZN(_02641_ ) );
INV_X1 _10383_ ( .A(\ID_EX_csr [1] ), .ZN(_02642_ ) );
OAI221_X1 _10384_ ( .A(_02641_ ), .B1(_02639_ ), .B2(\ID_EX_csr [4] ), .C1(fanout_net_7 ), .C2(_02642_ ), .ZN(_02643_ ) );
INV_X1 _10385_ ( .A(\EX_LS_dest_csreg_mem [11] ), .ZN(_02644_ ) );
INV_X1 _10386_ ( .A(\ID_EX_csr [2] ), .ZN(_02645_ ) );
AOI22_X1 _10387_ ( .A1(_02644_ ), .A2(\ID_EX_csr [11] ), .B1(_02645_ ), .B2(\EX_LS_dest_csreg_mem [2] ), .ZN(_02646_ ) );
INV_X1 _10388_ ( .A(fanout_net_7 ), .ZN(_02647_ ) );
OAI221_X1 _10389_ ( .A(_02646_ ), .B1(\EX_LS_dest_csreg_mem [2] ), .B2(_02645_ ), .C1(_02647_ ), .C2(\ID_EX_csr [1] ), .ZN(_02648_ ) );
XOR2_X1 _10390_ ( .A(\EX_LS_dest_csreg_mem [9] ), .B(\ID_EX_csr [9] ), .Z(_02649_ ) );
INV_X1 _10391_ ( .A(\EX_LS_dest_csreg_mem [10] ), .ZN(_02650_ ) );
OAI22_X1 _10392_ ( .A1(_02650_ ), .A2(\ID_EX_csr [10] ), .B1(_02640_ ), .B2(\EX_LS_dest_csreg_mem [8] ), .ZN(_02651_ ) );
NOR4_X1 _10393_ ( .A1(_02643_ ), .A2(_02648_ ), .A3(_02649_ ), .A4(_02651_ ), .ZN(_02652_ ) );
XNOR2_X1 _10394_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_02653_ ) );
INV_X1 _10395_ ( .A(\EX_LS_dest_csreg_mem [3] ), .ZN(_02654_ ) );
AOI22_X1 _10396_ ( .A1(_02650_ ), .A2(\ID_EX_csr [10] ), .B1(_02654_ ), .B2(\ID_EX_csr [3] ), .ZN(_02655_ ) );
XNOR2_X1 _10397_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_02656_ ) );
INV_X1 _10398_ ( .A(\ID_EX_csr [11] ), .ZN(_02657_ ) );
INV_X1 _10399_ ( .A(\ID_EX_csr [3] ), .ZN(_02658_ ) );
AOI22_X1 _10400_ ( .A1(\EX_LS_dest_csreg_mem [11] ), .A2(_02657_ ), .B1(_02658_ ), .B2(\EX_LS_dest_csreg_mem [3] ), .ZN(_02659_ ) );
AND4_X1 _10401_ ( .A1(_01676_ ), .A2(_02655_ ), .A3(_02656_ ), .A4(_02659_ ), .ZN(_02660_ ) );
XNOR2_X1 _10402_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_02661_ ) );
XNOR2_X1 _10403_ ( .A(fanout_net_6 ), .B(\ID_EX_csr [0] ), .ZN(_02662_ ) );
AND4_X2 _10404_ ( .A1(_02653_ ), .A2(_02660_ ), .A3(_02661_ ), .A4(_02662_ ), .ZN(_02663_ ) );
AND2_X1 _10405_ ( .A1(_02652_ ), .A2(_02663_ ), .ZN(_02664_ ) );
INV_X2 _10406_ ( .A(_02664_ ), .ZN(_02665_ ) );
AND2_X1 _10407_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_02666_ ) );
AND3_X1 _10408_ ( .A1(_02666_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_02667_ ) );
NOR3_X1 _10409_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .A3(\ID_EX_csr [5] ), .ZN(_02668_ ) );
AND3_X1 _10410_ ( .A1(_02667_ ), .A2(\ID_EX_csr [4] ), .A3(_02668_ ), .ZN(_02669_ ) );
INV_X1 _10411_ ( .A(\ID_EX_csr [0] ), .ZN(_02670_ ) );
NOR2_X1 _10412_ ( .A1(_02670_ ), .A2(\ID_EX_csr [1] ), .ZN(_02671_ ) );
NOR2_X1 _10413_ ( .A1(\ID_EX_csr [3] ), .A2(\ID_EX_csr [2] ), .ZN(_02672_ ) );
AND2_X1 _10414_ ( .A1(_02671_ ), .A2(_02672_ ), .ZN(_02673_ ) );
AND2_X1 _10415_ ( .A1(_02669_ ), .A2(_02673_ ), .ZN(_02674_ ) );
BUF_X4 _10416_ ( .A(_02674_ ), .Z(_02675_ ) );
INV_X1 _10417_ ( .A(_02675_ ), .ZN(_02676_ ) );
AND3_X2 _10418_ ( .A1(_02671_ ), .A2(_02658_ ), .A3(\ID_EX_csr [2] ), .ZN(_02677_ ) );
BUF_X2 _10419_ ( .A(_02677_ ), .Z(_02678_ ) );
INV_X1 _10420_ ( .A(\ID_EX_csr [4] ), .ZN(_02679_ ) );
AND2_X2 _10421_ ( .A1(_02668_ ), .A2(_02679_ ), .ZN(_02680_ ) );
BUF_X4 _10422_ ( .A(_02680_ ), .Z(_02681_ ) );
BUF_X4 _10423_ ( .A(_02681_ ), .Z(_02682_ ) );
BUF_X4 _10424_ ( .A(_02682_ ), .Z(_02683_ ) );
NOR2_X1 _10425_ ( .A1(\ID_EX_csr [10] ), .A2(\ID_EX_csr [11] ), .ZN(_02684_ ) );
AND2_X1 _10426_ ( .A1(_02666_ ), .A2(_02684_ ), .ZN(_02685_ ) );
BUF_X4 _10427_ ( .A(_02685_ ), .Z(_02686_ ) );
BUF_X4 _10428_ ( .A(_02686_ ), .Z(_02687_ ) );
BUF_X2 _10429_ ( .A(_02687_ ), .Z(_02688_ ) );
NAND4_X1 _10430_ ( .A1(_02678_ ), .A2(_02683_ ), .A3(\mtvec [30] ), .A4(_02688_ ), .ZN(_02689_ ) );
BUF_X4 _10431_ ( .A(_02673_ ), .Z(_02690_ ) );
BUF_X4 _10432_ ( .A(_02690_ ), .Z(_02691_ ) );
INV_X1 _10433_ ( .A(\ID_EX_csr [6] ), .ZN(_02692_ ) );
NOR2_X1 _10434_ ( .A1(_02692_ ), .A2(\ID_EX_csr [7] ), .ZN(_02693_ ) );
NOR2_X1 _10435_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_02694_ ) );
AND2_X1 _10436_ ( .A1(_02693_ ), .A2(_02694_ ), .ZN(_02695_ ) );
BUF_X4 _10437_ ( .A(_02695_ ), .Z(_02696_ ) );
BUF_X4 _10438_ ( .A(_02696_ ), .Z(_02697_ ) );
BUF_X4 _10439_ ( .A(_02697_ ), .Z(_02698_ ) );
NAND4_X1 _10440_ ( .A1(_02691_ ), .A2(_02698_ ), .A3(\mepc [30] ), .A4(_02688_ ), .ZN(_02699_ ) );
BUF_X4 _10441_ ( .A(_02686_ ), .Z(_02700_ ) );
BUF_X4 _10442_ ( .A(_02700_ ), .Z(_02701_ ) );
AND3_X2 _10443_ ( .A1(_02672_ ), .A2(_02642_ ), .A3(_02670_ ), .ZN(_02702_ ) );
BUF_X4 _10444_ ( .A(_02702_ ), .Z(_02703_ ) );
NAND4_X1 _10445_ ( .A1(_02682_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_02701_ ), .A4(_02703_ ), .ZN(_02704_ ) );
BUF_X4 _10446_ ( .A(_02696_ ), .Z(_02705_ ) );
NOR2_X1 _10447_ ( .A1(_02642_ ), .A2(\ID_EX_csr [0] ), .ZN(_02706_ ) );
AND2_X2 _10448_ ( .A1(_02706_ ), .A2(_02672_ ), .ZN(_02707_ ) );
BUF_X2 _10449_ ( .A(_02707_ ), .Z(_02708_ ) );
BUF_X4 _10450_ ( .A(_02700_ ), .Z(_02709_ ) );
NAND4_X1 _10451_ ( .A1(_02705_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][30] ), .A4(_02709_ ), .ZN(_02710_ ) );
AND2_X1 _10452_ ( .A1(_02704_ ), .A2(_02710_ ), .ZN(_02711_ ) );
NAND4_X1 _10453_ ( .A1(_02676_ ), .A2(_02689_ ), .A3(_02699_ ), .A4(_02711_ ), .ZN(_02712_ ) );
NAND2_X1 _10454_ ( .A1(_02665_ ), .A2(_02712_ ), .ZN(_02713_ ) );
BUF_X2 _10455_ ( .A(_02652_ ), .Z(_02714_ ) );
BUF_X4 _10456_ ( .A(_02714_ ), .Z(_02715_ ) );
BUF_X2 _10457_ ( .A(_02663_ ), .Z(_02716_ ) );
BUF_X4 _10458_ ( .A(_02716_ ), .Z(_02717_ ) );
NAND3_X1 _10459_ ( .A1(_02715_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_02717_ ), .ZN(_02718_ ) );
AND2_X1 _10460_ ( .A1(_02713_ ), .A2(_02718_ ), .ZN(_02719_ ) );
BUF_X4 _10461_ ( .A(_01652_ ), .Z(_02720_ ) );
NOR2_X1 _10462_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_02721_ ) );
XOR2_X1 _10463_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_02722_ ) );
NOR2_X1 _10464_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_02723_ ) );
XOR2_X1 _10465_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_02724_ ) );
XOR2_X1 _10466_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_02725_ ) );
AND2_X1 _10467_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_02726_ ) );
AND2_X1 _10468_ ( .A1(_02725_ ), .A2(_02726_ ), .ZN(_02727_ ) );
AND2_X1 _10469_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_02728_ ) );
OAI21_X1 _10470_ ( .A(_02724_ ), .B1(_02727_ ), .B2(_02728_ ), .ZN(_02729_ ) );
NAND2_X1 _10471_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_02730_ ) );
NAND2_X1 _10472_ ( .A1(_02729_ ), .A2(_02730_ ), .ZN(_02731_ ) );
OAI21_X1 _10473_ ( .A(_02731_ ), .B1(\ID_EX_pc [3] ), .B2(\ID_EX_imm [3] ), .ZN(_02732_ ) );
AND2_X1 _10474_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_02733_ ) );
INV_X1 _10475_ ( .A(_02733_ ), .ZN(_02734_ ) );
NAND2_X1 _10476_ ( .A1(_02732_ ), .A2(_02734_ ), .ZN(_02735_ ) );
XOR2_X1 _10477_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_02736_ ) );
NAND2_X1 _10478_ ( .A1(_02735_ ), .A2(_02736_ ), .ZN(_02737_ ) );
NAND2_X1 _10479_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_02738_ ) );
AOI21_X1 _10480_ ( .A(_02723_ ), .B1(_02737_ ), .B2(_02738_ ), .ZN(_02739_ ) );
AND2_X1 _10481_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_02740_ ) );
OAI21_X1 _10482_ ( .A(_02722_ ), .B1(_02739_ ), .B2(_02740_ ), .ZN(_02741_ ) );
NAND2_X1 _10483_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_02742_ ) );
AOI21_X1 _10484_ ( .A(_02721_ ), .B1(_02741_ ), .B2(_02742_ ), .ZN(_02743_ ) );
AND2_X1 _10485_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_02744_ ) );
OR2_X1 _10486_ ( .A1(_02743_ ), .A2(_02744_ ), .ZN(_02745_ ) );
XOR2_X1 _10487_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_02746_ ) );
XOR2_X1 _10488_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_02747_ ) );
AND2_X1 _10489_ ( .A1(_02746_ ), .A2(_02747_ ), .ZN(_02748_ ) );
XOR2_X1 _10490_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_02749_ ) );
XOR2_X1 _10491_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_02750_ ) );
AND2_X1 _10492_ ( .A1(_02749_ ), .A2(_02750_ ), .ZN(_02751_ ) );
AND3_X1 _10493_ ( .A1(_02745_ ), .A2(_02748_ ), .A3(_02751_ ), .ZN(_02752_ ) );
AND2_X1 _10494_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_02753_ ) );
AND2_X1 _10495_ ( .A1(_02746_ ), .A2(_02753_ ), .ZN(_02754_ ) );
AOI21_X1 _10496_ ( .A(_02754_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_02755_ ) );
AND2_X1 _10497_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_02756_ ) );
AND2_X1 _10498_ ( .A1(_02750_ ), .A2(_02756_ ), .ZN(_02757_ ) );
AOI21_X1 _10499_ ( .A(_02757_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_02758_ ) );
INV_X1 _10500_ ( .A(_02748_ ), .ZN(_02759_ ) );
OAI21_X1 _10501_ ( .A(_02755_ ), .B1(_02758_ ), .B2(_02759_ ), .ZN(_02760_ ) );
OR2_X1 _10502_ ( .A1(_02752_ ), .A2(_02760_ ), .ZN(_02761_ ) );
XOR2_X1 _10503_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_02762_ ) );
XOR2_X1 _10504_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_02763_ ) );
AND2_X1 _10505_ ( .A1(_02762_ ), .A2(_02763_ ), .ZN(_02764_ ) );
XOR2_X1 _10506_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .Z(_02765_ ) );
XOR2_X1 _10507_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_02766_ ) );
AND2_X1 _10508_ ( .A1(_02765_ ), .A2(_02766_ ), .ZN(_02767_ ) );
AND3_X1 _10509_ ( .A1(_02761_ ), .A2(_02764_ ), .A3(_02767_ ), .ZN(_02768_ ) );
AND2_X1 _10510_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_02769_ ) );
AND2_X1 _10511_ ( .A1(_02762_ ), .A2(_02769_ ), .ZN(_02770_ ) );
AOI21_X1 _10512_ ( .A(_02770_ ), .B1(\ID_EX_pc [15] ), .B2(\ID_EX_imm [15] ), .ZN(_02771_ ) );
AND3_X1 _10513_ ( .A1(_02765_ ), .A2(\ID_EX_pc [12] ), .A3(\ID_EX_imm [12] ), .ZN(_02772_ ) );
AOI21_X1 _10514_ ( .A(_02772_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_02773_ ) );
INV_X1 _10515_ ( .A(_02764_ ), .ZN(_02774_ ) );
OAI21_X1 _10516_ ( .A(_02771_ ), .B1(_02773_ ), .B2(_02774_ ), .ZN(_02775_ ) );
OR2_X1 _10517_ ( .A1(_02768_ ), .A2(_02775_ ), .ZN(_02776_ ) );
XOR2_X1 _10518_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_02777_ ) );
XOR2_X1 _10519_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_02778_ ) );
AND2_X1 _10520_ ( .A1(_02777_ ), .A2(_02778_ ), .ZN(_02779_ ) );
XOR2_X1 _10521_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_02780_ ) );
XOR2_X1 _10522_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_02781_ ) );
AND2_X1 _10523_ ( .A1(_02780_ ), .A2(_02781_ ), .ZN(_02782_ ) );
AND3_X1 _10524_ ( .A1(_02776_ ), .A2(_02779_ ), .A3(_02782_ ), .ZN(_02783_ ) );
AND2_X1 _10525_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_02784_ ) );
AND2_X1 _10526_ ( .A1(_02777_ ), .A2(_02784_ ), .ZN(_02785_ ) );
AOI21_X1 _10527_ ( .A(_02785_ ), .B1(\ID_EX_pc [19] ), .B2(\ID_EX_imm [19] ), .ZN(_02786_ ) );
AND2_X1 _10528_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_02787_ ) );
AND2_X1 _10529_ ( .A1(_02781_ ), .A2(_02787_ ), .ZN(_02788_ ) );
AOI21_X1 _10530_ ( .A(_02788_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_02789_ ) );
INV_X1 _10531_ ( .A(_02779_ ), .ZN(_02790_ ) );
OAI21_X1 _10532_ ( .A(_02786_ ), .B1(_02789_ ), .B2(_02790_ ), .ZN(_02791_ ) );
OR2_X1 _10533_ ( .A1(_02783_ ), .A2(_02791_ ), .ZN(_02792_ ) );
XOR2_X1 _10534_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_02793_ ) );
XOR2_X1 _10535_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_02794_ ) );
XOR2_X1 _10536_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_02795_ ) );
XOR2_X1 _10537_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_02796_ ) );
AND2_X1 _10538_ ( .A1(_02795_ ), .A2(_02796_ ), .ZN(_02797_ ) );
NAND4_X1 _10539_ ( .A1(_02792_ ), .A2(_02793_ ), .A3(_02794_ ), .A4(_02797_ ), .ZN(_02798_ ) );
AND2_X1 _10540_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_02799_ ) );
AND2_X1 _10541_ ( .A1(_02796_ ), .A2(_02799_ ), .ZN(_02800_ ) );
AOI21_X1 _10542_ ( .A(_02800_ ), .B1(\ID_EX_pc [21] ), .B2(\ID_EX_imm [21] ), .ZN(_02801_ ) );
NAND2_X1 _10543_ ( .A1(_02793_ ), .A2(_02794_ ), .ZN(_02802_ ) );
NOR2_X1 _10544_ ( .A1(_02801_ ), .A2(_02802_ ), .ZN(_02803_ ) );
AND2_X1 _10545_ ( .A1(\ID_EX_pc [23] ), .A2(\ID_EX_imm [23] ), .ZN(_02804_ ) );
AND2_X1 _10546_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_02805_ ) );
AND2_X1 _10547_ ( .A1(_02793_ ), .A2(_02805_ ), .ZN(_02806_ ) );
NOR3_X1 _10548_ ( .A1(_02803_ ), .A2(_02804_ ), .A3(_02806_ ), .ZN(_02807_ ) );
NAND2_X1 _10549_ ( .A1(_02798_ ), .A2(_02807_ ), .ZN(_02808_ ) );
XOR2_X1 _10550_ ( .A(\ID_EX_pc [25] ), .B(\ID_EX_imm [25] ), .Z(_02809_ ) );
XOR2_X1 _10551_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_02810_ ) );
NAND3_X1 _10552_ ( .A1(_02808_ ), .A2(_02809_ ), .A3(_02810_ ), .ZN(_02811_ ) );
AND2_X1 _10553_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_02812_ ) );
AND2_X1 _10554_ ( .A1(_02809_ ), .A2(_02812_ ), .ZN(_02813_ ) );
AOI21_X1 _10555_ ( .A(_02813_ ), .B1(\ID_EX_pc [25] ), .B2(\ID_EX_imm [25] ), .ZN(_02814_ ) );
NAND2_X1 _10556_ ( .A1(_02811_ ), .A2(_02814_ ), .ZN(_02815_ ) );
XOR2_X1 _10557_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_02816_ ) );
XOR2_X1 _10558_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_02817_ ) );
NAND3_X1 _10559_ ( .A1(_02815_ ), .A2(_02816_ ), .A3(_02817_ ), .ZN(_02818_ ) );
AND3_X1 _10560_ ( .A1(_02816_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_02819_ ) );
AOI21_X1 _10561_ ( .A(_02819_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_02820_ ) );
NAND2_X1 _10562_ ( .A1(_02818_ ), .A2(_02820_ ), .ZN(_02821_ ) );
XOR2_X1 _10563_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_02822_ ) );
NAND2_X1 _10564_ ( .A1(_02821_ ), .A2(_02822_ ), .ZN(_02823_ ) );
NAND2_X1 _10565_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_02824_ ) );
INV_X1 _10566_ ( .A(\ID_EX_pc [29] ), .ZN(_02825_ ) );
AOI22_X1 _10567_ ( .A1(_02823_ ), .A2(_02824_ ), .B1(_02825_ ), .B2(_02540_ ), .ZN(_02826_ ) );
AND2_X1 _10568_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_02827_ ) );
OR2_X1 _10569_ ( .A1(_02826_ ), .A2(_02827_ ), .ZN(_02828_ ) );
XOR2_X1 _10570_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_02829_ ) );
XOR2_X1 _10571_ ( .A(_02828_ ), .B(_02829_ ), .Z(_02830_ ) );
INV_X1 _10572_ ( .A(_02830_ ), .ZN(_02831_ ) );
INV_X2 _10573_ ( .A(fanout_net_8 ), .ZN(_02832_ ) );
BUF_X4 _10574_ ( .A(_02832_ ), .Z(_02833_ ) );
AOI21_X1 _10575_ ( .A(_02720_ ), .B1(_02831_ ), .B2(_02833_ ), .ZN(_02834_ ) );
BUF_X4 _10576_ ( .A(_02832_ ), .Z(_02835_ ) );
OAI21_X1 _10577_ ( .A(_02834_ ), .B1(_02583_ ), .B2(_02835_ ), .ZN(_02836_ ) );
INV_X1 _10578_ ( .A(_02578_ ), .ZN(_02837_ ) );
BUF_X4 _10579_ ( .A(_02837_ ), .Z(_02838_ ) );
AND2_X1 _10580_ ( .A1(_02836_ ), .A2(_02838_ ), .ZN(_02839_ ) );
BUF_X4 _10581_ ( .A(_02720_ ), .Z(_02840_ ) );
AND2_X1 _10582_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_02841_ ) );
AND2_X1 _10583_ ( .A1(_02841_ ), .A2(\ID_EX_pc [4] ), .ZN(_02842_ ) );
AND2_X1 _10584_ ( .A1(_02842_ ), .A2(\ID_EX_pc [5] ), .ZN(_02843_ ) );
AND2_X1 _10585_ ( .A1(_02843_ ), .A2(\ID_EX_pc [6] ), .ZN(_02844_ ) );
AND2_X1 _10586_ ( .A1(_02844_ ), .A2(\ID_EX_pc [7] ), .ZN(_02845_ ) );
AND2_X1 _10587_ ( .A1(_02845_ ), .A2(\ID_EX_pc [8] ), .ZN(_02846_ ) );
AND2_X2 _10588_ ( .A1(_02846_ ), .A2(\ID_EX_pc [9] ), .ZN(_02847_ ) );
AND3_X1 _10589_ ( .A1(_02847_ ), .A2(\ID_EX_pc [11] ), .A3(\ID_EX_pc [10] ), .ZN(_02848_ ) );
AND3_X1 _10590_ ( .A1(_02848_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_02849_ ) );
AND3_X1 _10591_ ( .A1(_02849_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_02850_ ) );
AND3_X1 _10592_ ( .A1(_02850_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_02851_ ) );
AND3_X1 _10593_ ( .A1(_02851_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_02852_ ) );
AND3_X1 _10594_ ( .A1(_02852_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_02853_ ) );
AND3_X1 _10595_ ( .A1(_02853_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_02854_ ) );
AND3_X1 _10596_ ( .A1(_02854_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_02855_ ) );
AND3_X1 _10597_ ( .A1(_02855_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_02856_ ) );
NAND3_X1 _10598_ ( .A1(_02856_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_02857_ ) );
XNOR2_X1 _10599_ ( .A(_02857_ ), .B(\ID_EX_pc [30] ), .ZN(_02858_ ) );
NOR2_X1 _10600_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_8 ), .ZN(_02859_ ) );
AND2_X1 _10601_ ( .A1(_02859_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_02860_ ) );
INV_X1 _10602_ ( .A(_02860_ ), .ZN(_02861_ ) );
INV_X32 _10603_ ( .A(fanout_net_25 ), .ZN(_02862_ ) );
BUF_X4 _10604_ ( .A(_02862_ ), .Z(_02863_ ) );
BUF_X8 _10605_ ( .A(_02863_ ), .Z(_02864_ ) );
OR2_X1 _10606_ ( .A1(_02864_ ), .A2(\myreg.Reg[11][17] ), .ZN(_02865_ ) );
OAI211_X1 _10607_ ( .A(_02865_ ), .B(fanout_net_33 ), .C1(fanout_net_25 ), .C2(\myreg.Reg[10][17] ), .ZN(_02866_ ) );
INV_X2 _10608_ ( .A(fanout_net_36 ), .ZN(_02867_ ) );
BUF_X4 _10609_ ( .A(_02867_ ), .Z(_02868_ ) );
BUF_X4 _10610_ ( .A(_02868_ ), .Z(_02869_ ) );
OR2_X1 _10611_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[8][17] ), .ZN(_02870_ ) );
INV_X2 _10612_ ( .A(fanout_net_33 ), .ZN(_02871_ ) );
BUF_X4 _10613_ ( .A(_02871_ ), .Z(_02872_ ) );
BUF_X4 _10614_ ( .A(_02872_ ), .Z(_02873_ ) );
BUF_X4 _10615_ ( .A(_02863_ ), .Z(_02874_ ) );
BUF_X2 _10616_ ( .A(_02874_ ), .Z(_02875_ ) );
OAI211_X1 _10617_ ( .A(_02870_ ), .B(_02873_ ), .C1(_02875_ ), .C2(\myreg.Reg[9][17] ), .ZN(_02876_ ) );
NAND3_X1 _10618_ ( .A1(_02866_ ), .A2(_02869_ ), .A3(_02876_ ), .ZN(_02877_ ) );
MUX2_X1 _10619_ ( .A(\myreg.Reg[14][17] ), .B(\myreg.Reg[15][17] ), .S(fanout_net_25 ), .Z(_02878_ ) );
MUX2_X1 _10620_ ( .A(\myreg.Reg[12][17] ), .B(\myreg.Reg[13][17] ), .S(fanout_net_25 ), .Z(_02879_ ) );
BUF_X4 _10621_ ( .A(_02871_ ), .Z(_02880_ ) );
BUF_X4 _10622_ ( .A(_02880_ ), .Z(_02881_ ) );
MUX2_X1 _10623_ ( .A(_02878_ ), .B(_02879_ ), .S(_02881_ ), .Z(_02882_ ) );
BUF_X4 _10624_ ( .A(_02868_ ), .Z(_02883_ ) );
OAI211_X1 _10625_ ( .A(fanout_net_37 ), .B(_02877_ ), .C1(_02882_ ), .C2(_02883_ ), .ZN(_02884_ ) );
MUX2_X1 _10626_ ( .A(\myreg.Reg[0][17] ), .B(\myreg.Reg[1][17] ), .S(fanout_net_25 ), .Z(_02885_ ) );
AND2_X1 _10627_ ( .A1(_02885_ ), .A2(_02873_ ), .ZN(_02886_ ) );
MUX2_X1 _10628_ ( .A(\myreg.Reg[2][17] ), .B(\myreg.Reg[3][17] ), .S(fanout_net_25 ), .Z(_02887_ ) );
AOI211_X1 _10629_ ( .A(fanout_net_36 ), .B(_02886_ ), .C1(fanout_net_33 ), .C2(_02887_ ), .ZN(_02888_ ) );
INV_X1 _10630_ ( .A(fanout_net_37 ), .ZN(_02889_ ) );
BUF_X4 _10631_ ( .A(_02889_ ), .Z(_02890_ ) );
MUX2_X1 _10632_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_25 ), .Z(_02891_ ) );
MUX2_X1 _10633_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_25 ), .Z(_02892_ ) );
MUX2_X1 _10634_ ( .A(_02891_ ), .B(_02892_ ), .S(_02881_ ), .Z(_02893_ ) );
OAI21_X1 _10635_ ( .A(_02890_ ), .B1(_02893_ ), .B2(_02883_ ), .ZN(_02894_ ) );
OAI21_X1 _10636_ ( .A(_02884_ ), .B1(_02888_ ), .B2(_02894_ ), .ZN(_02895_ ) );
INV_X1 _10637_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .ZN(_02896_ ) );
BUF_X2 _10638_ ( .A(_02896_ ), .Z(_02897_ ) );
BUF_X4 _10639_ ( .A(_02897_ ), .Z(_02898_ ) );
BUF_X4 _10640_ ( .A(_02898_ ), .Z(_02899_ ) );
XNOR2_X1 _10641_ ( .A(\EX_LS_dest_reg [1] ), .B(\ID_EX_rs2 [1] ), .ZN(_02900_ ) );
XOR2_X2 _10642_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .Z(_02901_ ) );
INV_X2 _10643_ ( .A(_02901_ ), .ZN(_02902_ ) );
XNOR2_X1 _10644_ ( .A(\EX_LS_dest_reg [3] ), .B(\ID_EX_rs2 [3] ), .ZN(_02903_ ) );
XNOR2_X1 _10645_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_02904_ ) );
AND4_X4 _10646_ ( .A1(_02900_ ), .A2(_02902_ ), .A3(_02903_ ), .A4(_02904_ ), .ZN(_02905_ ) );
AND2_X1 _10647_ ( .A1(_01665_ ), .A2(_01664_ ), .ZN(_02906_ ) );
INV_X1 _10648_ ( .A(_02906_ ), .ZN(_02907_ ) );
XNOR2_X2 _10649_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_02908_ ) );
NAND4_X4 _10650_ ( .A1(_02905_ ), .A2(_02012_ ), .A3(_02907_ ), .A4(_02908_ ), .ZN(_02909_ ) );
BUF_X8 _10651_ ( .A(_02909_ ), .Z(_02910_ ) );
BUF_X16 _10652_ ( .A(_02910_ ), .Z(_02911_ ) );
BUF_X32 _10653_ ( .A(_02911_ ), .Z(_02912_ ) );
OAI21_X2 _10654_ ( .A(_02895_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_02913_ ) );
INV_X1 _10655_ ( .A(\ID_EX_rs2 [2] ), .ZN(_02914_ ) );
NOR2_X1 _10656_ ( .A1(_02914_ ), .A2(\EX_LS_dest_reg [2] ), .ZN(_02915_ ) );
NOR3_X1 _10657_ ( .A1(_02901_ ), .A2(_02896_ ), .A3(_02915_ ), .ZN(_02916_ ) );
AND3_X1 _10658_ ( .A1(_02916_ ), .A2(_02908_ ), .A3(_02900_ ), .ZN(_02917_ ) );
NAND2_X1 _10659_ ( .A1(_02914_ ), .A2(\EX_LS_dest_reg [2] ), .ZN(_02918_ ) );
AND4_X4 _10660_ ( .A1(_02907_ ), .A2(_02917_ ), .A3(_02903_ ), .A4(_02918_ ), .ZN(_02919_ ) );
NAND3_X1 _10661_ ( .A1(_02919_ ), .A2(\EX_LS_result_reg [17] ), .A3(_02037_ ), .ZN(_02920_ ) );
AND2_X1 _10662_ ( .A1(_02913_ ), .A2(_02920_ ), .ZN(_02921_ ) );
INV_X4 _10663_ ( .A(_01942_ ), .ZN(_02922_ ) );
XNOR2_X1 _10664_ ( .A(_02921_ ), .B(_02922_ ), .ZN(_02923_ ) );
BUF_X8 _10665_ ( .A(_02910_ ), .Z(_02924_ ) );
INV_X1 _10666_ ( .A(\EX_LS_result_reg [16] ), .ZN(_02925_ ) );
BUF_X2 _10667_ ( .A(_02897_ ), .Z(_02926_ ) );
OR3_X1 _10668_ ( .A1(_02924_ ), .A2(_02925_ ), .A3(_02926_ ), .ZN(_02927_ ) );
OR2_X1 _10669_ ( .A1(_02864_ ), .A2(\myreg.Reg[1][16] ), .ZN(_02928_ ) );
BUF_X4 _10670_ ( .A(_02880_ ), .Z(_02929_ ) );
BUF_X4 _10671_ ( .A(_02929_ ), .Z(_02930_ ) );
OAI211_X1 _10672_ ( .A(_02928_ ), .B(_02930_ ), .C1(fanout_net_25 ), .C2(\myreg.Reg[0][16] ), .ZN(_02931_ ) );
OR2_X1 _10673_ ( .A1(_02864_ ), .A2(\myreg.Reg[3][16] ), .ZN(_02932_ ) );
OAI211_X1 _10674_ ( .A(_02932_ ), .B(fanout_net_33 ), .C1(fanout_net_25 ), .C2(\myreg.Reg[2][16] ), .ZN(_02933_ ) );
NAND3_X1 _10675_ ( .A1(_02931_ ), .A2(_02933_ ), .A3(_02869_ ), .ZN(_02934_ ) );
MUX2_X1 _10676_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_25 ), .Z(_02935_ ) );
MUX2_X1 _10677_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_25 ), .Z(_02936_ ) );
MUX2_X1 _10678_ ( .A(_02935_ ), .B(_02936_ ), .S(_02873_ ), .Z(_02937_ ) );
BUF_X4 _10679_ ( .A(_02869_ ), .Z(_02938_ ) );
OAI211_X1 _10680_ ( .A(_02890_ ), .B(_02934_ ), .C1(_02937_ ), .C2(_02938_ ), .ZN(_02939_ ) );
OR2_X1 _10681_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[14][16] ), .ZN(_02940_ ) );
BUF_X4 _10682_ ( .A(_02864_ ), .Z(_02941_ ) );
OAI211_X1 _10683_ ( .A(_02940_ ), .B(fanout_net_33 ), .C1(_02941_ ), .C2(\myreg.Reg[15][16] ), .ZN(_02942_ ) );
OR2_X1 _10684_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[12][16] ), .ZN(_02943_ ) );
OAI211_X1 _10685_ ( .A(_02943_ ), .B(_02873_ ), .C1(_02941_ ), .C2(\myreg.Reg[13][16] ), .ZN(_02944_ ) );
NAND3_X1 _10686_ ( .A1(_02942_ ), .A2(_02944_ ), .A3(fanout_net_36 ), .ZN(_02945_ ) );
MUX2_X1 _10687_ ( .A(\myreg.Reg[8][16] ), .B(\myreg.Reg[9][16] ), .S(fanout_net_25 ), .Z(_02946_ ) );
MUX2_X1 _10688_ ( .A(\myreg.Reg[10][16] ), .B(\myreg.Reg[11][16] ), .S(fanout_net_25 ), .Z(_02947_ ) );
MUX2_X1 _10689_ ( .A(_02946_ ), .B(_02947_ ), .S(fanout_net_33 ), .Z(_02948_ ) );
OAI211_X1 _10690_ ( .A(fanout_net_37 ), .B(_02945_ ), .C1(_02948_ ), .C2(fanout_net_36 ), .ZN(_02949_ ) );
NAND2_X1 _10691_ ( .A1(_02939_ ), .A2(_02949_ ), .ZN(_02950_ ) );
OAI21_X4 _10692_ ( .A(_02950_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_02951_ ) );
AND2_X1 _10693_ ( .A1(_02927_ ), .A2(_02951_ ), .ZN(_02952_ ) );
INV_X1 _10694_ ( .A(_01965_ ), .ZN(_02953_ ) );
XNOR2_X1 _10695_ ( .A(_02952_ ), .B(_02953_ ), .ZN(_02954_ ) );
AND2_X1 _10696_ ( .A1(_02923_ ), .A2(_02954_ ), .ZN(_02955_ ) );
OR2_X1 _10697_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[8][19] ), .ZN(_02956_ ) );
OAI211_X1 _10698_ ( .A(_02956_ ), .B(_02930_ ), .C1(_02941_ ), .C2(\myreg.Reg[9][19] ), .ZN(_02957_ ) );
OR2_X1 _10699_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[10][19] ), .ZN(_02958_ ) );
OAI211_X1 _10700_ ( .A(_02958_ ), .B(fanout_net_33 ), .C1(_02941_ ), .C2(\myreg.Reg[11][19] ), .ZN(_02959_ ) );
NAND3_X1 _10701_ ( .A1(_02957_ ), .A2(_02959_ ), .A3(_02883_ ), .ZN(_02960_ ) );
MUX2_X1 _10702_ ( .A(\myreg.Reg[14][19] ), .B(\myreg.Reg[15][19] ), .S(fanout_net_25 ), .Z(_02961_ ) );
MUX2_X1 _10703_ ( .A(\myreg.Reg[12][19] ), .B(\myreg.Reg[13][19] ), .S(fanout_net_25 ), .Z(_02962_ ) );
MUX2_X1 _10704_ ( .A(_02961_ ), .B(_02962_ ), .S(_02930_ ), .Z(_02963_ ) );
OAI211_X1 _10705_ ( .A(fanout_net_37 ), .B(_02960_ ), .C1(_02963_ ), .C2(_02938_ ), .ZN(_02964_ ) );
MUX2_X1 _10706_ ( .A(\myreg.Reg[0][19] ), .B(\myreg.Reg[1][19] ), .S(fanout_net_25 ), .Z(_02965_ ) );
AND2_X1 _10707_ ( .A1(_02965_ ), .A2(_02930_ ), .ZN(_02966_ ) );
MUX2_X1 _10708_ ( .A(\myreg.Reg[2][19] ), .B(\myreg.Reg[3][19] ), .S(fanout_net_25 ), .Z(_02967_ ) );
AOI211_X1 _10709_ ( .A(fanout_net_36 ), .B(_02966_ ), .C1(fanout_net_33 ), .C2(_02967_ ), .ZN(_02968_ ) );
MUX2_X1 _10710_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_25 ), .Z(_02969_ ) );
MUX2_X1 _10711_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_25 ), .Z(_02970_ ) );
MUX2_X1 _10712_ ( .A(_02969_ ), .B(_02970_ ), .S(_02930_ ), .Z(_02971_ ) );
OAI21_X1 _10713_ ( .A(_02890_ ), .B1(_02971_ ), .B2(_02938_ ), .ZN(_02972_ ) );
OAI21_X1 _10714_ ( .A(_02964_ ), .B1(_02968_ ), .B2(_02972_ ), .ZN(_02973_ ) );
OAI21_X1 _10715_ ( .A(_02973_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_02974_ ) );
NAND3_X1 _10716_ ( .A1(_02919_ ), .A2(\EX_LS_result_reg [19] ), .A3(_02037_ ), .ZN(_02975_ ) );
AND2_X1 _10717_ ( .A1(_02974_ ), .A2(_02975_ ), .ZN(_02976_ ) );
INV_X1 _10718_ ( .A(_01918_ ), .ZN(_02977_ ) );
XNOR2_X2 _10719_ ( .A(_02976_ ), .B(_02977_ ), .ZN(_02978_ ) );
OR2_X1 _10720_ ( .A1(_02875_ ), .A2(\myreg.Reg[9][18] ), .ZN(_02979_ ) );
BUF_X4 _10721_ ( .A(_02881_ ), .Z(_02980_ ) );
OAI211_X1 _10722_ ( .A(_02979_ ), .B(_02980_ ), .C1(fanout_net_25 ), .C2(\myreg.Reg[8][18] ), .ZN(_02981_ ) );
BUF_X4 _10723_ ( .A(_02862_ ), .Z(_02982_ ) );
BUF_X2 _10724_ ( .A(_02982_ ), .Z(_02983_ ) );
OR2_X1 _10725_ ( .A1(_02983_ ), .A2(\myreg.Reg[11][18] ), .ZN(_02984_ ) );
OAI211_X1 _10726_ ( .A(_02984_ ), .B(fanout_net_33 ), .C1(fanout_net_25 ), .C2(\myreg.Reg[10][18] ), .ZN(_02985_ ) );
NAND3_X1 _10727_ ( .A1(_02981_ ), .A2(_02985_ ), .A3(_02883_ ), .ZN(_02986_ ) );
MUX2_X1 _10728_ ( .A(\myreg.Reg[14][18] ), .B(\myreg.Reg[15][18] ), .S(fanout_net_25 ), .Z(_02987_ ) );
MUX2_X1 _10729_ ( .A(\myreg.Reg[12][18] ), .B(\myreg.Reg[13][18] ), .S(fanout_net_25 ), .Z(_02988_ ) );
MUX2_X1 _10730_ ( .A(_02987_ ), .B(_02988_ ), .S(_02980_ ), .Z(_02989_ ) );
OAI211_X1 _10731_ ( .A(fanout_net_37 ), .B(_02986_ ), .C1(_02989_ ), .C2(_02938_ ), .ZN(_02990_ ) );
MUX2_X1 _10732_ ( .A(\myreg.Reg[2][18] ), .B(\myreg.Reg[3][18] ), .S(fanout_net_25 ), .Z(_02991_ ) );
AND2_X1 _10733_ ( .A1(_02991_ ), .A2(fanout_net_33 ), .ZN(_02992_ ) );
BUF_X4 _10734_ ( .A(_02980_ ), .Z(_02993_ ) );
MUX2_X1 _10735_ ( .A(\myreg.Reg[0][18] ), .B(\myreg.Reg[1][18] ), .S(fanout_net_26 ), .Z(_02994_ ) );
AOI211_X1 _10736_ ( .A(fanout_net_36 ), .B(_02992_ ), .C1(_02993_ ), .C2(_02994_ ), .ZN(_02995_ ) );
BUF_X4 _10737_ ( .A(_02890_ ), .Z(_02996_ ) );
MUX2_X1 _10738_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_26 ), .Z(_02997_ ) );
MUX2_X1 _10739_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_26 ), .Z(_02998_ ) );
MUX2_X1 _10740_ ( .A(_02997_ ), .B(_02998_ ), .S(_02980_ ), .Z(_02999_ ) );
OAI21_X1 _10741_ ( .A(_02996_ ), .B1(_02999_ ), .B2(_02938_ ), .ZN(_03000_ ) );
OAI21_X1 _10742_ ( .A(_02990_ ), .B1(_02995_ ), .B2(_03000_ ), .ZN(_03001_ ) );
OAI21_X1 _10743_ ( .A(_03001_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_03002_ ) );
NAND3_X1 _10744_ ( .A1(_02919_ ), .A2(\EX_LS_result_reg [18] ), .A3(_02037_ ), .ZN(_03003_ ) );
AND2_X1 _10745_ ( .A1(_03002_ ), .A2(_03003_ ), .ZN(_03004_ ) );
INV_X1 _10746_ ( .A(_01895_ ), .ZN(_03005_ ) );
XNOR2_X2 _10747_ ( .A(_03004_ ), .B(_03005_ ), .ZN(_03006_ ) );
AND3_X2 _10748_ ( .A1(_02955_ ), .A2(_02978_ ), .A3(_03006_ ), .ZN(_03007_ ) );
INV_X1 _10749_ ( .A(_03007_ ), .ZN(_03008_ ) );
NAND3_X1 _10750_ ( .A1(_02919_ ), .A2(\EX_LS_result_reg [22] ), .A3(_02037_ ), .ZN(_03009_ ) );
NOR2_X1 _10751_ ( .A1(_02864_ ), .A2(\myreg.Reg[11][22] ), .ZN(_03010_ ) );
OAI21_X1 _10752_ ( .A(fanout_net_33 ), .B1(fanout_net_26 ), .B2(\myreg.Reg[10][22] ), .ZN(_03011_ ) );
NOR2_X1 _10753_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[8][22] ), .ZN(_03012_ ) );
OAI21_X1 _10754_ ( .A(_02872_ ), .B1(_02864_ ), .B2(\myreg.Reg[9][22] ), .ZN(_03013_ ) );
OAI221_X1 _10755_ ( .A(_02868_ ), .B1(_03010_ ), .B2(_03011_ ), .C1(_03012_ ), .C2(_03013_ ), .ZN(_03014_ ) );
MUX2_X1 _10756_ ( .A(\myreg.Reg[12][22] ), .B(\myreg.Reg[13][22] ), .S(fanout_net_26 ), .Z(_03015_ ) );
MUX2_X1 _10757_ ( .A(\myreg.Reg[14][22] ), .B(\myreg.Reg[15][22] ), .S(fanout_net_26 ), .Z(_03016_ ) );
MUX2_X1 _10758_ ( .A(_03015_ ), .B(_03016_ ), .S(fanout_net_33 ), .Z(_03017_ ) );
OAI211_X1 _10759_ ( .A(fanout_net_37 ), .B(_03014_ ), .C1(_03017_ ), .C2(_02869_ ), .ZN(_03018_ ) );
BUF_X4 _10760_ ( .A(_02889_ ), .Z(_03019_ ) );
OR2_X1 _10761_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[4][22] ), .ZN(_03020_ ) );
BUF_X4 _10762_ ( .A(_02982_ ), .Z(_03021_ ) );
OAI211_X1 _10763_ ( .A(_03020_ ), .B(_02929_ ), .C1(_03021_ ), .C2(\myreg.Reg[5][22] ), .ZN(_03022_ ) );
OR2_X1 _10764_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[6][22] ), .ZN(_03023_ ) );
OAI211_X1 _10765_ ( .A(_03023_ ), .B(fanout_net_33 ), .C1(_02864_ ), .C2(\myreg.Reg[7][22] ), .ZN(_03024_ ) );
NAND3_X1 _10766_ ( .A1(_03022_ ), .A2(_03024_ ), .A3(fanout_net_36 ), .ZN(_03025_ ) );
MUX2_X1 _10767_ ( .A(\myreg.Reg[2][22] ), .B(\myreg.Reg[3][22] ), .S(fanout_net_26 ), .Z(_03026_ ) );
MUX2_X1 _10768_ ( .A(\myreg.Reg[0][22] ), .B(\myreg.Reg[1][22] ), .S(fanout_net_26 ), .Z(_03027_ ) );
MUX2_X1 _10769_ ( .A(_03026_ ), .B(_03027_ ), .S(_02872_ ), .Z(_03028_ ) );
OAI211_X1 _10770_ ( .A(_03019_ ), .B(_03025_ ), .C1(_03028_ ), .C2(fanout_net_36 ), .ZN(_03029_ ) );
NAND2_X1 _10771_ ( .A1(_03018_ ), .A2(_03029_ ), .ZN(_03030_ ) );
OAI21_X2 _10772_ ( .A(_03030_ ), .B1(_02926_ ), .B2(_02924_ ), .ZN(_03031_ ) );
AND2_X1 _10773_ ( .A1(_03009_ ), .A2(_03031_ ), .ZN(_03032_ ) );
INV_X4 _10774_ ( .A(_01793_ ), .ZN(_03033_ ) );
XNOR2_X1 _10775_ ( .A(_03032_ ), .B(_03033_ ), .ZN(_03034_ ) );
INV_X1 _10776_ ( .A(\EX_LS_result_reg [23] ), .ZN(_03035_ ) );
OR3_X4 _10777_ ( .A1(_02910_ ), .A2(_03035_ ), .A3(_02897_ ), .ZN(_03036_ ) );
OR2_X1 _10778_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[0][23] ), .ZN(_03037_ ) );
OAI211_X1 _10779_ ( .A(_03037_ ), .B(_02880_ ), .C1(_02863_ ), .C2(\myreg.Reg[1][23] ), .ZN(_03038_ ) );
OR2_X1 _10780_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[2][23] ), .ZN(_03039_ ) );
OAI211_X1 _10781_ ( .A(_03039_ ), .B(fanout_net_33 ), .C1(_02863_ ), .C2(\myreg.Reg[3][23] ), .ZN(_03040_ ) );
NAND3_X1 _10782_ ( .A1(_03038_ ), .A2(_03040_ ), .A3(_02867_ ), .ZN(_03041_ ) );
MUX2_X1 _10783_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_26 ), .Z(_03042_ ) );
MUX2_X1 _10784_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_26 ), .Z(_03043_ ) );
MUX2_X1 _10785_ ( .A(_03042_ ), .B(_03043_ ), .S(_02871_ ), .Z(_03044_ ) );
OAI211_X1 _10786_ ( .A(_02889_ ), .B(_03041_ ), .C1(_03044_ ), .C2(_02867_ ), .ZN(_03045_ ) );
OR2_X1 _10787_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[14][23] ), .ZN(_03046_ ) );
OAI211_X1 _10788_ ( .A(_03046_ ), .B(fanout_net_33 ), .C1(_02863_ ), .C2(\myreg.Reg[15][23] ), .ZN(_03047_ ) );
OR2_X1 _10789_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[12][23] ), .ZN(_03048_ ) );
OAI211_X1 _10790_ ( .A(_03048_ ), .B(_02871_ ), .C1(_02863_ ), .C2(\myreg.Reg[13][23] ), .ZN(_03049_ ) );
NAND3_X1 _10791_ ( .A1(_03047_ ), .A2(_03049_ ), .A3(fanout_net_36 ), .ZN(_03050_ ) );
MUX2_X1 _10792_ ( .A(\myreg.Reg[8][23] ), .B(\myreg.Reg[9][23] ), .S(fanout_net_26 ), .Z(_03051_ ) );
MUX2_X1 _10793_ ( .A(\myreg.Reg[10][23] ), .B(\myreg.Reg[11][23] ), .S(fanout_net_26 ), .Z(_03052_ ) );
MUX2_X1 _10794_ ( .A(_03051_ ), .B(_03052_ ), .S(fanout_net_33 ), .Z(_03053_ ) );
OAI211_X1 _10795_ ( .A(fanout_net_37 ), .B(_03050_ ), .C1(_03053_ ), .C2(fanout_net_36 ), .ZN(_03054_ ) );
NAND2_X1 _10796_ ( .A1(_03045_ ), .A2(_03054_ ), .ZN(_03055_ ) );
OAI21_X1 _10797_ ( .A(_03055_ ), .B1(_02897_ ), .B2(_02910_ ), .ZN(_03056_ ) );
AND2_X2 _10798_ ( .A1(_03036_ ), .A2(_03056_ ), .ZN(_03057_ ) );
INV_X4 _10799_ ( .A(_01816_ ), .ZN(_03058_ ) );
XNOR2_X1 _10800_ ( .A(_03057_ ), .B(_03058_ ), .ZN(_03059_ ) );
AND2_X1 _10801_ ( .A1(_03034_ ), .A2(_03059_ ), .ZN(_03060_ ) );
NOR2_X4 _10802_ ( .A1(_02910_ ), .A2(_02897_ ), .ZN(_03061_ ) );
OR2_X1 _10803_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[0][20] ), .ZN(_03062_ ) );
OAI211_X1 _10804_ ( .A(_03062_ ), .B(_02930_ ), .C1(_02941_ ), .C2(\myreg.Reg[1][20] ), .ZN(_03063_ ) );
OR2_X1 _10805_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[2][20] ), .ZN(_03064_ ) );
OAI211_X1 _10806_ ( .A(_03064_ ), .B(fanout_net_33 ), .C1(_02941_ ), .C2(\myreg.Reg[3][20] ), .ZN(_03065_ ) );
NAND3_X1 _10807_ ( .A1(_03063_ ), .A2(_03065_ ), .A3(_02883_ ), .ZN(_03066_ ) );
MUX2_X1 _10808_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_26 ), .Z(_03067_ ) );
MUX2_X1 _10809_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_26 ), .Z(_03068_ ) );
MUX2_X1 _10810_ ( .A(_03067_ ), .B(_03068_ ), .S(_02873_ ), .Z(_03069_ ) );
OAI211_X1 _10811_ ( .A(_02890_ ), .B(_03066_ ), .C1(_03069_ ), .C2(_02938_ ), .ZN(_03070_ ) );
OR2_X1 _10812_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[14][20] ), .ZN(_03071_ ) );
OAI211_X1 _10813_ ( .A(_03071_ ), .B(fanout_net_33 ), .C1(_02941_ ), .C2(\myreg.Reg[15][20] ), .ZN(_03072_ ) );
OR2_X1 _10814_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[12][20] ), .ZN(_03073_ ) );
OAI211_X1 _10815_ ( .A(_03073_ ), .B(_02930_ ), .C1(_02941_ ), .C2(\myreg.Reg[13][20] ), .ZN(_03074_ ) );
NAND3_X1 _10816_ ( .A1(_03072_ ), .A2(_03074_ ), .A3(fanout_net_36 ), .ZN(_03075_ ) );
MUX2_X1 _10817_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_26 ), .Z(_03076_ ) );
MUX2_X1 _10818_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_26 ), .Z(_03077_ ) );
MUX2_X1 _10819_ ( .A(_03076_ ), .B(_03077_ ), .S(fanout_net_33 ), .Z(_03078_ ) );
OAI211_X1 _10820_ ( .A(fanout_net_37 ), .B(_03075_ ), .C1(_03078_ ), .C2(fanout_net_36 ), .ZN(_03079_ ) );
AOI21_X1 _10821_ ( .A(_03061_ ), .B1(_03070_ ), .B2(_03079_ ), .ZN(_03080_ ) );
INV_X1 _10822_ ( .A(\EX_LS_result_reg [20] ), .ZN(_03081_ ) );
NOR3_X1 _10823_ ( .A1(_02924_ ), .A2(_03081_ ), .A3(_02926_ ), .ZN(_03082_ ) );
NOR2_X1 _10824_ ( .A1(_03080_ ), .A2(_03082_ ), .ZN(_03083_ ) );
INV_X1 _10825_ ( .A(_01869_ ), .ZN(_03084_ ) );
XNOR2_X1 _10826_ ( .A(_03083_ ), .B(_03084_ ), .ZN(_03085_ ) );
INV_X1 _10827_ ( .A(\EX_LS_result_reg [21] ), .ZN(_03086_ ) );
OR3_X1 _10828_ ( .A1(_02924_ ), .A2(_03086_ ), .A3(_02926_ ), .ZN(_03087_ ) );
OR2_X1 _10829_ ( .A1(\myreg.Reg[0][21] ), .A2(fanout_net_26 ), .ZN(_03088_ ) );
OAI211_X1 _10830_ ( .A(_03088_ ), .B(_02873_ ), .C1(\myreg.Reg[1][21] ), .C2(_02875_ ), .ZN(_03089_ ) );
OR2_X1 _10831_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[2][21] ), .ZN(_03090_ ) );
OAI211_X1 _10832_ ( .A(_03090_ ), .B(fanout_net_33 ), .C1(_02875_ ), .C2(\myreg.Reg[3][21] ), .ZN(_03091_ ) );
NAND3_X1 _10833_ ( .A1(_03089_ ), .A2(_03091_ ), .A3(_02869_ ), .ZN(_03092_ ) );
MUX2_X1 _10834_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_26 ), .Z(_03093_ ) );
MUX2_X1 _10835_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_27 ), .Z(_03094_ ) );
MUX2_X1 _10836_ ( .A(_03093_ ), .B(_03094_ ), .S(_02881_ ), .Z(_03095_ ) );
OAI211_X1 _10837_ ( .A(_02890_ ), .B(_03092_ ), .C1(_03095_ ), .C2(_02883_ ), .ZN(_03096_ ) );
OR2_X1 _10838_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[14][21] ), .ZN(_03097_ ) );
OAI211_X1 _10839_ ( .A(_03097_ ), .B(fanout_net_33 ), .C1(_02875_ ), .C2(\myreg.Reg[15][21] ), .ZN(_03098_ ) );
OR2_X1 _10840_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[12][21] ), .ZN(_03099_ ) );
OAI211_X1 _10841_ ( .A(_03099_ ), .B(_02873_ ), .C1(_02875_ ), .C2(\myreg.Reg[13][21] ), .ZN(_03100_ ) );
NAND3_X1 _10842_ ( .A1(_03098_ ), .A2(_03100_ ), .A3(fanout_net_36 ), .ZN(_03101_ ) );
MUX2_X1 _10843_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_27 ), .Z(_03102_ ) );
MUX2_X1 _10844_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_27 ), .Z(_03103_ ) );
MUX2_X1 _10845_ ( .A(_03102_ ), .B(_03103_ ), .S(fanout_net_33 ), .Z(_03104_ ) );
OAI211_X1 _10846_ ( .A(fanout_net_37 ), .B(_03101_ ), .C1(_03104_ ), .C2(fanout_net_36 ), .ZN(_03105_ ) );
NAND2_X1 _10847_ ( .A1(_03096_ ), .A2(_03105_ ), .ZN(_03106_ ) );
OAI21_X4 _10848_ ( .A(_03106_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_03107_ ) );
AND2_X1 _10849_ ( .A1(_03087_ ), .A2(_03107_ ), .ZN(_03108_ ) );
XNOR2_X2 _10850_ ( .A(_03108_ ), .B(_02403_ ), .ZN(_03109_ ) );
NAND3_X1 _10851_ ( .A1(_03060_ ), .A2(_03085_ ), .A3(_03109_ ), .ZN(_03110_ ) );
NOR2_X2 _10852_ ( .A1(_03008_ ), .A2(_03110_ ), .ZN(_03111_ ) );
NAND3_X1 _10853_ ( .A1(_02919_ ), .A2(\EX_LS_result_reg [14] ), .A3(_02037_ ), .ZN(_03112_ ) );
BUF_X4 _10854_ ( .A(_02867_ ), .Z(_03113_ ) );
NOR2_X1 _10855_ ( .A1(_03021_ ), .A2(\myreg.Reg[11][14] ), .ZN(_03114_ ) );
OAI21_X1 _10856_ ( .A(fanout_net_33 ), .B1(fanout_net_27 ), .B2(\myreg.Reg[10][14] ), .ZN(_03115_ ) );
NOR2_X1 _10857_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[8][14] ), .ZN(_03116_ ) );
OAI21_X1 _10858_ ( .A(_02929_ ), .B1(_03021_ ), .B2(\myreg.Reg[9][14] ), .ZN(_03117_ ) );
OAI221_X1 _10859_ ( .A(_03113_ ), .B1(_03114_ ), .B2(_03115_ ), .C1(_03116_ ), .C2(_03117_ ), .ZN(_03118_ ) );
MUX2_X1 _10860_ ( .A(\myreg.Reg[12][14] ), .B(\myreg.Reg[13][14] ), .S(fanout_net_27 ), .Z(_03119_ ) );
MUX2_X1 _10861_ ( .A(\myreg.Reg[14][14] ), .B(\myreg.Reg[15][14] ), .S(fanout_net_27 ), .Z(_03120_ ) );
MUX2_X1 _10862_ ( .A(_03119_ ), .B(_03120_ ), .S(fanout_net_33 ), .Z(_03121_ ) );
OAI211_X1 _10863_ ( .A(fanout_net_37 ), .B(_03118_ ), .C1(_03121_ ), .C2(_02869_ ), .ZN(_03122_ ) );
OR2_X1 _10864_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[4][14] ), .ZN(_03123_ ) );
OAI211_X1 _10865_ ( .A(_03123_ ), .B(_02881_ ), .C1(_02983_ ), .C2(\myreg.Reg[5][14] ), .ZN(_03124_ ) );
OR2_X1 _10866_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[6][14] ), .ZN(_03125_ ) );
OAI211_X1 _10867_ ( .A(_03125_ ), .B(fanout_net_33 ), .C1(_02983_ ), .C2(\myreg.Reg[7][14] ), .ZN(_03126_ ) );
NAND3_X1 _10868_ ( .A1(_03124_ ), .A2(_03126_ ), .A3(fanout_net_36 ), .ZN(_03127_ ) );
MUX2_X1 _10869_ ( .A(\myreg.Reg[2][14] ), .B(\myreg.Reg[3][14] ), .S(fanout_net_27 ), .Z(_03128_ ) );
MUX2_X1 _10870_ ( .A(\myreg.Reg[0][14] ), .B(\myreg.Reg[1][14] ), .S(fanout_net_27 ), .Z(_03129_ ) );
MUX2_X1 _10871_ ( .A(_03128_ ), .B(_03129_ ), .S(_02929_ ), .Z(_03130_ ) );
OAI211_X1 _10872_ ( .A(_02890_ ), .B(_03127_ ), .C1(_03130_ ), .C2(fanout_net_36 ), .ZN(_03131_ ) );
NAND2_X1 _10873_ ( .A1(_03122_ ), .A2(_03131_ ), .ZN(_03132_ ) );
OAI21_X1 _10874_ ( .A(_03132_ ), .B1(_02926_ ), .B2(_02924_ ), .ZN(_03133_ ) );
AND2_X1 _10875_ ( .A1(_03112_ ), .A2(_03133_ ), .ZN(_03134_ ) );
INV_X1 _10876_ ( .A(_02332_ ), .ZN(_03135_ ) );
XNOR2_X1 _10877_ ( .A(_03134_ ), .B(_03135_ ), .ZN(_03136_ ) );
INV_X1 _10878_ ( .A(_03136_ ), .ZN(_03137_ ) );
INV_X1 _10879_ ( .A(\EX_LS_result_reg [15] ), .ZN(_03138_ ) );
OR3_X1 _10880_ ( .A1(_02910_ ), .A2(_03138_ ), .A3(_02897_ ), .ZN(_03139_ ) );
OR2_X1 _10881_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[0][15] ), .ZN(_03140_ ) );
BUF_X4 _10882_ ( .A(_02863_ ), .Z(_03141_ ) );
OAI211_X1 _10883_ ( .A(_03140_ ), .B(_02872_ ), .C1(_03141_ ), .C2(\myreg.Reg[1][15] ), .ZN(_03142_ ) );
OR2_X1 _10884_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[2][15] ), .ZN(_03143_ ) );
OAI211_X1 _10885_ ( .A(_03143_ ), .B(fanout_net_33 ), .C1(_02874_ ), .C2(\myreg.Reg[3][15] ), .ZN(_03144_ ) );
NAND3_X1 _10886_ ( .A1(_03142_ ), .A2(_03144_ ), .A3(_02868_ ), .ZN(_03145_ ) );
MUX2_X1 _10887_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_27 ), .Z(_03146_ ) );
MUX2_X1 _10888_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_27 ), .Z(_03147_ ) );
MUX2_X1 _10889_ ( .A(_03146_ ), .B(_03147_ ), .S(_02880_ ), .Z(_03148_ ) );
OAI211_X1 _10890_ ( .A(_03019_ ), .B(_03145_ ), .C1(_03148_ ), .C2(_03113_ ), .ZN(_03149_ ) );
OR2_X1 _10891_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[14][15] ), .ZN(_03150_ ) );
OAI211_X1 _10892_ ( .A(_03150_ ), .B(fanout_net_33 ), .C1(_02874_ ), .C2(\myreg.Reg[15][15] ), .ZN(_03151_ ) );
OR2_X1 _10893_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[12][15] ), .ZN(_03152_ ) );
BUF_X4 _10894_ ( .A(_02871_ ), .Z(_03153_ ) );
OAI211_X1 _10895_ ( .A(_03152_ ), .B(_03153_ ), .C1(_02874_ ), .C2(\myreg.Reg[13][15] ), .ZN(_03154_ ) );
NAND3_X1 _10896_ ( .A1(_03151_ ), .A2(_03154_ ), .A3(fanout_net_36 ), .ZN(_03155_ ) );
MUX2_X1 _10897_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_27 ), .Z(_03156_ ) );
MUX2_X1 _10898_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_27 ), .Z(_03157_ ) );
MUX2_X1 _10899_ ( .A(_03156_ ), .B(_03157_ ), .S(fanout_net_33 ), .Z(_03158_ ) );
OAI211_X1 _10900_ ( .A(fanout_net_37 ), .B(_03155_ ), .C1(_03158_ ), .C2(fanout_net_36 ), .ZN(_03159_ ) );
NAND2_X1 _10901_ ( .A1(_03149_ ), .A2(_03159_ ), .ZN(_03160_ ) );
OAI21_X4 _10902_ ( .A(_03160_ ), .B1(_02898_ ), .B2(_02911_ ), .ZN(_03161_ ) );
AND2_X1 _10903_ ( .A1(_03139_ ), .A2(_03161_ ), .ZN(_03162_ ) );
XNOR2_X1 _10904_ ( .A(_03162_ ), .B(_02309_ ), .ZN(_03163_ ) );
NOR2_X1 _10905_ ( .A1(_03137_ ), .A2(_03163_ ), .ZN(_03164_ ) );
INV_X1 _10906_ ( .A(\EX_LS_result_reg [12] ), .ZN(_03165_ ) );
OR3_X1 _10907_ ( .A1(_02911_ ), .A2(_03165_ ), .A3(_02898_ ), .ZN(_03166_ ) );
OR2_X1 _10908_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[0][12] ), .ZN(_03167_ ) );
OAI211_X1 _10909_ ( .A(_03167_ ), .B(_02881_ ), .C1(_02983_ ), .C2(\myreg.Reg[1][12] ), .ZN(_03168_ ) );
OR2_X1 _10910_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[2][12] ), .ZN(_03169_ ) );
OAI211_X1 _10911_ ( .A(_03169_ ), .B(fanout_net_33 ), .C1(_03021_ ), .C2(\myreg.Reg[3][12] ), .ZN(_03170_ ) );
NAND3_X1 _10912_ ( .A1(_03168_ ), .A2(_03170_ ), .A3(_03113_ ), .ZN(_03171_ ) );
MUX2_X1 _10913_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_27 ), .Z(_03172_ ) );
MUX2_X1 _10914_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_27 ), .Z(_03173_ ) );
MUX2_X1 _10915_ ( .A(_03172_ ), .B(_03173_ ), .S(_02929_ ), .Z(_03174_ ) );
OAI211_X1 _10916_ ( .A(_03019_ ), .B(_03171_ ), .C1(_03174_ ), .C2(_02869_ ), .ZN(_03175_ ) );
OR2_X1 _10917_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[14][12] ), .ZN(_03176_ ) );
OAI211_X1 _10918_ ( .A(_03176_ ), .B(fanout_net_33 ), .C1(_02983_ ), .C2(\myreg.Reg[15][12] ), .ZN(_03177_ ) );
OR2_X1 _10919_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[12][12] ), .ZN(_03178_ ) );
OAI211_X1 _10920_ ( .A(_03178_ ), .B(_02929_ ), .C1(_03021_ ), .C2(\myreg.Reg[13][12] ), .ZN(_03179_ ) );
NAND3_X1 _10921_ ( .A1(_03177_ ), .A2(_03179_ ), .A3(fanout_net_36 ), .ZN(_03180_ ) );
MUX2_X1 _10922_ ( .A(\myreg.Reg[8][12] ), .B(\myreg.Reg[9][12] ), .S(fanout_net_27 ), .Z(_03181_ ) );
MUX2_X1 _10923_ ( .A(\myreg.Reg[10][12] ), .B(\myreg.Reg[11][12] ), .S(fanout_net_27 ), .Z(_03182_ ) );
MUX2_X1 _10924_ ( .A(_03181_ ), .B(_03182_ ), .S(fanout_net_34 ), .Z(_03183_ ) );
OAI211_X1 _10925_ ( .A(fanout_net_37 ), .B(_03180_ ), .C1(_03183_ ), .C2(fanout_net_36 ), .ZN(_03184_ ) );
NAND2_X1 _10926_ ( .A1(_03175_ ), .A2(_03184_ ), .ZN(_03185_ ) );
OAI21_X1 _10927_ ( .A(_03185_ ), .B1(_02926_ ), .B2(_02924_ ), .ZN(_03186_ ) );
AND2_X1 _10928_ ( .A1(_03166_ ), .A2(_03186_ ), .ZN(_03187_ ) );
INV_X1 _10929_ ( .A(_02380_ ), .ZN(_03188_ ) );
XNOR2_X1 _10930_ ( .A(_03187_ ), .B(_03188_ ), .ZN(_03189_ ) );
INV_X1 _10931_ ( .A(\EX_LS_result_reg [13] ), .ZN(_03190_ ) );
OR3_X1 _10932_ ( .A1(_02924_ ), .A2(_03190_ ), .A3(_02926_ ), .ZN(_03191_ ) );
OR2_X1 _10933_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[0][13] ), .ZN(_03192_ ) );
OAI211_X1 _10934_ ( .A(_03192_ ), .B(_02873_ ), .C1(_02941_ ), .C2(\myreg.Reg[1][13] ), .ZN(_03193_ ) );
OR2_X1 _10935_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[2][13] ), .ZN(_03194_ ) );
OAI211_X1 _10936_ ( .A(_03194_ ), .B(fanout_net_34 ), .C1(_02875_ ), .C2(\myreg.Reg[3][13] ), .ZN(_03195_ ) );
NAND3_X1 _10937_ ( .A1(_03193_ ), .A2(_03195_ ), .A3(_02869_ ), .ZN(_03196_ ) );
MUX2_X1 _10938_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_28 ), .Z(_03197_ ) );
MUX2_X1 _10939_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_28 ), .Z(_03198_ ) );
MUX2_X1 _10940_ ( .A(_03197_ ), .B(_03198_ ), .S(_02873_ ), .Z(_03199_ ) );
OAI211_X1 _10941_ ( .A(_02890_ ), .B(_03196_ ), .C1(_03199_ ), .C2(_02883_ ), .ZN(_03200_ ) );
OR2_X1 _10942_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[14][13] ), .ZN(_03201_ ) );
OAI211_X1 _10943_ ( .A(_03201_ ), .B(fanout_net_34 ), .C1(_02875_ ), .C2(\myreg.Reg[15][13] ), .ZN(_03202_ ) );
OR2_X1 _10944_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[12][13] ), .ZN(_03203_ ) );
OAI211_X1 _10945_ ( .A(_03203_ ), .B(_02873_ ), .C1(_02875_ ), .C2(\myreg.Reg[13][13] ), .ZN(_03204_ ) );
NAND3_X1 _10946_ ( .A1(_03202_ ), .A2(_03204_ ), .A3(fanout_net_36 ), .ZN(_03205_ ) );
MUX2_X1 _10947_ ( .A(\myreg.Reg[8][13] ), .B(\myreg.Reg[9][13] ), .S(fanout_net_28 ), .Z(_03206_ ) );
MUX2_X1 _10948_ ( .A(\myreg.Reg[10][13] ), .B(\myreg.Reg[11][13] ), .S(fanout_net_28 ), .Z(_03207_ ) );
MUX2_X1 _10949_ ( .A(_03206_ ), .B(_03207_ ), .S(fanout_net_34 ), .Z(_03208_ ) );
OAI211_X1 _10950_ ( .A(fanout_net_37 ), .B(_03205_ ), .C1(_03208_ ), .C2(fanout_net_36 ), .ZN(_03209_ ) );
NAND2_X1 _10951_ ( .A1(_03200_ ), .A2(_03209_ ), .ZN(_03210_ ) );
OAI21_X2 _10952_ ( .A(_03210_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_03211_ ) );
AND2_X1 _10953_ ( .A1(_03191_ ), .A2(_03211_ ), .ZN(_03212_ ) );
NAND2_X2 _10954_ ( .A1(_02354_ ), .A2(_02356_ ), .ZN(_03213_ ) );
INV_X1 _10955_ ( .A(_03213_ ), .ZN(_03214_ ) );
XNOR2_X2 _10956_ ( .A(_03212_ ), .B(_03214_ ), .ZN(_03215_ ) );
AND2_X1 _10957_ ( .A1(_03189_ ), .A2(_03215_ ), .ZN(_03216_ ) );
AND2_X1 _10958_ ( .A1(_03164_ ), .A2(_03216_ ), .ZN(_03217_ ) );
INV_X1 _10959_ ( .A(\EX_LS_result_reg [11] ), .ZN(_03218_ ) );
OR3_X1 _10960_ ( .A1(_02911_ ), .A2(_03218_ ), .A3(_02897_ ), .ZN(_03219_ ) );
OR2_X1 _10961_ ( .A1(_02863_ ), .A2(\myreg.Reg[3][11] ), .ZN(_03220_ ) );
OAI211_X1 _10962_ ( .A(_03220_ ), .B(fanout_net_34 ), .C1(fanout_net_28 ), .C2(\myreg.Reg[2][11] ), .ZN(_03221_ ) );
OR2_X1 _10963_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[0][11] ), .ZN(_03222_ ) );
OAI211_X1 _10964_ ( .A(_03222_ ), .B(_02929_ ), .C1(_02864_ ), .C2(\myreg.Reg[1][11] ), .ZN(_03223_ ) );
NAND3_X1 _10965_ ( .A1(_03221_ ), .A2(_02868_ ), .A3(_03223_ ), .ZN(_03224_ ) );
MUX2_X1 _10966_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_28 ), .Z(_03225_ ) );
MUX2_X1 _10967_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_28 ), .Z(_03226_ ) );
MUX2_X1 _10968_ ( .A(_03225_ ), .B(_03226_ ), .S(_02872_ ), .Z(_03227_ ) );
OAI211_X1 _10969_ ( .A(_03019_ ), .B(_03224_ ), .C1(_03227_ ), .C2(_02869_ ), .ZN(_03228_ ) );
OR2_X1 _10970_ ( .A1(_02863_ ), .A2(\myreg.Reg[13][11] ), .ZN(_03229_ ) );
OAI211_X1 _10971_ ( .A(_03229_ ), .B(_02929_ ), .C1(fanout_net_28 ), .C2(\myreg.Reg[12][11] ), .ZN(_03230_ ) );
OR2_X1 _10972_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[14][11] ), .ZN(_03231_ ) );
OAI211_X1 _10973_ ( .A(_03231_ ), .B(fanout_net_34 ), .C1(_02864_ ), .C2(\myreg.Reg[15][11] ), .ZN(_03232_ ) );
NAND3_X1 _10974_ ( .A1(_03230_ ), .A2(fanout_net_36 ), .A3(_03232_ ), .ZN(_03233_ ) );
MUX2_X1 _10975_ ( .A(\myreg.Reg[8][11] ), .B(\myreg.Reg[9][11] ), .S(fanout_net_28 ), .Z(_03234_ ) );
MUX2_X1 _10976_ ( .A(\myreg.Reg[10][11] ), .B(\myreg.Reg[11][11] ), .S(fanout_net_28 ), .Z(_03235_ ) );
MUX2_X1 _10977_ ( .A(_03234_ ), .B(_03235_ ), .S(fanout_net_34 ), .Z(_03236_ ) );
OAI211_X1 _10978_ ( .A(fanout_net_37 ), .B(_03233_ ), .C1(_03236_ ), .C2(fanout_net_36 ), .ZN(_03237_ ) );
NAND2_X1 _10979_ ( .A1(_03228_ ), .A2(_03237_ ), .ZN(_03238_ ) );
OAI21_X1 _10980_ ( .A(_03238_ ), .B1(_02926_ ), .B2(_02924_ ), .ZN(_03239_ ) );
AND2_X1 _10981_ ( .A1(_03219_ ), .A2(_03239_ ), .ZN(_03240_ ) );
INV_X1 _10982_ ( .A(_02272_ ), .ZN(_03241_ ) );
XNOR2_X2 _10983_ ( .A(_03240_ ), .B(_03241_ ), .ZN(_03242_ ) );
INV_X1 _10984_ ( .A(\EX_LS_result_reg [10] ), .ZN(_03243_ ) );
OR3_X1 _10985_ ( .A1(_02911_ ), .A2(_03243_ ), .A3(_02898_ ), .ZN(_03244_ ) );
NOR2_X1 _10986_ ( .A1(_03021_ ), .A2(\myreg.Reg[11][10] ), .ZN(_03245_ ) );
OAI21_X1 _10987_ ( .A(fanout_net_34 ), .B1(fanout_net_28 ), .B2(\myreg.Reg[10][10] ), .ZN(_03246_ ) );
NOR2_X1 _10988_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[8][10] ), .ZN(_03247_ ) );
OAI21_X1 _10989_ ( .A(_02881_ ), .B1(_03021_ ), .B2(\myreg.Reg[9][10] ), .ZN(_03248_ ) );
OAI221_X1 _10990_ ( .A(_03113_ ), .B1(_03245_ ), .B2(_03246_ ), .C1(_03247_ ), .C2(_03248_ ), .ZN(_03249_ ) );
MUX2_X1 _10991_ ( .A(\myreg.Reg[12][10] ), .B(\myreg.Reg[13][10] ), .S(fanout_net_28 ), .Z(_03250_ ) );
MUX2_X1 _10992_ ( .A(\myreg.Reg[14][10] ), .B(\myreg.Reg[15][10] ), .S(fanout_net_28 ), .Z(_03251_ ) );
MUX2_X1 _10993_ ( .A(_03250_ ), .B(_03251_ ), .S(fanout_net_34 ), .Z(_03252_ ) );
OAI211_X1 _10994_ ( .A(fanout_net_37 ), .B(_03249_ ), .C1(_03252_ ), .C2(_02883_ ), .ZN(_03253_ ) );
OR2_X1 _10995_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[4][10] ), .ZN(_03254_ ) );
OAI211_X1 _10996_ ( .A(_03254_ ), .B(_02881_ ), .C1(_02983_ ), .C2(\myreg.Reg[5][10] ), .ZN(_03255_ ) );
OR2_X1 _10997_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[6][10] ), .ZN(_03256_ ) );
OAI211_X1 _10998_ ( .A(_03256_ ), .B(fanout_net_34 ), .C1(_02983_ ), .C2(\myreg.Reg[7][10] ), .ZN(_03257_ ) );
NAND3_X1 _10999_ ( .A1(_03255_ ), .A2(_03257_ ), .A3(fanout_net_36 ), .ZN(_03258_ ) );
MUX2_X1 _11000_ ( .A(\myreg.Reg[2][10] ), .B(\myreg.Reg[3][10] ), .S(fanout_net_28 ), .Z(_03259_ ) );
MUX2_X1 _11001_ ( .A(\myreg.Reg[0][10] ), .B(\myreg.Reg[1][10] ), .S(fanout_net_28 ), .Z(_03260_ ) );
MUX2_X1 _11002_ ( .A(_03259_ ), .B(_03260_ ), .S(_02929_ ), .Z(_03261_ ) );
OAI211_X1 _11003_ ( .A(_02890_ ), .B(_03258_ ), .C1(_03261_ ), .C2(fanout_net_36 ), .ZN(_03262_ ) );
NAND2_X1 _11004_ ( .A1(_03253_ ), .A2(_03262_ ), .ZN(_03263_ ) );
OAI21_X1 _11005_ ( .A(_03263_ ), .B1(_02899_ ), .B2(_02924_ ), .ZN(_03264_ ) );
AND2_X1 _11006_ ( .A1(_03244_ ), .A2(_03264_ ), .ZN(_03265_ ) );
INV_X1 _11007_ ( .A(_02249_ ), .ZN(_03266_ ) );
XNOR2_X1 _11008_ ( .A(_03265_ ), .B(_03266_ ), .ZN(_03267_ ) );
AND2_X2 _11009_ ( .A1(_03242_ ), .A2(_03267_ ), .ZN(_03268_ ) );
INV_X1 _11010_ ( .A(\EX_LS_result_reg [9] ), .ZN(_03269_ ) );
OR3_X1 _11011_ ( .A1(_02911_ ), .A2(_03269_ ), .A3(_02898_ ), .ZN(_03270_ ) );
OR2_X1 _11012_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[0][9] ), .ZN(_03271_ ) );
OAI211_X1 _11013_ ( .A(_03271_ ), .B(_02881_ ), .C1(_02983_ ), .C2(\myreg.Reg[1][9] ), .ZN(_03272_ ) );
OR2_X1 _11014_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[2][9] ), .ZN(_03273_ ) );
OAI211_X1 _11015_ ( .A(_03273_ ), .B(fanout_net_34 ), .C1(_02983_ ), .C2(\myreg.Reg[3][9] ), .ZN(_03274_ ) );
NAND3_X1 _11016_ ( .A1(_03272_ ), .A2(_03274_ ), .A3(_03113_ ), .ZN(_03275_ ) );
MUX2_X1 _11017_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_28 ), .Z(_03276_ ) );
MUX2_X1 _11018_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_28 ), .Z(_03277_ ) );
MUX2_X1 _11019_ ( .A(_03276_ ), .B(_03277_ ), .S(_02929_ ), .Z(_03278_ ) );
OAI211_X1 _11020_ ( .A(_02890_ ), .B(_03275_ ), .C1(_03278_ ), .C2(_02869_ ), .ZN(_03279_ ) );
OR2_X1 _11021_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[14][9] ), .ZN(_03280_ ) );
OAI211_X1 _11022_ ( .A(_03280_ ), .B(fanout_net_34 ), .C1(_02983_ ), .C2(\myreg.Reg[15][9] ), .ZN(_03281_ ) );
OR2_X1 _11023_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[12][9] ), .ZN(_03282_ ) );
OAI211_X1 _11024_ ( .A(_03282_ ), .B(_02881_ ), .C1(_03021_ ), .C2(\myreg.Reg[13][9] ), .ZN(_03283_ ) );
NAND3_X1 _11025_ ( .A1(_03281_ ), .A2(_03283_ ), .A3(fanout_net_36 ), .ZN(_03284_ ) );
MUX2_X1 _11026_ ( .A(\myreg.Reg[8][9] ), .B(\myreg.Reg[9][9] ), .S(fanout_net_28 ), .Z(_03285_ ) );
MUX2_X1 _11027_ ( .A(\myreg.Reg[10][9] ), .B(\myreg.Reg[11][9] ), .S(fanout_net_29 ), .Z(_03286_ ) );
MUX2_X1 _11028_ ( .A(_03285_ ), .B(_03286_ ), .S(fanout_net_34 ), .Z(_03287_ ) );
OAI211_X1 _11029_ ( .A(fanout_net_37 ), .B(_03284_ ), .C1(_03287_ ), .C2(fanout_net_36 ), .ZN(_03288_ ) );
NAND2_X1 _11030_ ( .A1(_03279_ ), .A2(_03288_ ), .ZN(_03289_ ) );
OAI21_X1 _11031_ ( .A(_03289_ ), .B1(_02926_ ), .B2(_02924_ ), .ZN(_03290_ ) );
AND2_X1 _11032_ ( .A1(_03270_ ), .A2(_03290_ ), .ZN(_03291_ ) );
INV_X1 _11033_ ( .A(_02225_ ), .ZN(_03292_ ) );
XNOR2_X2 _11034_ ( .A(_03291_ ), .B(_03292_ ), .ZN(_03293_ ) );
OR2_X1 _11035_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][8] ), .ZN(_03294_ ) );
BUF_X4 _11036_ ( .A(_03021_ ), .Z(_03295_ ) );
OAI211_X1 _11037_ ( .A(_03294_ ), .B(_02980_ ), .C1(_03295_ ), .C2(\myreg.Reg[1][8] ), .ZN(_03296_ ) );
OR2_X1 _11038_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[2][8] ), .ZN(_03297_ ) );
OAI211_X1 _11039_ ( .A(_03297_ ), .B(fanout_net_34 ), .C1(_03295_ ), .C2(\myreg.Reg[3][8] ), .ZN(_03298_ ) );
NAND3_X1 _11040_ ( .A1(_03296_ ), .A2(_03298_ ), .A3(_02883_ ), .ZN(_03299_ ) );
MUX2_X1 _11041_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_29 ), .Z(_03300_ ) );
MUX2_X1 _11042_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_29 ), .Z(_03301_ ) );
MUX2_X1 _11043_ ( .A(_03300_ ), .B(_03301_ ), .S(_02930_ ), .Z(_03302_ ) );
OAI211_X1 _11044_ ( .A(_02996_ ), .B(_03299_ ), .C1(_03302_ ), .C2(_02938_ ), .ZN(_03303_ ) );
OR2_X1 _11045_ ( .A1(_03021_ ), .A2(\myreg.Reg[13][8] ), .ZN(_03304_ ) );
OAI211_X1 _11046_ ( .A(_03304_ ), .B(_02930_ ), .C1(fanout_net_29 ), .C2(\myreg.Reg[12][8] ), .ZN(_03305_ ) );
OR2_X1 _11047_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[14][8] ), .ZN(_03306_ ) );
OAI211_X1 _11048_ ( .A(_03306_ ), .B(fanout_net_34 ), .C1(_02941_ ), .C2(\myreg.Reg[15][8] ), .ZN(_03307_ ) );
NAND3_X1 _11049_ ( .A1(_03305_ ), .A2(fanout_net_36 ), .A3(_03307_ ), .ZN(_03308_ ) );
MUX2_X1 _11050_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_29 ), .Z(_03309_ ) );
MUX2_X1 _11051_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_29 ), .Z(_03310_ ) );
MUX2_X1 _11052_ ( .A(_03309_ ), .B(_03310_ ), .S(fanout_net_34 ), .Z(_03311_ ) );
OAI211_X1 _11053_ ( .A(fanout_net_37 ), .B(_03308_ ), .C1(_03311_ ), .C2(fanout_net_36 ), .ZN(_03312_ ) );
AOI21_X1 _11054_ ( .A(_03061_ ), .B1(_03303_ ), .B2(_03312_ ), .ZN(_03313_ ) );
INV_X1 _11055_ ( .A(\EX_LS_result_reg [8] ), .ZN(_03314_ ) );
NOR3_X1 _11056_ ( .A1(_02912_ ), .A2(_03314_ ), .A3(_02926_ ), .ZN(_03315_ ) );
NOR2_X1 _11057_ ( .A1(_03313_ ), .A2(_03315_ ), .ZN(_03316_ ) );
INV_X1 _11058_ ( .A(_02202_ ), .ZN(_03317_ ) );
XNOR2_X1 _11059_ ( .A(_03316_ ), .B(_03317_ ), .ZN(_03318_ ) );
AND3_X1 _11060_ ( .A1(_03268_ ), .A2(_03293_ ), .A3(_03318_ ), .ZN(_03319_ ) );
NAND3_X1 _11061_ ( .A1(_02919_ ), .A2(\EX_LS_result_reg [7] ), .A3(_02012_ ), .ZN(_03320_ ) );
NOR2_X1 _11062_ ( .A1(_02862_ ), .A2(\myreg.Reg[11][7] ), .ZN(_03321_ ) );
OAI21_X1 _11063_ ( .A(fanout_net_34 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[10][7] ), .ZN(_03322_ ) );
NOR2_X1 _11064_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][7] ), .ZN(_03323_ ) );
OAI21_X1 _11065_ ( .A(_02871_ ), .B1(_02862_ ), .B2(\myreg.Reg[9][7] ), .ZN(_03324_ ) );
OAI221_X1 _11066_ ( .A(_02867_ ), .B1(_03321_ ), .B2(_03322_ ), .C1(_03323_ ), .C2(_03324_ ), .ZN(_03325_ ) );
MUX2_X1 _11067_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_29 ), .Z(_03326_ ) );
MUX2_X1 _11068_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_29 ), .Z(_03327_ ) );
MUX2_X1 _11069_ ( .A(_03326_ ), .B(_03327_ ), .S(fanout_net_34 ), .Z(_03328_ ) );
OAI211_X1 _11070_ ( .A(fanout_net_37 ), .B(_03325_ ), .C1(_03328_ ), .C2(_02867_ ), .ZN(_03329_ ) );
OR2_X1 _11071_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[4][7] ), .ZN(_03330_ ) );
OAI211_X1 _11072_ ( .A(_03330_ ), .B(_02871_ ), .C1(_02862_ ), .C2(\myreg.Reg[5][7] ), .ZN(_03331_ ) );
OR2_X1 _11073_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[6][7] ), .ZN(_03332_ ) );
OAI211_X1 _11074_ ( .A(_03332_ ), .B(fanout_net_34 ), .C1(_02862_ ), .C2(\myreg.Reg[7][7] ), .ZN(_03333_ ) );
NAND3_X1 _11075_ ( .A1(_03331_ ), .A2(_03333_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03334_ ) );
MUX2_X1 _11076_ ( .A(\myreg.Reg[2][7] ), .B(\myreg.Reg[3][7] ), .S(fanout_net_29 ), .Z(_03335_ ) );
MUX2_X1 _11077_ ( .A(\myreg.Reg[0][7] ), .B(\myreg.Reg[1][7] ), .S(fanout_net_29 ), .Z(_03336_ ) );
MUX2_X1 _11078_ ( .A(_03335_ ), .B(_03336_ ), .S(_02871_ ), .Z(_03337_ ) );
OAI211_X1 _11079_ ( .A(_02889_ ), .B(_03334_ ), .C1(_03337_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03338_ ) );
NAND2_X1 _11080_ ( .A1(_03329_ ), .A2(_03338_ ), .ZN(_03339_ ) );
OAI21_X1 _11081_ ( .A(_03339_ ), .B1(_02896_ ), .B2(_02909_ ), .ZN(_03340_ ) );
AND2_X2 _11082_ ( .A1(_03320_ ), .A2(_03340_ ), .ZN(_03341_ ) );
INV_X2 _11083_ ( .A(_02149_ ), .ZN(_03342_ ) );
XNOR2_X2 _11084_ ( .A(_03341_ ), .B(_03342_ ), .ZN(_03343_ ) );
INV_X1 _11085_ ( .A(_02171_ ), .ZN(_03344_ ) );
INV_X1 _11086_ ( .A(\EX_LS_dest_reg [3] ), .ZN(_03345_ ) );
INV_X1 _11087_ ( .A(\ID_EX_rs2 [1] ), .ZN(_03346_ ) );
AOI22_X1 _11088_ ( .A1(_03345_ ), .A2(\ID_EX_rs2 [3] ), .B1(_03346_ ), .B2(\EX_LS_dest_reg [1] ), .ZN(_03347_ ) );
NAND3_X1 _11089_ ( .A1(_02908_ ), .A2(_02904_ ), .A3(_03347_ ), .ZN(_03348_ ) );
NOR2_X1 _11090_ ( .A1(_03345_ ), .A2(\ID_EX_rs2 [3] ), .ZN(_03349_ ) );
NOR3_X1 _11091_ ( .A1(_03348_ ), .A2(_02896_ ), .A3(_03349_ ), .ZN(_03350_ ) );
NAND3_X1 _11092_ ( .A1(_02012_ ), .A2(_03350_ ), .A3(_02902_ ), .ZN(_03351_ ) );
OAI21_X1 _11093_ ( .A(_02907_ ), .B1(\EX_LS_dest_reg [1] ), .B2(_03346_ ), .ZN(_03352_ ) );
OR3_X4 _11094_ ( .A1(_03351_ ), .A2(\EX_LS_result_reg [6] ), .A3(_03352_ ), .ZN(_03353_ ) );
OR2_X1 _11095_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[4][6] ), .ZN(_03354_ ) );
OAI211_X1 _11096_ ( .A(_03354_ ), .B(_02872_ ), .C1(_03141_ ), .C2(\myreg.Reg[5][6] ), .ZN(_03355_ ) );
OR2_X1 _11097_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[6][6] ), .ZN(_03356_ ) );
OAI211_X1 _11098_ ( .A(_03356_ ), .B(fanout_net_34 ), .C1(_03141_ ), .C2(\myreg.Reg[7][6] ), .ZN(_03357_ ) );
NAND3_X1 _11099_ ( .A1(_03355_ ), .A2(_03357_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03358_ ) );
MUX2_X1 _11100_ ( .A(\myreg.Reg[2][6] ), .B(\myreg.Reg[3][6] ), .S(fanout_net_29 ), .Z(_03359_ ) );
MUX2_X1 _11101_ ( .A(\myreg.Reg[0][6] ), .B(\myreg.Reg[1][6] ), .S(fanout_net_29 ), .Z(_03360_ ) );
MUX2_X1 _11102_ ( .A(_03359_ ), .B(_03360_ ), .S(_03153_ ), .Z(_03361_ ) );
OAI211_X1 _11103_ ( .A(_03019_ ), .B(_03358_ ), .C1(_03361_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03362_ ) );
NOR2_X1 _11104_ ( .A1(_02982_ ), .A2(\myreg.Reg[11][6] ), .ZN(_03363_ ) );
OAI21_X1 _11105_ ( .A(fanout_net_34 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[10][6] ), .ZN(_03364_ ) );
NOR2_X1 _11106_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][6] ), .ZN(_03365_ ) );
OAI21_X1 _11107_ ( .A(_03153_ ), .B1(_02982_ ), .B2(\myreg.Reg[9][6] ), .ZN(_03366_ ) );
OAI221_X1 _11108_ ( .A(_02867_ ), .B1(_03363_ ), .B2(_03364_ ), .C1(_03365_ ), .C2(_03366_ ), .ZN(_03367_ ) );
MUX2_X1 _11109_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(fanout_net_29 ), .Z(_03368_ ) );
MUX2_X1 _11110_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(fanout_net_29 ), .Z(_03369_ ) );
MUX2_X1 _11111_ ( .A(_03368_ ), .B(_03369_ ), .S(fanout_net_34 ), .Z(_03370_ ) );
OAI211_X1 _11112_ ( .A(fanout_net_37 ), .B(_03367_ ), .C1(_03370_ ), .C2(_03113_ ), .ZN(_03371_ ) );
OAI211_X1 _11113_ ( .A(_03362_ ), .B(_03371_ ), .C1(_03351_ ), .C2(_03352_ ), .ZN(_03372_ ) );
NAND2_X1 _11114_ ( .A1(_03353_ ), .A2(_03372_ ), .ZN(_03373_ ) );
XNOR2_X1 _11115_ ( .A(_03344_ ), .B(_03373_ ), .ZN(_03374_ ) );
AND2_X1 _11116_ ( .A1(_03343_ ), .A2(_03374_ ), .ZN(_03375_ ) );
NAND3_X1 _11117_ ( .A1(_02919_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02037_ ), .ZN(_03376_ ) );
NOR2_X1 _11118_ ( .A1(_02982_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03377_ ) );
OAI21_X1 _11119_ ( .A(fanout_net_34 ), .B1(fanout_net_29 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03378_ ) );
NOR2_X1 _11120_ ( .A1(fanout_net_29 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03379_ ) );
OAI21_X1 _11121_ ( .A(_02880_ ), .B1(_02982_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03380_ ) );
OAI221_X1 _11122_ ( .A(_02867_ ), .B1(_03377_ ), .B2(_03378_ ), .C1(_03379_ ), .C2(_03380_ ), .ZN(_03381_ ) );
MUX2_X1 _11123_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_03382_ ) );
MUX2_X1 _11124_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_03383_ ) );
MUX2_X1 _11125_ ( .A(_03382_ ), .B(_03383_ ), .S(fanout_net_34 ), .Z(_03384_ ) );
OAI211_X1 _11126_ ( .A(fanout_net_37 ), .B(_03381_ ), .C1(_03384_ ), .C2(_03113_ ), .ZN(_03385_ ) );
OR2_X1 _11127_ ( .A1(fanout_net_29 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03386_ ) );
OAI211_X1 _11128_ ( .A(_03386_ ), .B(_03153_ ), .C1(_02874_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03387_ ) );
OR2_X1 _11129_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03388_ ) );
OAI211_X1 _11130_ ( .A(_03388_ ), .B(fanout_net_34 ), .C1(_02874_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03389_ ) );
NAND3_X1 _11131_ ( .A1(_03387_ ), .A2(_03389_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03390_ ) );
MUX2_X1 _11132_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03391_ ) );
MUX2_X1 _11133_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03392_ ) );
MUX2_X1 _11134_ ( .A(_03391_ ), .B(_03392_ ), .S(_02880_ ), .Z(_03393_ ) );
OAI211_X1 _11135_ ( .A(_03019_ ), .B(_03390_ ), .C1(_03393_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03394_ ) );
NAND2_X1 _11136_ ( .A1(_03385_ ), .A2(_03394_ ), .ZN(_03395_ ) );
OAI21_X2 _11137_ ( .A(_03395_ ), .B1(_02898_ ), .B2(_02911_ ), .ZN(_03396_ ) );
AND2_X1 _11138_ ( .A1(_03376_ ), .A2(_03396_ ), .ZN(_03397_ ) );
XNOR2_X1 _11139_ ( .A(_03397_ ), .B(_02096_ ), .ZN(_03398_ ) );
NAND2_X1 _11140_ ( .A1(_03061_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_03399_ ) );
OR2_X1 _11141_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[0][4] ), .ZN(_03400_ ) );
OAI211_X1 _11142_ ( .A(_03400_ ), .B(_02872_ ), .C1(_03141_ ), .C2(\myreg.Reg[1][4] ), .ZN(_03401_ ) );
OR2_X1 _11143_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[2][4] ), .ZN(_03402_ ) );
OAI211_X1 _11144_ ( .A(_03402_ ), .B(fanout_net_34 ), .C1(_02874_ ), .C2(\myreg.Reg[3][4] ), .ZN(_03403_ ) );
NAND3_X1 _11145_ ( .A1(_03401_ ), .A2(_03403_ ), .A3(_02868_ ), .ZN(_03404_ ) );
MUX2_X1 _11146_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_30 ), .Z(_03405_ ) );
MUX2_X1 _11147_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_30 ), .Z(_03406_ ) );
MUX2_X1 _11148_ ( .A(_03405_ ), .B(_03406_ ), .S(_03153_ ), .Z(_03407_ ) );
OAI211_X1 _11149_ ( .A(_03019_ ), .B(_03404_ ), .C1(_03407_ ), .C2(_03113_ ), .ZN(_03408_ ) );
OR2_X1 _11150_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[14][4] ), .ZN(_03409_ ) );
OAI211_X1 _11151_ ( .A(_03409_ ), .B(fanout_net_34 ), .C1(_03141_ ), .C2(\myreg.Reg[15][4] ), .ZN(_03410_ ) );
OR2_X1 _11152_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[12][4] ), .ZN(_03411_ ) );
OAI211_X1 _11153_ ( .A(_03411_ ), .B(_03153_ ), .C1(_02874_ ), .C2(\myreg.Reg[13][4] ), .ZN(_03412_ ) );
NAND3_X1 _11154_ ( .A1(_03410_ ), .A2(_03412_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03413_ ) );
MUX2_X1 _11155_ ( .A(\myreg.Reg[8][4] ), .B(\myreg.Reg[9][4] ), .S(fanout_net_30 ), .Z(_03414_ ) );
MUX2_X1 _11156_ ( .A(\myreg.Reg[10][4] ), .B(\myreg.Reg[11][4] ), .S(fanout_net_30 ), .Z(_03415_ ) );
MUX2_X1 _11157_ ( .A(_03414_ ), .B(_03415_ ), .S(fanout_net_34 ), .Z(_03416_ ) );
OAI211_X1 _11158_ ( .A(fanout_net_37 ), .B(_03413_ ), .C1(_03416_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03417_ ) );
NAND2_X1 _11159_ ( .A1(_03408_ ), .A2(_03417_ ), .ZN(_03418_ ) );
OAI21_X2 _11160_ ( .A(_03418_ ), .B1(_02898_ ), .B2(_02911_ ), .ZN(_03419_ ) );
AND2_X1 _11161_ ( .A1(_03399_ ), .A2(_03419_ ), .ZN(_03420_ ) );
XNOR2_X2 _11162_ ( .A(_03420_ ), .B(_02123_ ), .ZN(_03421_ ) );
AND2_X1 _11163_ ( .A1(_03398_ ), .A2(_03421_ ), .ZN(_03422_ ) );
AND2_X2 _11164_ ( .A1(_03375_ ), .A2(_03422_ ), .ZN(_03423_ ) );
AND3_X1 _11165_ ( .A1(_03217_ ), .A2(_03319_ ), .A3(_03423_ ), .ZN(_03424_ ) );
OR2_X1 _11166_ ( .A1(_03351_ ), .A2(_03352_ ), .ZN(_03425_ ) );
OR2_X1 _11167_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03426_ ) );
BUF_X4 _11168_ ( .A(_03295_ ), .Z(_03427_ ) );
OAI211_X1 _11169_ ( .A(_03426_ ), .B(_02993_ ), .C1(_03427_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03428_ ) );
NAND2_X1 _11170_ ( .A1(_02412_ ), .A2(fanout_net_30 ), .ZN(_03429_ ) );
OAI211_X1 _11171_ ( .A(_03429_ ), .B(fanout_net_34 ), .C1(fanout_net_30 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03430_ ) );
BUF_X4 _11172_ ( .A(_02883_ ), .Z(_03431_ ) );
NAND3_X1 _11173_ ( .A1(_03428_ ), .A2(_03430_ ), .A3(_03431_ ), .ZN(_03432_ ) );
MUX2_X1 _11174_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03433_ ) );
MUX2_X1 _11175_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03434_ ) );
MUX2_X1 _11176_ ( .A(_03433_ ), .B(_03434_ ), .S(_02993_ ), .Z(_03435_ ) );
BUF_X4 _11177_ ( .A(_02938_ ), .Z(_03436_ ) );
OAI211_X1 _11178_ ( .A(fanout_net_37 ), .B(_03432_ ), .C1(_03435_ ), .C2(_03436_ ), .ZN(_03437_ ) );
OR2_X1 _11179_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03438_ ) );
OAI211_X1 _11180_ ( .A(_03438_ ), .B(_02993_ ), .C1(_03427_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03439_ ) );
NAND2_X1 _11181_ ( .A1(_02422_ ), .A2(fanout_net_30 ), .ZN(_03440_ ) );
OAI211_X1 _11182_ ( .A(_03440_ ), .B(fanout_net_34 ), .C1(fanout_net_30 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03441_ ) );
NAND3_X1 _11183_ ( .A1(_03439_ ), .A2(_03441_ ), .A3(_03431_ ), .ZN(_03442_ ) );
MUX2_X1 _11184_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03443_ ) );
MUX2_X1 _11185_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03444_ ) );
MUX2_X1 _11186_ ( .A(_03443_ ), .B(_03444_ ), .S(_02993_ ), .Z(_03445_ ) );
OAI211_X1 _11187_ ( .A(_02996_ ), .B(_03442_ ), .C1(_03445_ ), .C2(_03436_ ), .ZN(_03446_ ) );
NAND3_X1 _11188_ ( .A1(_03425_ ), .A2(_03437_ ), .A3(_03446_ ), .ZN(_03447_ ) );
INV_X1 _11189_ ( .A(\EX_LS_result_reg [24] ), .ZN(_03448_ ) );
OR3_X1 _11190_ ( .A1(_03351_ ), .A2(_03448_ ), .A3(_03352_ ), .ZN(_03449_ ) );
NAND2_X1 _11191_ ( .A1(_03447_ ), .A2(_03449_ ), .ZN(_03450_ ) );
XNOR2_X1 _11192_ ( .A(_03450_ ), .B(_02432_ ), .ZN(_03451_ ) );
OR2_X1 _11193_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03452_ ) );
OAI211_X1 _11194_ ( .A(_03452_ ), .B(_02993_ ), .C1(_03427_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03453_ ) );
OR2_X1 _11195_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03454_ ) );
BUF_X4 _11196_ ( .A(_03295_ ), .Z(_03455_ ) );
OAI211_X1 _11197_ ( .A(_03454_ ), .B(fanout_net_35 ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03456_ ) );
NAND3_X1 _11198_ ( .A1(_03453_ ), .A2(_03456_ ), .A3(_03431_ ), .ZN(_03457_ ) );
MUX2_X1 _11199_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03458_ ) );
MUX2_X1 _11200_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03459_ ) );
BUF_X4 _11201_ ( .A(_02930_ ), .Z(_03460_ ) );
MUX2_X1 _11202_ ( .A(_03458_ ), .B(_03459_ ), .S(_03460_ ), .Z(_03461_ ) );
OAI211_X1 _11203_ ( .A(fanout_net_37 ), .B(_03457_ ), .C1(_03461_ ), .C2(_03436_ ), .ZN(_03462_ ) );
OR2_X1 _11204_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03463_ ) );
OAI211_X1 _11205_ ( .A(_03463_ ), .B(_03460_ ), .C1(_03427_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03464_ ) );
OR2_X1 _11206_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03465_ ) );
OAI211_X1 _11207_ ( .A(_03465_ ), .B(fanout_net_35 ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03466_ ) );
NAND3_X1 _11208_ ( .A1(_03464_ ), .A2(_03466_ ), .A3(_03431_ ), .ZN(_03467_ ) );
MUX2_X1 _11209_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03468_ ) );
MUX2_X1 _11210_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_03469_ ) );
MUX2_X1 _11211_ ( .A(_03468_ ), .B(_03469_ ), .S(_03460_ ), .Z(_03470_ ) );
OAI211_X1 _11212_ ( .A(_02996_ ), .B(_03467_ ), .C1(_03470_ ), .C2(_03436_ ), .ZN(_03471_ ) );
NAND3_X1 _11213_ ( .A1(_03425_ ), .A2(_03462_ ), .A3(_03471_ ), .ZN(_03472_ ) );
INV_X1 _11214_ ( .A(\EX_LS_result_reg [25] ), .ZN(_03473_ ) );
OR3_X1 _11215_ ( .A1(_03351_ ), .A2(_03473_ ), .A3(_03352_ ), .ZN(_03474_ ) );
NAND2_X1 _11216_ ( .A1(_03472_ ), .A2(_03474_ ), .ZN(_03475_ ) );
INV_X1 _11217_ ( .A(_02456_ ), .ZN(_03476_ ) );
NAND2_X1 _11218_ ( .A1(_03475_ ), .A2(_03476_ ), .ZN(_03477_ ) );
NAND3_X1 _11219_ ( .A1(_03472_ ), .A2(_02456_ ), .A3(_03474_ ), .ZN(_03478_ ) );
AND2_X2 _11220_ ( .A1(_03477_ ), .A2(_03478_ ), .ZN(_03479_ ) );
AND2_X1 _11221_ ( .A1(_03451_ ), .A2(_03479_ ), .ZN(_03480_ ) );
OR2_X1 _11222_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03481_ ) );
OAI211_X1 _11223_ ( .A(_03481_ ), .B(_02993_ ), .C1(_03427_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03482_ ) );
OR2_X1 _11224_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03483_ ) );
OAI211_X1 _11225_ ( .A(_03483_ ), .B(fanout_net_35 ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03484_ ) );
NAND3_X1 _11226_ ( .A1(_03482_ ), .A2(_03484_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03485_ ) );
MUX2_X1 _11227_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03486_ ) );
MUX2_X1 _11228_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03487_ ) );
MUX2_X1 _11229_ ( .A(_03486_ ), .B(_03487_ ), .S(_03460_ ), .Z(_03488_ ) );
OAI211_X1 _11230_ ( .A(_02996_ ), .B(_03485_ ), .C1(_03488_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03489_ ) );
NOR2_X1 _11231_ ( .A1(_03455_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03490_ ) );
OAI21_X1 _11232_ ( .A(fanout_net_35 ), .B1(fanout_net_31 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03491_ ) );
MUX2_X1 _11233_ ( .A(_02476_ ), .B(_02477_ ), .S(fanout_net_31 ), .Z(_03492_ ) );
OAI221_X1 _11234_ ( .A(_03431_ ), .B1(_03490_ ), .B2(_03491_ ), .C1(_03492_ ), .C2(fanout_net_35 ), .ZN(_03493_ ) );
MUX2_X1 _11235_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03494_ ) );
MUX2_X1 _11236_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03495_ ) );
MUX2_X1 _11237_ ( .A(_03494_ ), .B(_03495_ ), .S(fanout_net_35 ), .Z(_03496_ ) );
OAI211_X1 _11238_ ( .A(fanout_net_37 ), .B(_03493_ ), .C1(_03496_ ), .C2(_03436_ ), .ZN(_03497_ ) );
NAND3_X1 _11239_ ( .A1(_03425_ ), .A2(_03489_ ), .A3(_03497_ ), .ZN(_03498_ ) );
INV_X1 _11240_ ( .A(\EX_LS_result_reg [27] ), .ZN(_03499_ ) );
OR3_X1 _11241_ ( .A1(_03351_ ), .A2(_03499_ ), .A3(_03352_ ), .ZN(_03500_ ) );
NAND2_X1 _11242_ ( .A1(_03498_ ), .A2(_03500_ ), .ZN(_03501_ ) );
NAND2_X1 _11243_ ( .A1(_02484_ ), .A2(_02486_ ), .ZN(_03502_ ) );
XNOR2_X1 _11244_ ( .A(_03501_ ), .B(_03502_ ), .ZN(_03503_ ) );
OR2_X1 _11245_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03504_ ) );
OAI211_X1 _11246_ ( .A(_03504_ ), .B(_03460_ ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03505_ ) );
OR2_X1 _11247_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03506_ ) );
OAI211_X1 _11248_ ( .A(_03506_ ), .B(fanout_net_35 ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03507_ ) );
NAND3_X1 _11249_ ( .A1(_03505_ ), .A2(_03507_ ), .A3(_03431_ ), .ZN(_03508_ ) );
MUX2_X1 _11250_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03509_ ) );
MUX2_X1 _11251_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03510_ ) );
MUX2_X1 _11252_ ( .A(_03509_ ), .B(_03510_ ), .S(_03460_ ), .Z(_03511_ ) );
OAI211_X1 _11253_ ( .A(fanout_net_37 ), .B(_03508_ ), .C1(_03511_ ), .C2(_03436_ ), .ZN(_03512_ ) );
OAI21_X1 _11254_ ( .A(_02980_ ), .B1(_03295_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03513_ ) );
NOR2_X1 _11255_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03514_ ) );
NOR2_X1 _11256_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03515_ ) );
OAI21_X1 _11257_ ( .A(fanout_net_35 ), .B1(_03295_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03516_ ) );
OAI221_X1 _11258_ ( .A(_03431_ ), .B1(_03513_ ), .B2(_03514_ ), .C1(_03515_ ), .C2(_03516_ ), .ZN(_03517_ ) );
MUX2_X1 _11259_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03518_ ) );
MUX2_X1 _11260_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03519_ ) );
MUX2_X1 _11261_ ( .A(_03518_ ), .B(_03519_ ), .S(_03460_ ), .Z(_03520_ ) );
OAI211_X1 _11262_ ( .A(_02996_ ), .B(_03517_ ), .C1(_03520_ ), .C2(_03436_ ), .ZN(_03521_ ) );
NAND3_X1 _11263_ ( .A1(_03425_ ), .A2(_03512_ ), .A3(_03521_ ), .ZN(_03522_ ) );
INV_X1 _11264_ ( .A(\EX_LS_result_reg [26] ), .ZN(_03523_ ) );
OR3_X1 _11265_ ( .A1(_03351_ ), .A2(_03523_ ), .A3(_03352_ ), .ZN(_03524_ ) );
NAND2_X1 _11266_ ( .A1(_03522_ ), .A2(_03524_ ), .ZN(_03525_ ) );
XNOR2_X1 _11267_ ( .A(_03525_ ), .B(_02510_ ), .ZN(_03526_ ) );
AND3_X1 _11268_ ( .A1(_03480_ ), .A2(_03503_ ), .A3(_03526_ ), .ZN(_03527_ ) );
NAND2_X1 _11269_ ( .A1(_03061_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_03528_ ) );
OR2_X1 _11270_ ( .A1(fanout_net_31 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03529_ ) );
OAI211_X1 _11271_ ( .A(_03529_ ), .B(_02980_ ), .C1(_03295_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03530_ ) );
OR2_X1 _11272_ ( .A1(fanout_net_31 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03531_ ) );
OAI211_X1 _11273_ ( .A(_03531_ ), .B(fanout_net_35 ), .C1(_03295_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03532_ ) );
NAND3_X1 _11274_ ( .A1(_03530_ ), .A2(_03532_ ), .A3(_02938_ ), .ZN(_03533_ ) );
MUX2_X1 _11275_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03534_ ) );
MUX2_X1 _11276_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03535_ ) );
MUX2_X1 _11277_ ( .A(_03534_ ), .B(_03535_ ), .S(_02980_ ), .Z(_03536_ ) );
OAI211_X1 _11278_ ( .A(_02996_ ), .B(_03533_ ), .C1(_03536_ ), .C2(_03431_ ), .ZN(_03537_ ) );
OR2_X1 _11279_ ( .A1(_02875_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03538_ ) );
OAI211_X1 _11280_ ( .A(_03538_ ), .B(fanout_net_35 ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03539_ ) );
OR2_X1 _11281_ ( .A1(fanout_net_31 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03540_ ) );
OAI211_X1 _11282_ ( .A(_03540_ ), .B(_02980_ ), .C1(_03295_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03541_ ) );
NAND3_X1 _11283_ ( .A1(_03539_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03541_ ), .ZN(_03542_ ) );
MUX2_X1 _11284_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03543_ ) );
MUX2_X1 _11285_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03544_ ) );
MUX2_X1 _11286_ ( .A(_03543_ ), .B(_03544_ ), .S(fanout_net_35 ), .Z(_03545_ ) );
OAI211_X1 _11287_ ( .A(fanout_net_37 ), .B(_03542_ ), .C1(_03545_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03546_ ) );
NAND2_X1 _11288_ ( .A1(_03537_ ), .A2(_03546_ ), .ZN(_03547_ ) );
OAI21_X1 _11289_ ( .A(_03547_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_03548_ ) );
AND2_X1 _11290_ ( .A1(_03528_ ), .A2(_03548_ ), .ZN(_03549_ ) );
XOR2_X2 _11291_ ( .A(_01732_ ), .B(_03549_ ), .Z(_03550_ ) );
NAND3_X1 _11292_ ( .A1(_02919_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02037_ ), .ZN(_03551_ ) );
NOR2_X1 _11293_ ( .A1(_03295_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03552_ ) );
OAI21_X1 _11294_ ( .A(fanout_net_35 ), .B1(fanout_net_31 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03553_ ) );
MUX2_X1 _11295_ ( .A(_02551_ ), .B(_02552_ ), .S(fanout_net_31 ), .Z(_03554_ ) );
OAI221_X1 _11296_ ( .A(_02938_ ), .B1(_03552_ ), .B2(_03553_ ), .C1(_03554_ ), .C2(fanout_net_35 ), .ZN(_03555_ ) );
MUX2_X1 _11297_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03556_ ) );
MUX2_X1 _11298_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03557_ ) );
MUX2_X1 _11299_ ( .A(_03556_ ), .B(_03557_ ), .S(fanout_net_35 ), .Z(_03558_ ) );
OAI211_X1 _11300_ ( .A(fanout_net_37 ), .B(_03555_ ), .C1(_03558_ ), .C2(_03431_ ), .ZN(_03559_ ) );
OR2_X1 _11301_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03560_ ) );
OAI211_X1 _11302_ ( .A(_03560_ ), .B(_03460_ ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03561_ ) );
OR2_X1 _11303_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03562_ ) );
OAI211_X1 _11304_ ( .A(_03562_ ), .B(fanout_net_35 ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03563_ ) );
NAND3_X1 _11305_ ( .A1(_03561_ ), .A2(_03563_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03564_ ) );
MUX2_X1 _11306_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_03565_ ) );
MUX2_X1 _11307_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03566_ ) );
MUX2_X1 _11308_ ( .A(_03565_ ), .B(_03566_ ), .S(_02980_ ), .Z(_03567_ ) );
OAI211_X1 _11309_ ( .A(_02996_ ), .B(_03564_ ), .C1(_03567_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03568_ ) );
NAND2_X1 _11310_ ( .A1(_03559_ ), .A2(_03568_ ), .ZN(_03569_ ) );
OAI21_X1 _11311_ ( .A(_03569_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_03570_ ) );
AND2_X1 _11312_ ( .A1(_03551_ ), .A2(_03570_ ), .ZN(_03571_ ) );
XNOR2_X1 _11313_ ( .A(_03571_ ), .B(_02571_ ), .ZN(_03572_ ) );
AND2_X1 _11314_ ( .A1(_03550_ ), .A2(_03572_ ), .ZN(_03573_ ) );
NAND3_X1 _11315_ ( .A1(_02919_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02037_ ), .ZN(_03574_ ) );
NOR2_X1 _11316_ ( .A1(_03455_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03575_ ) );
OAI21_X1 _11317_ ( .A(fanout_net_35 ), .B1(fanout_net_32 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03576_ ) );
MUX2_X1 _11318_ ( .A(_02520_ ), .B(_02521_ ), .S(fanout_net_32 ), .Z(_03577_ ) );
OAI221_X1 _11319_ ( .A(_03431_ ), .B1(_03575_ ), .B2(_03576_ ), .C1(_03577_ ), .C2(fanout_net_35 ), .ZN(_03578_ ) );
MUX2_X1 _11320_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03579_ ) );
MUX2_X1 _11321_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03580_ ) );
MUX2_X1 _11322_ ( .A(_03579_ ), .B(_03580_ ), .S(fanout_net_35 ), .Z(_03581_ ) );
OAI211_X1 _11323_ ( .A(fanout_net_37 ), .B(_03578_ ), .C1(_03581_ ), .C2(_03436_ ), .ZN(_03582_ ) );
OR2_X1 _11324_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03583_ ) );
OAI211_X1 _11325_ ( .A(_03583_ ), .B(_03460_ ), .C1(_03427_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03584_ ) );
OR2_X1 _11326_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03585_ ) );
OAI211_X1 _11327_ ( .A(_03585_ ), .B(fanout_net_35 ), .C1(_03455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03586_ ) );
NAND3_X1 _11328_ ( .A1(_03584_ ), .A2(_03586_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03587_ ) );
MUX2_X1 _11329_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03588_ ) );
MUX2_X1 _11330_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03589_ ) );
MUX2_X1 _11331_ ( .A(_03588_ ), .B(_03589_ ), .S(_03460_ ), .Z(_03590_ ) );
OAI211_X1 _11332_ ( .A(_02996_ ), .B(_03587_ ), .C1(_03590_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03591_ ) );
NAND2_X1 _11333_ ( .A1(_03582_ ), .A2(_03591_ ), .ZN(_03592_ ) );
OAI21_X1 _11334_ ( .A(_03592_ ), .B1(_02899_ ), .B2(_02912_ ), .ZN(_03593_ ) );
AND2_X1 _11335_ ( .A1(_03574_ ), .A2(_03593_ ), .ZN(_03594_ ) );
XNOR2_X1 _11336_ ( .A(_03594_ ), .B(_02539_ ), .ZN(_03595_ ) );
OR2_X1 _11337_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03596_ ) );
OAI211_X1 _11338_ ( .A(_03596_ ), .B(_02993_ ), .C1(_03427_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03597_ ) );
OR2_X1 _11339_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03598_ ) );
OAI211_X1 _11340_ ( .A(_03598_ ), .B(fanout_net_35 ), .C1(_03427_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03599_ ) );
NAND3_X1 _11341_ ( .A1(_03597_ ), .A2(_03599_ ), .A3(_03436_ ), .ZN(_03600_ ) );
MUX2_X1 _11342_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03601_ ) );
MUX2_X1 _11343_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03602_ ) );
MUX2_X1 _11344_ ( .A(_03601_ ), .B(_03602_ ), .S(_02993_ ), .Z(_03603_ ) );
OAI211_X1 _11345_ ( .A(_02996_ ), .B(_03600_ ), .C1(_03603_ ), .C2(_03436_ ), .ZN(_03604_ ) );
OR2_X1 _11346_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03605_ ) );
OAI211_X1 _11347_ ( .A(_03605_ ), .B(fanout_net_35 ), .C1(_03427_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03606_ ) );
OR2_X1 _11348_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03607_ ) );
OAI211_X1 _11349_ ( .A(_03607_ ), .B(_02993_ ), .C1(_03427_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03608_ ) );
NAND3_X1 _11350_ ( .A1(_03606_ ), .A2(_03608_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03609_ ) );
MUX2_X1 _11351_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03610_ ) );
MUX2_X1 _11352_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_03611_ ) );
MUX2_X1 _11353_ ( .A(_03610_ ), .B(_03611_ ), .S(fanout_net_35 ), .Z(_03612_ ) );
OAI211_X1 _11354_ ( .A(fanout_net_37 ), .B(_03609_ ), .C1(_03612_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03613_ ) );
AOI21_X1 _11355_ ( .A(_03061_ ), .B1(_03604_ ), .B2(_03613_ ), .ZN(_03614_ ) );
AND2_X1 _11356_ ( .A1(_03061_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_03615_ ) );
NOR2_X1 _11357_ ( .A1(_03614_ ), .A2(_03615_ ), .ZN(_03616_ ) );
XNOR2_X1 _11358_ ( .A(_03616_ ), .B(_01765_ ), .ZN(_03617_ ) );
AND2_X1 _11359_ ( .A1(_03595_ ), .A2(_03617_ ), .ZN(_03618_ ) );
AND3_X4 _11360_ ( .A1(_03527_ ), .A2(_03573_ ), .A3(_03618_ ), .ZN(_03619_ ) );
AND3_X1 _11361_ ( .A1(_03111_ ), .A2(_03424_ ), .A3(_03619_ ), .ZN(_03620_ ) );
INV_X1 _11362_ ( .A(\EX_LS_result_reg [1] ), .ZN(_03621_ ) );
OR3_X4 _11363_ ( .A1(_02910_ ), .A2(_03621_ ), .A3(_02897_ ), .ZN(_03622_ ) );
NOR2_X1 _11364_ ( .A1(_02982_ ), .A2(\myreg.Reg[11][1] ), .ZN(_03623_ ) );
OAI21_X1 _11365_ ( .A(fanout_net_35 ), .B1(fanout_net_32 ), .B2(\myreg.Reg[10][1] ), .ZN(_03624_ ) );
NOR2_X1 _11366_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][1] ), .ZN(_03625_ ) );
OAI21_X1 _11367_ ( .A(_02880_ ), .B1(_02982_ ), .B2(\myreg.Reg[9][1] ), .ZN(_03626_ ) );
OAI221_X1 _11368_ ( .A(_02867_ ), .B1(_03623_ ), .B2(_03624_ ), .C1(_03625_ ), .C2(_03626_ ), .ZN(_03627_ ) );
MUX2_X1 _11369_ ( .A(\myreg.Reg[12][1] ), .B(\myreg.Reg[13][1] ), .S(fanout_net_32 ), .Z(_03628_ ) );
MUX2_X1 _11370_ ( .A(\myreg.Reg[14][1] ), .B(\myreg.Reg[15][1] ), .S(fanout_net_32 ), .Z(_03629_ ) );
MUX2_X1 _11371_ ( .A(_03628_ ), .B(_03629_ ), .S(fanout_net_35 ), .Z(_03630_ ) );
OAI211_X1 _11372_ ( .A(fanout_net_37 ), .B(_03627_ ), .C1(_03630_ ), .C2(_02868_ ), .ZN(_03631_ ) );
OR2_X1 _11373_ ( .A1(_02862_ ), .A2(\myreg.Reg[5][1] ), .ZN(_03632_ ) );
OAI211_X1 _11374_ ( .A(_03632_ ), .B(_02880_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[4][1] ), .ZN(_03633_ ) );
OR2_X1 _11375_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[6][1] ), .ZN(_03634_ ) );
OAI211_X1 _11376_ ( .A(_03634_ ), .B(fanout_net_35 ), .C1(_02982_ ), .C2(\myreg.Reg[7][1] ), .ZN(_03635_ ) );
NAND3_X1 _11377_ ( .A1(_03633_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03635_ ), .ZN(_03636_ ) );
MUX2_X1 _11378_ ( .A(\myreg.Reg[2][1] ), .B(\myreg.Reg[3][1] ), .S(fanout_net_32 ), .Z(_03637_ ) );
MUX2_X1 _11379_ ( .A(\myreg.Reg[0][1] ), .B(\myreg.Reg[1][1] ), .S(fanout_net_32 ), .Z(_03638_ ) );
MUX2_X1 _11380_ ( .A(_03637_ ), .B(_03638_ ), .S(_02880_ ), .Z(_03639_ ) );
OAI211_X1 _11381_ ( .A(_02889_ ), .B(_03636_ ), .C1(_03639_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03640_ ) );
NAND2_X1 _11382_ ( .A1(_03631_ ), .A2(_03640_ ), .ZN(_03641_ ) );
OAI21_X1 _11383_ ( .A(_03641_ ), .B1(_02898_ ), .B2(_02910_ ), .ZN(_03642_ ) );
AND2_X1 _11384_ ( .A1(_03622_ ), .A2(_03642_ ), .ZN(_03643_ ) );
XNOR2_X2 _11385_ ( .A(_02041_ ), .B(_03643_ ), .ZN(_03644_ ) );
AND2_X2 _11386_ ( .A1(_02036_ ), .A2(_02038_ ), .ZN(_03645_ ) );
INV_X1 _11387_ ( .A(_03645_ ), .ZN(_03646_ ) );
INV_X1 _11388_ ( .A(\EX_LS_result_reg [0] ), .ZN(_03647_ ) );
OR3_X1 _11389_ ( .A1(_02910_ ), .A2(_03647_ ), .A3(_02897_ ), .ZN(_03648_ ) );
OR2_X1 _11390_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][0] ), .ZN(_03649_ ) );
OAI211_X1 _11391_ ( .A(_03649_ ), .B(_02872_ ), .C1(_03141_ ), .C2(\myreg.Reg[1][0] ), .ZN(_03650_ ) );
OR2_X1 _11392_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][0] ), .ZN(_03651_ ) );
OAI211_X1 _11393_ ( .A(_03651_ ), .B(fanout_net_35 ), .C1(_02874_ ), .C2(\myreg.Reg[3][0] ), .ZN(_03652_ ) );
NAND3_X1 _11394_ ( .A1(_03650_ ), .A2(_03652_ ), .A3(_02868_ ), .ZN(_03653_ ) );
MUX2_X1 _11395_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_32 ), .Z(_03654_ ) );
MUX2_X1 _11396_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_32 ), .Z(_03655_ ) );
MUX2_X1 _11397_ ( .A(_03654_ ), .B(_03655_ ), .S(_02880_ ), .Z(_03656_ ) );
OAI211_X1 _11398_ ( .A(_03019_ ), .B(_03653_ ), .C1(_03656_ ), .C2(_02868_ ), .ZN(_03657_ ) );
OR2_X1 _11399_ ( .A1(_02862_ ), .A2(\myreg.Reg[13][0] ), .ZN(_03658_ ) );
OAI211_X1 _11400_ ( .A(_03658_ ), .B(_03153_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[12][0] ), .ZN(_03659_ ) );
OR2_X1 _11401_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[14][0] ), .ZN(_03660_ ) );
OAI211_X1 _11402_ ( .A(_03660_ ), .B(fanout_net_35 ), .C1(_02874_ ), .C2(\myreg.Reg[15][0] ), .ZN(_03661_ ) );
NAND3_X1 _11403_ ( .A1(_03659_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03661_ ), .ZN(_03662_ ) );
MUX2_X1 _11404_ ( .A(\myreg.Reg[8][0] ), .B(\myreg.Reg[9][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03663_ ) );
MUX2_X1 _11405_ ( .A(\myreg.Reg[10][0] ), .B(\myreg.Reg[11][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03664_ ) );
MUX2_X1 _11406_ ( .A(_03663_ ), .B(_03664_ ), .S(fanout_net_35 ), .Z(_03665_ ) );
OAI211_X1 _11407_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03662_ ), .C1(_03665_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03666_ ) );
NAND2_X1 _11408_ ( .A1(_03657_ ), .A2(_03666_ ), .ZN(_03667_ ) );
OAI21_X4 _11409_ ( .A(_03667_ ), .B1(_02898_ ), .B2(_02911_ ), .ZN(_03668_ ) );
AND2_X1 _11410_ ( .A1(_03648_ ), .A2(_03668_ ), .ZN(_03669_ ) );
XNOR2_X1 _11411_ ( .A(_03646_ ), .B(_03669_ ), .ZN(_03670_ ) );
NAND2_X1 _11412_ ( .A1(_03644_ ), .A2(_03670_ ), .ZN(_03671_ ) );
OR3_X1 _11413_ ( .A1(_03351_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03352_ ), .ZN(_03672_ ) );
OR2_X1 _11414_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03673_ ) );
OAI211_X1 _11415_ ( .A(_03673_ ), .B(_02872_ ), .C1(_02864_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03674_ ) );
OR2_X1 _11416_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03675_ ) );
OAI211_X1 _11417_ ( .A(_03675_ ), .B(fanout_net_35 ), .C1(_03141_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03676_ ) );
NAND3_X1 _11418_ ( .A1(_03674_ ), .A2(_03676_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03677_ ) );
MUX2_X1 _11419_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03678_ ) );
MUX2_X1 _11420_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03679_ ) );
MUX2_X1 _11421_ ( .A(_03678_ ), .B(_03679_ ), .S(_03153_ ), .Z(_03680_ ) );
OAI211_X1 _11422_ ( .A(_03019_ ), .B(_03677_ ), .C1(_03680_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03681_ ) );
NOR2_X1 _11423_ ( .A1(_02982_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03682_ ) );
OAI21_X1 _11424_ ( .A(fanout_net_35 ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03683_ ) );
MUX2_X1 _11425_ ( .A(_02050_ ), .B(_02051_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03684_ ) );
OAI221_X1 _11426_ ( .A(_02867_ ), .B1(_03682_ ), .B2(_03683_ ), .C1(_03684_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_03685_ ) );
MUX2_X1 _11427_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03686_ ) );
MUX2_X1 _11428_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03687_ ) );
MUX2_X1 _11429_ ( .A(_03686_ ), .B(_03687_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03688_ ) );
OAI211_X1 _11430_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03685_ ), .C1(_03688_ ), .C2(_03113_ ), .ZN(_03689_ ) );
OAI211_X1 _11431_ ( .A(_03681_ ), .B(_03689_ ), .C1(_03351_ ), .C2(_03352_ ), .ZN(_03690_ ) );
NAND2_X1 _11432_ ( .A1(_03672_ ), .A2(_03690_ ), .ZN(_03691_ ) );
XNOR2_X1 _11433_ ( .A(_03691_ ), .B(_02069_ ), .ZN(_03692_ ) );
INV_X1 _11434_ ( .A(_03692_ ), .ZN(_03693_ ) );
INV_X1 _11435_ ( .A(\EX_LS_result_reg [2] ), .ZN(_03694_ ) );
OR3_X1 _11436_ ( .A1(_02910_ ), .A2(_03694_ ), .A3(_02897_ ), .ZN(_03695_ ) );
OR2_X1 _11437_ ( .A1(_02863_ ), .A2(\myreg.Reg[1][2] ), .ZN(_03696_ ) );
OAI211_X1 _11438_ ( .A(_03696_ ), .B(_02872_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[0][2] ), .ZN(_03697_ ) );
OR2_X1 _11439_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[2][2] ), .ZN(_03698_ ) );
OAI211_X1 _11440_ ( .A(_03698_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03141_ ), .C2(\myreg.Reg[3][2] ), .ZN(_03699_ ) );
NAND3_X1 _11441_ ( .A1(_03697_ ), .A2(_02868_ ), .A3(_03699_ ), .ZN(_03700_ ) );
MUX2_X1 _11442_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03701_ ) );
MUX2_X1 _11443_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03702_ ) );
MUX2_X1 _11444_ ( .A(_03701_ ), .B(_03702_ ), .S(_03153_ ), .Z(_03703_ ) );
OAI211_X1 _11445_ ( .A(_03019_ ), .B(_03700_ ), .C1(_03703_ ), .C2(_03113_ ), .ZN(_03704_ ) );
OR2_X1 _11446_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[14][2] ), .ZN(_03705_ ) );
OAI211_X1 _11447_ ( .A(_03705_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03141_ ), .C2(\myreg.Reg[15][2] ), .ZN(_03706_ ) );
OR2_X1 _11448_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[12][2] ), .ZN(_03707_ ) );
OAI211_X1 _11449_ ( .A(_03707_ ), .B(_03153_ ), .C1(_03141_ ), .C2(\myreg.Reg[13][2] ), .ZN(_03708_ ) );
NAND3_X1 _11450_ ( .A1(_03706_ ), .A2(_03708_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03709_ ) );
MUX2_X1 _11451_ ( .A(\myreg.Reg[8][2] ), .B(\myreg.Reg[9][2] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03710_ ) );
MUX2_X1 _11452_ ( .A(\myreg.Reg[10][2] ), .B(\myreg.Reg[11][2] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03711_ ) );
MUX2_X1 _11453_ ( .A(_03710_ ), .B(_03711_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03712_ ) );
OAI211_X1 _11454_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03709_ ), .C1(_03712_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03713_ ) );
NAND2_X1 _11455_ ( .A1(_03704_ ), .A2(_03713_ ), .ZN(_03714_ ) );
OAI21_X2 _11456_ ( .A(_03714_ ), .B1(_02898_ ), .B2(_02911_ ), .ZN(_03715_ ) );
AND2_X1 _11457_ ( .A1(_03695_ ), .A2(_03715_ ), .ZN(_03716_ ) );
INV_X1 _11458_ ( .A(_02045_ ), .ZN(_03717_ ) );
XNOR2_X1 _11459_ ( .A(_03716_ ), .B(_03717_ ), .ZN(_03718_ ) );
INV_X1 _11460_ ( .A(_03718_ ), .ZN(_03719_ ) );
NOR3_X1 _11461_ ( .A1(_03671_ ), .A2(_03693_ ), .A3(_03719_ ), .ZN(_03720_ ) );
AND2_X1 _11462_ ( .A1(_03620_ ), .A2(_03720_ ), .ZN(_03721_ ) );
NOR2_X1 _11463_ ( .A1(_02832_ ), .A2(\ID_EX_typ [1] ), .ZN(_03722_ ) );
AND2_X2 _11464_ ( .A1(_03722_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_03723_ ) );
INV_X1 _11465_ ( .A(_03723_ ), .ZN(_03724_ ) );
INV_X1 _11466_ ( .A(fanout_net_11 ), .ZN(_03725_ ) );
BUF_X4 _11467_ ( .A(_03725_ ), .Z(_03726_ ) );
BUF_X4 _11468_ ( .A(_03726_ ), .Z(_03727_ ) );
BUF_X2 _11469_ ( .A(_03727_ ), .Z(_03728_ ) );
OAI21_X1 _11470_ ( .A(_03728_ ), .B1(_03614_ ), .B2(_03615_ ), .ZN(_03729_ ) );
NAND2_X1 _11471_ ( .A1(fanout_net_11 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03730_ ) );
AND2_X2 _11472_ ( .A1(_03729_ ), .A2(_03730_ ), .ZN(_03731_ ) );
INV_X1 _11473_ ( .A(_01765_ ), .ZN(_03732_ ) );
XNOR2_X1 _11474_ ( .A(_03731_ ), .B(_03732_ ), .ZN(_03733_ ) );
INV_X1 _11475_ ( .A(_03733_ ), .ZN(_03734_ ) );
NAND3_X1 _11476_ ( .A1(_03574_ ), .A2(_03728_ ), .A3(_03593_ ), .ZN(_03735_ ) );
NAND2_X1 _11477_ ( .A1(_02544_ ), .A2(fanout_net_11 ), .ZN(_03736_ ) );
NAND2_X1 _11478_ ( .A1(_03735_ ), .A2(_03736_ ), .ZN(_03737_ ) );
INV_X1 _11479_ ( .A(_02539_ ), .ZN(_03738_ ) );
XNOR2_X1 _11480_ ( .A(_03737_ ), .B(_03738_ ), .ZN(_03739_ ) );
INV_X1 _11481_ ( .A(_03739_ ), .ZN(_03740_ ) );
NAND3_X1 _11482_ ( .A1(_03528_ ), .A2(_03548_ ), .A3(_03728_ ), .ZN(_03741_ ) );
OR2_X1 _11483_ ( .A1(_03728_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03742_ ) );
AND3_X1 _11484_ ( .A1(_01732_ ), .A2(_03741_ ), .A3(_03742_ ), .ZN(_03743_ ) );
AOI21_X1 _11485_ ( .A(_01732_ ), .B1(_03741_ ), .B2(_03742_ ), .ZN(_03744_ ) );
NOR2_X1 _11486_ ( .A1(_03743_ ), .A2(_03744_ ), .ZN(_03745_ ) );
NAND3_X1 _11487_ ( .A1(_03551_ ), .A2(_03728_ ), .A3(_03570_ ), .ZN(_03746_ ) );
INV_X1 _11488_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_03747_ ) );
NAND2_X1 _11489_ ( .A1(_03747_ ), .A2(fanout_net_11 ), .ZN(_03748_ ) );
AOI21_X1 _11490_ ( .A(_02571_ ), .B1(_03746_ ), .B2(_03748_ ), .ZN(_03749_ ) );
AND3_X1 _11491_ ( .A1(_03746_ ), .A2(_02571_ ), .A3(_03748_ ), .ZN(_03750_ ) );
NOR3_X1 _11492_ ( .A1(_03745_ ), .A2(_03749_ ), .A3(_03750_ ), .ZN(_03751_ ) );
NAND3_X1 _11493_ ( .A1(_03734_ ), .A2(_03740_ ), .A3(_03751_ ), .ZN(_03752_ ) );
NAND3_X1 _11494_ ( .A1(_03522_ ), .A2(_03727_ ), .A3(_03524_ ), .ZN(_03753_ ) );
NAND2_X1 _11495_ ( .A1(_02511_ ), .A2(fanout_net_11 ), .ZN(_03754_ ) );
NAND2_X1 _11496_ ( .A1(_03753_ ), .A2(_03754_ ), .ZN(_03755_ ) );
NOR2_X4 _11497_ ( .A1(_03755_ ), .A2(_02514_ ), .ZN(_03756_ ) );
AOI21_X1 _11498_ ( .A(_02510_ ), .B1(_03753_ ), .B2(_03754_ ), .ZN(_03757_ ) );
NOR2_X1 _11499_ ( .A1(_03756_ ), .A2(_03757_ ), .ZN(_03758_ ) );
INV_X2 _11500_ ( .A(_03758_ ), .ZN(_03759_ ) );
NAND3_X1 _11501_ ( .A1(_03498_ ), .A2(_03727_ ), .A3(_03500_ ), .ZN(_03760_ ) );
NAND2_X1 _11502_ ( .A1(_02485_ ), .A2(fanout_net_11 ), .ZN(_03761_ ) );
NAND2_X1 _11503_ ( .A1(_03760_ ), .A2(_03761_ ), .ZN(_03762_ ) );
INV_X1 _11504_ ( .A(_03502_ ), .ZN(_03763_ ) );
NOR2_X1 _11505_ ( .A1(_03762_ ), .A2(_03763_ ), .ZN(_03764_ ) );
AOI21_X1 _11506_ ( .A(_03502_ ), .B1(_03760_ ), .B2(_03761_ ), .ZN(_03765_ ) );
NOR2_X1 _11507_ ( .A1(_03764_ ), .A2(_03765_ ), .ZN(_03766_ ) );
INV_X1 _11508_ ( .A(_03766_ ), .ZN(_03767_ ) );
NAND2_X1 _11509_ ( .A1(_03759_ ), .A2(_03767_ ), .ZN(_03768_ ) );
NAND3_X1 _11510_ ( .A1(_03447_ ), .A2(_03728_ ), .A3(_03449_ ), .ZN(_03769_ ) );
NAND2_X1 _11511_ ( .A1(_02433_ ), .A2(fanout_net_11 ), .ZN(_03770_ ) );
NAND2_X1 _11512_ ( .A1(_03769_ ), .A2(_03770_ ), .ZN(_03771_ ) );
XNOR2_X1 _11513_ ( .A(_03771_ ), .B(_02432_ ), .ZN(_03772_ ) );
NAND3_X1 _11514_ ( .A1(_03472_ ), .A2(_03727_ ), .A3(_03474_ ), .ZN(_03773_ ) );
NAND2_X1 _11515_ ( .A1(_02457_ ), .A2(fanout_net_11 ), .ZN(_03774_ ) );
NAND2_X1 _11516_ ( .A1(_03773_ ), .A2(_03774_ ), .ZN(_03775_ ) );
NOR2_X1 _11517_ ( .A1(_03775_ ), .A2(_03476_ ), .ZN(_03776_ ) );
AOI21_X1 _11518_ ( .A(_02456_ ), .B1(_03773_ ), .B2(_03774_ ), .ZN(_03777_ ) );
NOR2_X1 _11519_ ( .A1(_03776_ ), .A2(_03777_ ), .ZN(_03778_ ) );
NOR3_X1 _11520_ ( .A1(_03768_ ), .A2(_03772_ ), .A3(_03778_ ), .ZN(_03779_ ) );
NAND3_X1 _11521_ ( .A1(_03009_ ), .A2(_03726_ ), .A3(_03031_ ), .ZN(_03780_ ) );
NAND2_X1 _11522_ ( .A1(_01794_ ), .A2(fanout_net_11 ), .ZN(_03781_ ) );
NAND2_X2 _11523_ ( .A1(_03780_ ), .A2(_03781_ ), .ZN(_03782_ ) );
XNOR2_X2 _11524_ ( .A(_03782_ ), .B(_01793_ ), .ZN(_03783_ ) );
INV_X2 _11525_ ( .A(_03783_ ), .ZN(_03784_ ) );
OR2_X4 _11526_ ( .A1(_03057_ ), .A2(fanout_net_11 ), .ZN(_03785_ ) );
NAND2_X1 _11527_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [23] ), .ZN(_03786_ ) );
AND2_X4 _11528_ ( .A1(_03785_ ), .A2(_03786_ ), .ZN(_03787_ ) );
NOR2_X4 _11529_ ( .A1(_03787_ ), .A2(_03058_ ), .ZN(_03788_ ) );
AND3_X4 _11530_ ( .A1(_03785_ ), .A2(_03058_ ), .A3(_03786_ ), .ZN(_03789_ ) );
OAI21_X4 _11531_ ( .A(_03784_ ), .B1(_03788_ ), .B2(_03789_ ), .ZN(_03790_ ) );
OAI21_X1 _11532_ ( .A(_03727_ ), .B1(_03080_ ), .B2(_03082_ ), .ZN(_03791_ ) );
NAND2_X1 _11533_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [20] ), .ZN(_03792_ ) );
AND2_X2 _11534_ ( .A1(_03791_ ), .A2(_03792_ ), .ZN(_03793_ ) );
XNOR2_X2 _11535_ ( .A(_03793_ ), .B(_01869_ ), .ZN(_03794_ ) );
NAND3_X1 _11536_ ( .A1(_03087_ ), .A2(_03107_ ), .A3(_03726_ ), .ZN(_03795_ ) );
NAND2_X1 _11537_ ( .A1(_01844_ ), .A2(fanout_net_11 ), .ZN(_03796_ ) );
NAND2_X2 _11538_ ( .A1(_03795_ ), .A2(_03796_ ), .ZN(_03797_ ) );
XNOR2_X2 _11539_ ( .A(_03797_ ), .B(_01843_ ), .ZN(_03798_ ) );
NOR3_X1 _11540_ ( .A1(_03790_ ), .A2(_03794_ ), .A3(_03798_ ), .ZN(_03799_ ) );
NAND3_X1 _11541_ ( .A1(_02974_ ), .A2(_03727_ ), .A3(_02975_ ), .ZN(_03800_ ) );
NAND2_X1 _11542_ ( .A1(_01919_ ), .A2(fanout_net_11 ), .ZN(_03801_ ) );
NAND2_X1 _11543_ ( .A1(_03800_ ), .A2(_03801_ ), .ZN(_03802_ ) );
NAND2_X1 _11544_ ( .A1(_03802_ ), .A2(_01918_ ), .ZN(_03803_ ) );
AOI21_X1 _11545_ ( .A(fanout_net_11 ), .B1(_02913_ ), .B2(_02920_ ), .ZN(_03804_ ) );
AND2_X1 _11546_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [17] ), .ZN(_03805_ ) );
NOR2_X2 _11547_ ( .A1(_03804_ ), .A2(_03805_ ), .ZN(_03806_ ) );
XNOR2_X1 _11548_ ( .A(_03806_ ), .B(_01942_ ), .ZN(_03807_ ) );
NAND3_X2 _11549_ ( .A1(_02927_ ), .A2(_02951_ ), .A3(_03727_ ), .ZN(_03808_ ) );
NAND2_X1 _11550_ ( .A1(_01966_ ), .A2(fanout_net_11 ), .ZN(_03809_ ) );
NAND2_X2 _11551_ ( .A1(_03808_ ), .A2(_03809_ ), .ZN(_03810_ ) );
INV_X1 _11552_ ( .A(_03810_ ), .ZN(_03811_ ) );
NOR3_X1 _11553_ ( .A1(_03807_ ), .A2(_02953_ ), .A3(_03811_ ), .ZN(_03812_ ) );
AOI21_X1 _11554_ ( .A(_03812_ ), .B1(_01942_ ), .B2(_03806_ ), .ZN(_03813_ ) );
XNOR2_X1 _11555_ ( .A(_03802_ ), .B(_01918_ ), .ZN(_03814_ ) );
INV_X1 _11556_ ( .A(_03814_ ), .ZN(_03815_ ) );
NAND3_X1 _11557_ ( .A1(_03002_ ), .A2(_03727_ ), .A3(_03003_ ), .ZN(_03816_ ) );
NAND2_X1 _11558_ ( .A1(_01896_ ), .A2(fanout_net_11 ), .ZN(_03817_ ) );
NAND2_X1 _11559_ ( .A1(_03816_ ), .A2(_03817_ ), .ZN(_03818_ ) );
XNOR2_X1 _11560_ ( .A(_03818_ ), .B(_01895_ ), .ZN(_03819_ ) );
INV_X1 _11561_ ( .A(_03819_ ), .ZN(_03820_ ) );
NAND2_X1 _11562_ ( .A1(_03815_ ), .A2(_03820_ ), .ZN(_03821_ ) );
OAI21_X1 _11563_ ( .A(_03803_ ), .B1(_03813_ ), .B2(_03821_ ), .ZN(_03822_ ) );
AND3_X1 _11564_ ( .A1(_03815_ ), .A2(_01895_ ), .A3(_03818_ ), .ZN(_03823_ ) );
OAI21_X1 _11565_ ( .A(_03799_ ), .B1(_03822_ ), .B2(_03823_ ), .ZN(_03824_ ) );
NAND2_X1 _11566_ ( .A1(_03797_ ), .A2(_01843_ ), .ZN(_03825_ ) );
AND2_X1 _11567_ ( .A1(_03797_ ), .A2(_02403_ ), .ZN(_03826_ ) );
NOR2_X1 _11568_ ( .A1(_03797_ ), .A2(_02403_ ), .ZN(_03827_ ) );
OAI211_X1 _11569_ ( .A(_01869_ ), .B(_03793_ ), .C1(_03826_ ), .C2(_03827_ ), .ZN(_03828_ ) );
AOI21_X1 _11570_ ( .A(_03790_ ), .B1(_03825_ ), .B2(_03828_ ), .ZN(_03829_ ) );
AOI21_X1 _11571_ ( .A(_03829_ ), .B1(_01816_ ), .B2(_03787_ ), .ZN(_03830_ ) );
AOI21_X1 _11572_ ( .A(fanout_net_11 ), .B1(_03139_ ), .B2(_03161_ ), .ZN(_03831_ ) );
AND2_X1 _11573_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [15] ), .ZN(_03832_ ) );
NOR2_X2 _11574_ ( .A1(_03831_ ), .A2(_03832_ ), .ZN(_03833_ ) );
XNOR2_X2 _11575_ ( .A(_03833_ ), .B(_02309_ ), .ZN(_03834_ ) );
INV_X1 _11576_ ( .A(_03834_ ), .ZN(_03835_ ) );
NAND3_X1 _11577_ ( .A1(_03112_ ), .A2(_03726_ ), .A3(_03133_ ), .ZN(_03836_ ) );
NAND2_X1 _11578_ ( .A1(_02333_ ), .A2(fanout_net_11 ), .ZN(_03837_ ) );
NAND2_X1 _11579_ ( .A1(_03836_ ), .A2(_03837_ ), .ZN(_03838_ ) );
XNOR2_X2 _11580_ ( .A(_03838_ ), .B(_02332_ ), .ZN(_03839_ ) );
INV_X1 _11581_ ( .A(_03839_ ), .ZN(_03840_ ) );
NAND3_X1 _11582_ ( .A1(_03166_ ), .A2(_03186_ ), .A3(_03726_ ), .ZN(_03841_ ) );
NAND2_X1 _11583_ ( .A1(_02381_ ), .A2(fanout_net_11 ), .ZN(_03842_ ) );
NAND2_X2 _11584_ ( .A1(_03841_ ), .A2(_03842_ ), .ZN(_03843_ ) );
XNOR2_X2 _11585_ ( .A(_03843_ ), .B(_02380_ ), .ZN(_03844_ ) );
INV_X2 _11586_ ( .A(_03844_ ), .ZN(_03845_ ) );
NAND3_X2 _11587_ ( .A1(_03835_ ), .A2(_03840_ ), .A3(_03845_ ), .ZN(_03846_ ) );
NAND3_X1 _11588_ ( .A1(_03191_ ), .A2(_03211_ ), .A3(_03727_ ), .ZN(_03847_ ) );
NAND2_X1 _11589_ ( .A1(_02355_ ), .A2(fanout_net_11 ), .ZN(_03848_ ) );
NAND2_X2 _11590_ ( .A1(_03847_ ), .A2(_03848_ ), .ZN(_03849_ ) );
XNOR2_X1 _11591_ ( .A(_03849_ ), .B(_03213_ ), .ZN(_03850_ ) );
NOR2_X2 _11592_ ( .A1(_03846_ ), .A2(_03850_ ), .ZN(_03851_ ) );
NAND3_X1 _11593_ ( .A1(_03244_ ), .A2(_03264_ ), .A3(_03726_ ), .ZN(_03852_ ) );
NAND2_X1 _11594_ ( .A1(_02250_ ), .A2(fanout_net_11 ), .ZN(_03853_ ) );
NAND2_X1 _11595_ ( .A1(_03852_ ), .A2(_03853_ ), .ZN(_03854_ ) );
XNOR2_X1 _11596_ ( .A(_03854_ ), .B(_02249_ ), .ZN(_03855_ ) );
NAND3_X1 _11597_ ( .A1(_03219_ ), .A2(_03239_ ), .A3(_03726_ ), .ZN(_03856_ ) );
NAND2_X1 _11598_ ( .A1(_02273_ ), .A2(fanout_net_11 ), .ZN(_03857_ ) );
NAND2_X1 _11599_ ( .A1(_03856_ ), .A2(_03857_ ), .ZN(_03858_ ) );
XNOR2_X1 _11600_ ( .A(_03858_ ), .B(_02272_ ), .ZN(_03859_ ) );
NOR2_X1 _11601_ ( .A1(_03855_ ), .A2(_03859_ ), .ZN(_03860_ ) );
NAND3_X1 _11602_ ( .A1(_03270_ ), .A2(_03290_ ), .A3(_03726_ ), .ZN(_03861_ ) );
NAND2_X1 _11603_ ( .A1(_02226_ ), .A2(fanout_net_11 ), .ZN(_03862_ ) );
NAND2_X1 _11604_ ( .A1(_03861_ ), .A2(_03862_ ), .ZN(_03863_ ) );
XNOR2_X1 _11605_ ( .A(_03863_ ), .B(_02225_ ), .ZN(_03864_ ) );
INV_X1 _11606_ ( .A(_03864_ ), .ZN(_03865_ ) );
OAI21_X1 _11607_ ( .A(_03727_ ), .B1(_03313_ ), .B2(_03315_ ), .ZN(_03866_ ) );
NAND2_X1 _11608_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [8] ), .ZN(_03867_ ) );
AND2_X1 _11609_ ( .A1(_03866_ ), .A2(_03867_ ), .ZN(_03868_ ) );
XNOR2_X1 _11610_ ( .A(_03868_ ), .B(_02202_ ), .ZN(_03869_ ) );
INV_X1 _11611_ ( .A(_03869_ ), .ZN(_03870_ ) );
NAND4_X1 _11612_ ( .A1(_03851_ ), .A2(_03860_ ), .A3(_03865_ ), .A4(_03870_ ), .ZN(_03871_ ) );
OR2_X4 _11613_ ( .A1(_03341_ ), .A2(fanout_net_11 ), .ZN(_03872_ ) );
NAND2_X1 _11614_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [7] ), .ZN(_03873_ ) );
AND2_X2 _11615_ ( .A1(_03872_ ), .A2(_03873_ ), .ZN(_03874_ ) );
NOR2_X2 _11616_ ( .A1(_03874_ ), .A2(_03342_ ), .ZN(_03875_ ) );
AND3_X1 _11617_ ( .A1(_03872_ ), .A2(_03342_ ), .A3(_03873_ ), .ZN(_03876_ ) );
NOR2_X4 _11618_ ( .A1(_03875_ ), .A2(_03876_ ), .ZN(_03877_ ) );
INV_X4 _11619_ ( .A(_03877_ ), .ZN(_03878_ ) );
NAND3_X1 _11620_ ( .A1(_03353_ ), .A2(_03725_ ), .A3(_03372_ ), .ZN(_03879_ ) );
NAND2_X1 _11621_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [6] ), .ZN(_03880_ ) );
AND2_X4 _11622_ ( .A1(_03879_ ), .A2(_03880_ ), .ZN(_03881_ ) );
XNOR2_X1 _11623_ ( .A(_03881_ ), .B(_02171_ ), .ZN(_03882_ ) );
INV_X1 _11624_ ( .A(_03882_ ), .ZN(_03883_ ) );
NAND3_X1 _11625_ ( .A1(_03399_ ), .A2(_03419_ ), .A3(_03725_ ), .ZN(_03884_ ) );
NAND2_X1 _11626_ ( .A1(_02119_ ), .A2(\ID_EX_typ [4] ), .ZN(_03885_ ) );
NAND2_X2 _11627_ ( .A1(_03884_ ), .A2(_03885_ ), .ZN(_03886_ ) );
NAND3_X1 _11628_ ( .A1(_03376_ ), .A2(_03725_ ), .A3(_03396_ ), .ZN(_03887_ ) );
NAND2_X1 _11629_ ( .A1(_02125_ ), .A2(\ID_EX_typ [4] ), .ZN(_03888_ ) );
NAND2_X4 _11630_ ( .A1(_03887_ ), .A2(_03888_ ), .ZN(_03889_ ) );
AND2_X1 _11631_ ( .A1(_03889_ ), .A2(_02096_ ), .ZN(_03890_ ) );
INV_X1 _11632_ ( .A(_02096_ ), .ZN(_03891_ ) );
AND3_X1 _11633_ ( .A1(_03891_ ), .A2(_03887_ ), .A3(_03888_ ), .ZN(_03892_ ) );
OAI211_X1 _11634_ ( .A(_02118_ ), .B(_03886_ ), .C1(_03890_ ), .C2(_03892_ ), .ZN(_03893_ ) );
OAI21_X1 _11635_ ( .A(_03893_ ), .B1(_03891_ ), .B2(_03889_ ), .ZN(_03894_ ) );
AND3_X1 _11636_ ( .A1(_03878_ ), .A2(_03883_ ), .A3(_03894_ ), .ZN(_03895_ ) );
XNOR2_X1 _11637_ ( .A(_03889_ ), .B(_03891_ ), .ZN(_03896_ ) );
INV_X1 _11638_ ( .A(_03896_ ), .ZN(_03897_ ) );
XNOR2_X1 _11639_ ( .A(_03886_ ), .B(_02118_ ), .ZN(_03898_ ) );
INV_X1 _11640_ ( .A(_03898_ ), .ZN(_03899_ ) );
NAND4_X1 _11641_ ( .A1(_03878_ ), .A2(_03883_ ), .A3(_03897_ ), .A4(_03899_ ), .ZN(_03900_ ) );
NAND3_X1 _11642_ ( .A1(_03672_ ), .A2(_03725_ ), .A3(_03690_ ), .ZN(_03901_ ) );
NAND2_X1 _11643_ ( .A1(\ID_EX_typ [4] ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_03902_ ) );
AND2_X1 _11644_ ( .A1(_03901_ ), .A2(_03902_ ), .ZN(_03903_ ) );
INV_X1 _11645_ ( .A(_02069_ ), .ZN(_03904_ ) );
XNOR2_X2 _11646_ ( .A(_03903_ ), .B(_03904_ ), .ZN(_03905_ ) );
NAND3_X2 _11647_ ( .A1(_03695_ ), .A2(_03715_ ), .A3(_03726_ ), .ZN(_03906_ ) );
NAND2_X1 _11648_ ( .A1(_01969_ ), .A2(\ID_EX_typ [4] ), .ZN(_03907_ ) );
NAND2_X4 _11649_ ( .A1(_03906_ ), .A2(_03907_ ), .ZN(_03908_ ) );
INV_X1 _11650_ ( .A(_03908_ ), .ZN(_03909_ ) );
NOR3_X1 _11651_ ( .A1(_03905_ ), .A2(_03717_ ), .A3(_03909_ ), .ZN(_03910_ ) );
BUF_X4 _11652_ ( .A(_03903_ ), .Z(_03911_ ) );
INV_X1 _11653_ ( .A(_03911_ ), .ZN(_03912_ ) );
AOI21_X1 _11654_ ( .A(_03910_ ), .B1(_02069_ ), .B2(_03912_ ), .ZN(_03913_ ) );
XNOR2_X2 _11655_ ( .A(_03908_ ), .B(_02045_ ), .ZN(_03914_ ) );
INV_X1 _11656_ ( .A(_03914_ ), .ZN(_03915_ ) );
AND2_X1 _11657_ ( .A1(_03911_ ), .A2(_02069_ ), .ZN(_03916_ ) );
NOR2_X1 _11658_ ( .A1(_03911_ ), .A2(_02069_ ), .ZN(_03917_ ) );
NAND3_X2 _11659_ ( .A1(_03648_ ), .A2(_03668_ ), .A3(_03725_ ), .ZN(_03918_ ) );
INV_X1 _11660_ ( .A(\ID_EX_imm [0] ), .ZN(_03919_ ) );
NAND2_X1 _11661_ ( .A1(_03919_ ), .A2(\ID_EX_typ [4] ), .ZN(_03920_ ) );
NAND2_X2 _11662_ ( .A1(_03918_ ), .A2(_03920_ ), .ZN(_03921_ ) );
NOR2_X1 _11663_ ( .A1(_03921_ ), .A2(_03645_ ), .ZN(_03922_ ) );
NAND3_X1 _11664_ ( .A1(_03622_ ), .A2(_03642_ ), .A3(_03726_ ), .ZN(_03923_ ) );
NAND2_X1 _11665_ ( .A1(_02015_ ), .A2(\ID_EX_typ [4] ), .ZN(_03924_ ) );
AND3_X1 _11666_ ( .A1(_03923_ ), .A2(_02014_ ), .A3(_03924_ ), .ZN(_03925_ ) );
INV_X1 _11667_ ( .A(_03925_ ), .ZN(_03926_ ) );
NAND2_X1 _11668_ ( .A1(_03923_ ), .A2(_03924_ ), .ZN(_03927_ ) );
NAND2_X1 _11669_ ( .A1(_03927_ ), .A2(_02041_ ), .ZN(_03928_ ) );
AOI21_X1 _11670_ ( .A(_03922_ ), .B1(_03926_ ), .B2(_03928_ ), .ZN(_03929_ ) );
AOI21_X1 _11671_ ( .A(_02041_ ), .B1(_03923_ ), .B2(_03924_ ), .ZN(_03930_ ) );
OAI221_X1 _11672_ ( .A(_03915_ ), .B1(_03916_ ), .B2(_03917_ ), .C1(_03929_ ), .C2(_03930_ ), .ZN(_03931_ ) );
AOI21_X1 _11673_ ( .A(_03900_ ), .B1(_03913_ ), .B2(_03931_ ), .ZN(_03932_ ) );
AOI211_X1 _11674_ ( .A(_03895_ ), .B(_03932_ ), .C1(_02149_ ), .C2(_03874_ ), .ZN(_03933_ ) );
NAND3_X1 _11675_ ( .A1(_03878_ ), .A2(_02171_ ), .A3(_03881_ ), .ZN(_03934_ ) );
AOI21_X1 _11676_ ( .A(_03871_ ), .B1(_03933_ ), .B2(_03934_ ), .ZN(_03935_ ) );
INV_X1 _11677_ ( .A(_03838_ ), .ZN(_03936_ ) );
NOR3_X1 _11678_ ( .A1(_03834_ ), .A2(_03135_ ), .A3(_03936_ ), .ZN(_03937_ ) );
AND2_X1 _11679_ ( .A1(_03863_ ), .A2(_03292_ ), .ZN(_03938_ ) );
NOR2_X1 _11680_ ( .A1(_03863_ ), .A2(_03292_ ), .ZN(_03939_ ) );
OAI211_X1 _11681_ ( .A(_02202_ ), .B(_03868_ ), .C1(_03938_ ), .C2(_03939_ ), .ZN(_03940_ ) );
INV_X1 _11682_ ( .A(_03863_ ), .ZN(_03941_ ) );
OAI21_X1 _11683_ ( .A(_03940_ ), .B1(_03292_ ), .B2(_03941_ ), .ZN(_03942_ ) );
NAND2_X1 _11684_ ( .A1(_03942_ ), .A2(_03860_ ), .ZN(_03943_ ) );
NAND2_X1 _11685_ ( .A1(_03858_ ), .A2(_02272_ ), .ZN(_03944_ ) );
NAND2_X1 _11686_ ( .A1(_03943_ ), .A2(_03944_ ), .ZN(_03945_ ) );
INV_X1 _11687_ ( .A(_03854_ ), .ZN(_03946_ ) );
NOR3_X1 _11688_ ( .A1(_03859_ ), .A2(_03266_ ), .A3(_03946_ ), .ZN(_03947_ ) );
OAI21_X1 _11689_ ( .A(_03851_ ), .B1(_03945_ ), .B2(_03947_ ), .ZN(_03948_ ) );
NOR2_X1 _11690_ ( .A1(_03834_ ), .A2(_03839_ ), .ZN(_03949_ ) );
INV_X1 _11691_ ( .A(_03843_ ), .ZN(_03950_ ) );
NOR3_X1 _11692_ ( .A1(_03850_ ), .A2(_03188_ ), .A3(_03950_ ), .ZN(_03951_ ) );
AOI21_X1 _11693_ ( .A(_03214_ ), .B1(_03847_ ), .B2(_03848_ ), .ZN(_03952_ ) );
OAI21_X1 _11694_ ( .A(_03949_ ), .B1(_03951_ ), .B2(_03952_ ), .ZN(_03953_ ) );
INV_X1 _11695_ ( .A(_02309_ ), .ZN(_03954_ ) );
OR3_X1 _11696_ ( .A1(_03831_ ), .A2(_03954_ ), .A3(_03832_ ), .ZN(_03955_ ) );
NAND3_X1 _11697_ ( .A1(_03948_ ), .A2(_03953_ ), .A3(_03955_ ), .ZN(_03956_ ) );
NOR3_X2 _11698_ ( .A1(_03935_ ), .A2(_03937_ ), .A3(_03956_ ), .ZN(_03957_ ) );
XNOR2_X1 _11699_ ( .A(_03810_ ), .B(_01965_ ), .ZN(_03958_ ) );
OR4_X2 _11700_ ( .A1(_03790_ ), .A2(_03794_ ), .A3(_03798_ ), .A4(_03958_ ), .ZN(_03959_ ) );
OR3_X4 _11701_ ( .A1(_03959_ ), .A2(_03821_ ), .A3(_03807_ ), .ZN(_03960_ ) );
OAI211_X1 _11702_ ( .A(_03824_ ), .B(_03830_ ), .C1(_03957_ ), .C2(_03960_ ), .ZN(_03961_ ) );
NOR2_X1 _11703_ ( .A1(_03788_ ), .A2(_03789_ ), .ZN(_03962_ ) );
INV_X1 _11704_ ( .A(_03782_ ), .ZN(_03963_ ) );
NOR3_X1 _11705_ ( .A1(_03962_ ), .A2(_03033_ ), .A3(_03963_ ), .ZN(_03964_ ) );
OAI21_X1 _11706_ ( .A(_03779_ ), .B1(_03961_ ), .B2(_03964_ ), .ZN(_03965_ ) );
NAND2_X1 _11707_ ( .A1(_03775_ ), .A2(_02456_ ), .ZN(_03966_ ) );
OAI211_X1 _11708_ ( .A(_02432_ ), .B(_03771_ ), .C1(_03776_ ), .C2(_03777_ ), .ZN(_03967_ ) );
AOI21_X1 _11709_ ( .A(_03768_ ), .B1(_03966_ ), .B2(_03967_ ), .ZN(_03968_ ) );
AOI21_X1 _11710_ ( .A(_03968_ ), .B1(_03502_ ), .B2(_03762_ ), .ZN(_03969_ ) );
NAND3_X1 _11711_ ( .A1(_03767_ ), .A2(_02510_ ), .A3(_03755_ ), .ZN(_03970_ ) );
AND2_X1 _11712_ ( .A1(_03969_ ), .A2(_03970_ ), .ZN(_03971_ ) );
AOI21_X1 _11713_ ( .A(_03752_ ), .B1(_03965_ ), .B2(_03971_ ), .ZN(_03972_ ) );
INV_X1 _11714_ ( .A(_03972_ ), .ZN(_03973_ ) );
OR3_X1 _11715_ ( .A1(_03739_ ), .A2(_03732_ ), .A3(_03731_ ), .ZN(_03974_ ) );
OAI21_X1 _11716_ ( .A(_03974_ ), .B1(_03738_ ), .B2(_03737_ ), .ZN(_03975_ ) );
NAND2_X1 _11717_ ( .A1(_03975_ ), .A2(_03751_ ), .ZN(_03976_ ) );
NOR2_X1 _11718_ ( .A1(_03750_ ), .A2(_03749_ ), .ZN(_03977_ ) );
NAND2_X1 _11719_ ( .A1(_03741_ ), .A2(_03742_ ), .ZN(_03978_ ) );
NOR2_X1 _11720_ ( .A1(_03978_ ), .A2(_01732_ ), .ZN(_03979_ ) );
AOI21_X1 _11721_ ( .A(_03749_ ), .B1(_03977_ ), .B2(_03979_ ), .ZN(_03980_ ) );
AND3_X4 _11722_ ( .A1(_03973_ ), .A2(_03976_ ), .A3(_03980_ ), .ZN(_03981_ ) );
INV_X1 _11723_ ( .A(\ID_EX_typ [2] ), .ZN(_03982_ ) );
NOR3_X1 _11724_ ( .A1(_03982_ ), .A2(\ID_EX_typ [1] ), .A3(fanout_net_8 ), .ZN(_03983_ ) );
AND2_X4 _11725_ ( .A1(_03981_ ), .A2(_03983_ ), .ZN(_03984_ ) );
AND2_X1 _11726_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_8 ), .ZN(_03985_ ) );
AND2_X2 _11727_ ( .A1(_03985_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_03986_ ) );
INV_X1 _11728_ ( .A(_03986_ ), .ZN(_03987_ ) );
AND3_X1 _11729_ ( .A1(_02045_ ), .A2(_03695_ ), .A3(_03715_ ), .ZN(_03988_ ) );
INV_X1 _11730_ ( .A(_03988_ ), .ZN(_03989_ ) );
NOR2_X1 _11731_ ( .A1(_03669_ ), .A2(_03645_ ), .ZN(_03990_ ) );
INV_X1 _11732_ ( .A(_03990_ ), .ZN(_03991_ ) );
AND2_X1 _11733_ ( .A1(_03644_ ), .A2(_03991_ ), .ZN(_03992_ ) );
AOI21_X1 _11734_ ( .A(_03992_ ), .B1(_02014_ ), .B2(_03643_ ), .ZN(_03993_ ) );
OAI221_X2 _11735_ ( .A(_03989_ ), .B1(_03904_ ), .B2(_03691_ ), .C1(_03993_ ), .C2(_03719_ ), .ZN(_03994_ ) );
NAND3_X1 _11736_ ( .A1(_03691_ ), .A2(_02068_ ), .A3(_02067_ ), .ZN(_03995_ ) );
NAND3_X2 _11737_ ( .A1(_03994_ ), .A2(_03995_ ), .A3(_03423_ ), .ZN(_03996_ ) );
AND3_X1 _11738_ ( .A1(_03343_ ), .A2(_02171_ ), .A3(_03373_ ), .ZN(_03997_ ) );
AND3_X1 _11739_ ( .A1(_02118_ ), .A2(_03399_ ), .A3(_03419_ ), .ZN(_03998_ ) );
NAND2_X1 _11740_ ( .A1(_03398_ ), .A2(_03998_ ), .ZN(_03999_ ) );
OAI21_X1 _11741_ ( .A(_03999_ ), .B1(_03891_ ), .B2(_03397_ ), .ZN(_04000_ ) );
AOI221_X4 _11742_ ( .A(_03997_ ), .B1(_02149_ ), .B2(_03341_ ), .C1(_04000_ ), .C2(_03375_ ), .ZN(_04001_ ) );
AND2_X4 _11743_ ( .A1(_03996_ ), .A2(_04001_ ), .ZN(_04002_ ) );
INV_X4 _11744_ ( .A(_04002_ ), .ZN(_04003_ ) );
NAND3_X2 _11745_ ( .A1(_04003_ ), .A2(_03217_ ), .A3(_03319_ ), .ZN(_04004_ ) );
AND2_X1 _11746_ ( .A1(_03134_ ), .A2(_02332_ ), .ZN(_04005_ ) );
INV_X1 _11747_ ( .A(_04005_ ), .ZN(_04006_ ) );
NOR2_X1 _11748_ ( .A1(_04006_ ), .A2(_03163_ ), .ZN(_04007_ ) );
NOR2_X1 _11749_ ( .A1(_03212_ ), .A2(_03213_ ), .ZN(_04008_ ) );
INV_X1 _11750_ ( .A(_04008_ ), .ZN(_04009_ ) );
AND2_X1 _11751_ ( .A1(_03187_ ), .A2(_02380_ ), .ZN(_04010_ ) );
AND2_X1 _11752_ ( .A1(_03212_ ), .A2(_03213_ ), .ZN(_04011_ ) );
OAI21_X1 _11753_ ( .A(_04009_ ), .B1(_04010_ ), .B2(_04011_ ), .ZN(_04012_ ) );
OR3_X1 _11754_ ( .A1(_03137_ ), .A2(_04012_ ), .A3(_03163_ ), .ZN(_04013_ ) );
INV_X1 _11755_ ( .A(_03217_ ), .ZN(_04014_ ) );
NAND3_X1 _11756_ ( .A1(_03293_ ), .A2(_02202_ ), .A3(_03316_ ), .ZN(_04015_ ) );
NAND2_X1 _11757_ ( .A1(_03291_ ), .A2(_02225_ ), .ZN(_04016_ ) );
NAND2_X1 _11758_ ( .A1(_04015_ ), .A2(_04016_ ), .ZN(_04017_ ) );
NAND2_X1 _11759_ ( .A1(_04017_ ), .A2(_03268_ ), .ZN(_04018_ ) );
NAND3_X1 _11760_ ( .A1(_02272_ ), .A2(_03219_ ), .A3(_03239_ ), .ZN(_04019_ ) );
AND2_X1 _11761_ ( .A1(_03265_ ), .A2(_02249_ ), .ZN(_04020_ ) );
NAND2_X1 _11762_ ( .A1(_03242_ ), .A2(_04020_ ), .ZN(_04021_ ) );
AND3_X2 _11763_ ( .A1(_04018_ ), .A2(_04019_ ), .A3(_04021_ ), .ZN(_04022_ ) );
OAI21_X2 _11764_ ( .A(_04013_ ), .B1(_04014_ ), .B2(_04022_ ), .ZN(_04023_ ) );
AOI211_X2 _11765_ ( .A(_04007_ ), .B(_04023_ ), .C1(_02309_ ), .C2(_03162_ ), .ZN(_04024_ ) );
AND2_X2 _11766_ ( .A1(_04004_ ), .A2(_04024_ ), .ZN(_04025_ ) );
AND2_X1 _11767_ ( .A1(_03111_ ), .A2(_03619_ ), .ZN(_04026_ ) );
INV_X1 _11768_ ( .A(_04026_ ), .ZN(_04027_ ) );
OR2_X2 _11769_ ( .A1(_04025_ ), .A2(_04027_ ), .ZN(_04028_ ) );
INV_X1 _11770_ ( .A(_02571_ ), .ZN(_04029_ ) );
NOR2_X1 _11771_ ( .A1(_04029_ ), .A2(_03571_ ), .ZN(_04030_ ) );
NOR2_X1 _11772_ ( .A1(_01732_ ), .A2(_03549_ ), .ZN(_04031_ ) );
AOI21_X1 _11773_ ( .A(_04030_ ), .B1(_03572_ ), .B2(_04031_ ), .ZN(_04032_ ) );
NAND4_X1 _11774_ ( .A1(_03479_ ), .A2(_02432_ ), .A3(_03447_ ), .A4(_03449_ ), .ZN(_04033_ ) );
NAND2_X1 _11775_ ( .A1(_04033_ ), .A2(_03478_ ), .ZN(_04034_ ) );
AND3_X1 _11776_ ( .A1(_04034_ ), .A2(_03503_ ), .A3(_03526_ ), .ZN(_04035_ ) );
NOR2_X1 _11777_ ( .A1(_03501_ ), .A2(_03763_ ), .ZN(_04036_ ) );
NOR2_X1 _11778_ ( .A1(_03525_ ), .A2(_02514_ ), .ZN(_04037_ ) );
AND2_X1 _11779_ ( .A1(_03503_ ), .A2(_04037_ ), .ZN(_04038_ ) );
NOR3_X1 _11780_ ( .A1(_04035_ ), .A2(_04036_ ), .A3(_04038_ ), .ZN(_04039_ ) );
AND2_X1 _11781_ ( .A1(_03573_ ), .A2(_03618_ ), .ZN(_04040_ ) );
INV_X1 _11782_ ( .A(_04040_ ), .ZN(_04041_ ) );
OAI21_X1 _11783_ ( .A(_04032_ ), .B1(_04039_ ), .B2(_04041_ ), .ZN(_04042_ ) );
AND3_X1 _11784_ ( .A1(_03738_ ), .A2(_03593_ ), .A3(_03574_ ), .ZN(_04043_ ) );
NOR2_X1 _11785_ ( .A1(_03616_ ), .A2(_03732_ ), .ZN(_04044_ ) );
INV_X1 _11786_ ( .A(_04044_ ), .ZN(_04045_ ) );
OR2_X1 _11787_ ( .A1(_03594_ ), .A2(_03738_ ), .ZN(_04046_ ) );
AOI21_X1 _11788_ ( .A(_04043_ ), .B1(_04045_ ), .B2(_04046_ ), .ZN(_04047_ ) );
AND2_X1 _11789_ ( .A1(_02952_ ), .A2(_01965_ ), .ZN(_04048_ ) );
INV_X1 _11790_ ( .A(_04048_ ), .ZN(_04049_ ) );
AND2_X1 _11791_ ( .A1(_02921_ ), .A2(_01942_ ), .ZN(_04050_ ) );
NOR2_X1 _11792_ ( .A1(_02921_ ), .A2(_01942_ ), .ZN(_04051_ ) );
NOR3_X1 _11793_ ( .A1(_04049_ ), .A2(_04050_ ), .A3(_04051_ ), .ZN(_04052_ ) );
OAI211_X1 _11794_ ( .A(_02978_ ), .B(_03006_ ), .C1(_04052_ ), .C2(_04050_ ), .ZN(_04053_ ) );
NAND3_X1 _11795_ ( .A1(_02974_ ), .A2(_01918_ ), .A3(_02975_ ), .ZN(_04054_ ) );
NAND3_X1 _11796_ ( .A1(_02978_ ), .A2(_01895_ ), .A3(_03004_ ), .ZN(_04055_ ) );
AND3_X2 _11797_ ( .A1(_04053_ ), .A2(_04054_ ), .A3(_04055_ ), .ZN(_04056_ ) );
NOR2_X1 _11798_ ( .A1(_04056_ ), .A2(_03110_ ), .ZN(_04057_ ) );
AND2_X1 _11799_ ( .A1(_03032_ ), .A2(_01793_ ), .ZN(_04058_ ) );
AND2_X1 _11800_ ( .A1(_03059_ ), .A2(_04058_ ), .ZN(_04059_ ) );
AOI21_X1 _11801_ ( .A(_04059_ ), .B1(_01816_ ), .B2(_03057_ ), .ZN(_04060_ ) );
INV_X1 _11802_ ( .A(_04060_ ), .ZN(_04061_ ) );
NAND3_X1 _11803_ ( .A1(_03109_ ), .A2(_01869_ ), .A3(_03083_ ), .ZN(_04062_ ) );
INV_X1 _11804_ ( .A(_03108_ ), .ZN(_04063_ ) );
OAI21_X1 _11805_ ( .A(_04062_ ), .B1(_02403_ ), .B2(_04063_ ), .ZN(_04064_ ) );
AND2_X2 _11806_ ( .A1(_03060_ ), .A2(_04064_ ), .ZN(_04065_ ) );
NOR3_X1 _11807_ ( .A1(_04057_ ), .A2(_04061_ ), .A3(_04065_ ), .ZN(_04066_ ) );
INV_X1 _11808_ ( .A(_04066_ ), .ZN(_04067_ ) );
AOI221_X4 _11809_ ( .A(_04042_ ), .B1(_03573_ ), .B2(_04047_ ), .C1(_04067_ ), .C2(_03619_ ), .ZN(_04068_ ) );
AOI21_X1 _11810_ ( .A(_03987_ ), .B1(_04028_ ), .B2(_04068_ ), .ZN(_04069_ ) );
AND2_X2 _11811_ ( .A1(_03722_ ), .A2(\ID_EX_typ [2] ), .ZN(_04070_ ) );
AND3_X1 _11812_ ( .A1(_04028_ ), .A2(_04068_ ), .A3(_04070_ ), .ZN(_04071_ ) );
OR4_X4 _11813_ ( .A1(_03984_ ), .A2(_04069_ ), .A3(_03723_ ), .A4(_04071_ ), .ZN(_04072_ ) );
INV_X1 _11814_ ( .A(\ID_EX_typ [1] ), .ZN(_04073_ ) );
NOR2_X1 _11815_ ( .A1(_04073_ ), .A2(fanout_net_8 ), .ZN(_04074_ ) );
AND2_X2 _11816_ ( .A1(_04074_ ), .A2(_03982_ ), .ZN(_04075_ ) );
INV_X1 _11817_ ( .A(_04075_ ), .ZN(_04076_ ) );
NOR2_X1 _11818_ ( .A1(_03981_ ), .A2(_04076_ ), .ZN(_04077_ ) );
OAI221_X2 _11819_ ( .A(_02861_ ), .B1(_03721_ ), .B2(_03724_ ), .C1(_04072_ ), .C2(_04077_ ), .ZN(_04078_ ) );
AND4_X1 _11820_ ( .A1(_03217_ ), .A2(_03720_ ), .A3(_03319_ ), .A4(_03423_ ), .ZN(_04079_ ) );
NAND3_X1 _11821_ ( .A1(_03111_ ), .A2(_04079_ ), .A3(_03619_ ), .ZN(_04080_ ) );
NAND2_X1 _11822_ ( .A1(_04080_ ), .A2(_02860_ ), .ZN(_04081_ ) );
AOI21_X1 _11823_ ( .A(_02858_ ), .B1(_04078_ ), .B2(_04081_ ), .ZN(_04082_ ) );
AND2_X4 _11824_ ( .A1(_04078_ ), .A2(_04081_ ), .ZN(_04083_ ) );
BUF_X8 _11825_ ( .A(_04083_ ), .Z(_04084_ ) );
AOI211_X1 _11826_ ( .A(fanout_net_10 ), .B(_04082_ ), .C1(_02831_ ), .C2(_04084_ ), .ZN(_04085_ ) );
INV_X1 _11827_ ( .A(fanout_net_10 ), .ZN(_04086_ ) );
XNOR2_X1 _11828_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_04087_ ) );
AND2_X1 _11829_ ( .A1(_02661_ ), .A2(_04087_ ), .ZN(_04088_ ) );
XNOR2_X1 _11830_ ( .A(fanout_net_7 ), .B(\ID_EX_csr [1] ), .ZN(_04089_ ) );
AND2_X1 _11831_ ( .A1(_02662_ ), .A2(_04089_ ), .ZN(_04090_ ) );
XNOR2_X1 _11832_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_04091_ ) );
XNOR2_X1 _11833_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_04092_ ) );
AND2_X1 _11834_ ( .A1(_04091_ ), .A2(_04092_ ), .ZN(_04093_ ) );
AND2_X1 _11835_ ( .A1(_02653_ ), .A2(_02656_ ), .ZN(_04094_ ) );
AND4_X1 _11836_ ( .A1(_04088_ ), .A2(_04090_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04095_ ) );
XOR2_X1 _11837_ ( .A(\EX_LS_dest_csreg_mem [8] ), .B(\ID_EX_csr [8] ), .Z(_04096_ ) );
NOR2_X1 _11838_ ( .A1(_02649_ ), .A2(_04096_ ), .ZN(_04097_ ) );
XNOR2_X1 _11839_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_04098_ ) );
XOR2_X1 _11840_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .Z(_04099_ ) );
INV_X1 _11841_ ( .A(_04099_ ), .ZN(_04100_ ) );
NAND4_X1 _11842_ ( .A1(_04095_ ), .A2(_04097_ ), .A3(_04098_ ), .A4(_04100_ ), .ZN(_04101_ ) );
NOR2_X1 _11843_ ( .A1(_04101_ ), .A2(_01677_ ), .ZN(_04102_ ) );
NAND2_X1 _11844_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [30] ), .ZN(_04103_ ) );
AND4_X1 _11845_ ( .A1(\ID_EX_csr [4] ), .A2(_02668_ ), .A3(_02671_ ), .A4(_02672_ ), .ZN(_04104_ ) );
NAND2_X1 _11846_ ( .A1(_04104_ ), .A2(_02667_ ), .ZN(_04105_ ) );
BUF_X2 _11847_ ( .A(_02696_ ), .Z(_04106_ ) );
BUF_X4 _11848_ ( .A(_02700_ ), .Z(_04107_ ) );
NAND4_X1 _11849_ ( .A1(_04106_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][30] ), .A4(_04107_ ), .ZN(_04108_ ) );
AND2_X1 _11850_ ( .A1(_04105_ ), .A2(_04108_ ), .ZN(_04109_ ) );
AND4_X1 _11851_ ( .A1(_02694_ ), .A2(_02671_ ), .A3(_02693_ ), .A4(_02672_ ), .ZN(_04110_ ) );
BUF_X4 _11852_ ( .A(_04110_ ), .Z(_04111_ ) );
BUF_X4 _11853_ ( .A(_02700_ ), .Z(_04112_ ) );
BUF_X4 _11854_ ( .A(_04112_ ), .Z(_04113_ ) );
NAND3_X1 _11855_ ( .A1(_04111_ ), .A2(\mepc [30] ), .A3(_04113_ ), .ZN(_04114_ ) );
BUF_X4 _11856_ ( .A(_02701_ ), .Z(_04115_ ) );
NAND4_X1 _11857_ ( .A1(_02678_ ), .A2(_02683_ ), .A3(\mtvec [30] ), .A4(_04115_ ), .ZN(_04116_ ) );
BUF_X2 _11858_ ( .A(_02702_ ), .Z(_04117_ ) );
NAND4_X1 _11859_ ( .A1(_02683_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_04115_ ), .A4(_04117_ ), .ZN(_04118_ ) );
NAND4_X1 _11860_ ( .A1(_04109_ ), .A2(_04114_ ), .A3(_04116_ ), .A4(_04118_ ), .ZN(_04119_ ) );
CLKBUF_X2 _11861_ ( .A(_04101_ ), .Z(_04120_ ) );
CLKBUF_X2 _11862_ ( .A(_01677_ ), .Z(_04121_ ) );
OAI21_X1 _11863_ ( .A(_04119_ ), .B1(_04120_ ), .B2(_04121_ ), .ZN(_04122_ ) );
AOI21_X1 _11864_ ( .A(_04086_ ), .B1(_04103_ ), .B2(_04122_ ), .ZN(_04123_ ) );
OAI21_X1 _11865_ ( .A(_02840_ ), .B1(_04085_ ), .B2(_04123_ ), .ZN(_04124_ ) );
AOI221_X1 _11866_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_02719_ ), .C1(_02839_ ), .C2(_04124_ ), .ZN(_00120_ ) );
BUF_X4 _11867_ ( .A(_02578_ ), .Z(_04125_ ) );
NAND2_X1 _11868_ ( .A1(_02823_ ), .A2(_02824_ ), .ZN(_04126_ ) );
XNOR2_X1 _11869_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .ZN(_04127_ ) );
XOR2_X1 _11870_ ( .A(_04126_ ), .B(_04127_ ), .Z(_04128_ ) );
INV_X1 _11871_ ( .A(_04128_ ), .ZN(_04129_ ) );
OAI21_X1 _11872_ ( .A(_01649_ ), .B1(_04129_ ), .B2(fanout_net_8 ), .ZN(_04130_ ) );
AOI21_X1 _11873_ ( .A(_04130_ ), .B1(_02618_ ), .B2(fanout_net_8 ), .ZN(_04131_ ) );
NOR2_X1 _11874_ ( .A1(_02665_ ), .A2(\EX_LS_result_csreg_mem [29] ), .ZN(_04132_ ) );
BUF_X2 _11875_ ( .A(_02680_ ), .Z(_04133_ ) );
BUF_X2 _11876_ ( .A(_02686_ ), .Z(_04134_ ) );
NAND4_X1 _11877_ ( .A1(_02677_ ), .A2(_04133_ ), .A3(\mtvec [29] ), .A4(_04134_ ), .ZN(_04135_ ) );
BUF_X4 _11878_ ( .A(_02702_ ), .Z(_04136_ ) );
NAND4_X1 _11879_ ( .A1(_04133_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_02687_ ), .A4(_04136_ ), .ZN(_04137_ ) );
BUF_X4 _11880_ ( .A(_02695_ ), .Z(_04138_ ) );
NAND4_X1 _11881_ ( .A1(_02690_ ), .A2(_04138_ ), .A3(\mepc [29] ), .A4(_02687_ ), .ZN(_04139_ ) );
BUF_X4 _11882_ ( .A(_02707_ ), .Z(_04140_ ) );
NAND4_X1 _11883_ ( .A1(_04138_ ), .A2(_04140_ ), .A3(\mycsreg.CSReg[3][29] ), .A4(_02687_ ), .ZN(_04141_ ) );
NAND4_X1 _11884_ ( .A1(_04135_ ), .A2(_04137_ ), .A3(_04139_ ), .A4(_04141_ ), .ZN(_04142_ ) );
AOI211_X1 _11885_ ( .A(_02675_ ), .B(_04142_ ), .C1(_02714_ ), .C2(_02716_ ), .ZN(_04143_ ) );
NOR2_X1 _11886_ ( .A1(_04132_ ), .A2(_04143_ ), .ZN(_04144_ ) );
AND4_X1 _11887_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_04145_ ) );
AND2_X1 _11888_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_04146_ ) );
AND4_X1 _11889_ ( .A1(\ID_EX_pc [13] ), .A2(_04145_ ), .A3(\ID_EX_pc [12] ), .A4(_04146_ ), .ZN(_04147_ ) );
AND2_X1 _11890_ ( .A1(_02847_ ), .A2(_04147_ ), .ZN(_04148_ ) );
AND4_X1 _11891_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_04149_ ) );
AND2_X1 _11892_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_04150_ ) );
AND4_X1 _11893_ ( .A1(\ID_EX_pc [21] ), .A2(_04149_ ), .A3(\ID_EX_pc [20] ), .A4(_04150_ ), .ZN(_04151_ ) );
NAND2_X1 _11894_ ( .A1(_04148_ ), .A2(_04151_ ), .ZN(_04152_ ) );
INV_X1 _11895_ ( .A(\ID_EX_pc [27] ), .ZN(_04153_ ) );
INV_X1 _11896_ ( .A(\ID_EX_pc [26] ), .ZN(_04154_ ) );
NOR3_X1 _11897_ ( .A1(_04152_ ), .A2(_04153_ ), .A3(_04154_ ), .ZN(_04155_ ) );
NAND2_X1 _11898_ ( .A1(_04155_ ), .A2(\ID_EX_pc [28] ), .ZN(_04156_ ) );
XNOR2_X1 _11899_ ( .A(_04156_ ), .B(\ID_EX_pc [29] ), .ZN(_04157_ ) );
MUX2_X1 _11900_ ( .A(_04157_ ), .B(_04129_ ), .S(_04083_ ), .Z(_04158_ ) );
BUF_X4 _11901_ ( .A(_04086_ ), .Z(_04159_ ) );
MUX2_X2 _11902_ ( .A(_04144_ ), .B(_04158_ ), .S(_04159_ ), .Z(_04160_ ) );
BUF_X4 _11903_ ( .A(_02840_ ), .Z(_04161_ ) );
AOI211_X1 _11904_ ( .A(_04125_ ), .B(_04131_ ), .C1(_04160_ ), .C2(_04161_ ), .ZN(_04162_ ) );
BUF_X4 _11905_ ( .A(_04125_ ), .Z(_04163_ ) );
INV_X1 _11906_ ( .A(_04144_ ), .ZN(_04164_ ) );
AOI211_X1 _11907_ ( .A(fanout_net_2 ), .B(_04162_ ), .C1(_04163_ ), .C2(_04164_ ), .ZN(_00121_ ) );
NOR2_X1 _11908_ ( .A1(_02664_ ), .A2(_02674_ ), .ZN(_04165_ ) );
AND2_X1 _11909_ ( .A1(_02669_ ), .A2(_02707_ ), .ZN(_04166_ ) );
INV_X1 _11910_ ( .A(_04166_ ), .ZN(_04167_ ) );
BUF_X4 _11911_ ( .A(_04167_ ), .Z(_04168_ ) );
BUF_X2 _11912_ ( .A(_02677_ ), .Z(_04169_ ) );
BUF_X2 _11913_ ( .A(_02686_ ), .Z(_04170_ ) );
NAND4_X1 _11914_ ( .A1(_04169_ ), .A2(_04133_ ), .A3(\mtvec [20] ), .A4(_04170_ ), .ZN(_04171_ ) );
BUF_X4 _11915_ ( .A(_02696_ ), .Z(_04172_ ) );
BUF_X2 _11916_ ( .A(_02707_ ), .Z(_04173_ ) );
BUF_X4 _11917_ ( .A(_02686_ ), .Z(_04174_ ) );
NAND4_X1 _11918_ ( .A1(_04172_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][20] ), .A4(_04174_ ), .ZN(_04175_ ) );
NAND4_X1 _11919_ ( .A1(_04133_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_04134_ ), .A4(_04136_ ), .ZN(_04176_ ) );
NAND4_X1 _11920_ ( .A1(_02690_ ), .A2(_04138_ ), .A3(\mepc [20] ), .A4(_04134_ ), .ZN(_04177_ ) );
AND4_X1 _11921_ ( .A1(_04171_ ), .A2(_04175_ ), .A3(_04176_ ), .A4(_04177_ ), .ZN(_04178_ ) );
NAND3_X1 _11922_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04178_ ), .ZN(_04179_ ) );
AND3_X1 _11923_ ( .A1(_04097_ ), .A2(_01676_ ), .A3(_04098_ ), .ZN(_04180_ ) );
AND3_X2 _11924_ ( .A1(_04180_ ), .A2(_04088_ ), .A3(_04090_ ), .ZN(_04181_ ) );
INV_X1 _11925_ ( .A(\EX_LS_result_csreg_mem [20] ), .ZN(_04182_ ) );
AND3_X2 _11926_ ( .A1(_04093_ ), .A2(_04094_ ), .A3(_04100_ ), .ZN(_04183_ ) );
NAND3_X1 _11927_ ( .A1(_04181_ ), .A2(_04182_ ), .A3(_04183_ ), .ZN(_04184_ ) );
AND2_X1 _11928_ ( .A1(_04179_ ), .A2(_04184_ ), .ZN(_04185_ ) );
INV_X1 _11929_ ( .A(_04185_ ), .ZN(_04186_ ) );
NAND3_X1 _11930_ ( .A1(_02847_ ), .A2(_04147_ ), .A3(_04150_ ), .ZN(_04187_ ) );
XNOR2_X1 _11931_ ( .A(_04187_ ), .B(\ID_EX_pc [20] ), .ZN(_04188_ ) );
BUF_X4 _11932_ ( .A(_04078_ ), .Z(_04189_ ) );
BUF_X4 _11933_ ( .A(_04081_ ), .Z(_04190_ ) );
AOI21_X1 _11934_ ( .A(_04188_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04191_ ) );
BUF_X4 _11935_ ( .A(_04084_ ), .Z(_04192_ ) );
XNOR2_X1 _11936_ ( .A(_02792_ ), .B(_02795_ ), .ZN(_04193_ ) );
AOI211_X1 _11937_ ( .A(fanout_net_10 ), .B(_04191_ ), .C1(_04192_ ), .C2(_04193_ ), .ZN(_04194_ ) );
AND3_X1 _11938_ ( .A1(_04179_ ), .A2(fanout_net_10 ), .A3(_04184_ ), .ZN(_04195_ ) );
OAI21_X1 _11939_ ( .A(_01654_ ), .B1(_04194_ ), .B2(_04195_ ), .ZN(_04196_ ) );
AOI21_X1 _11940_ ( .A(_02720_ ), .B1(_04193_ ), .B2(_02833_ ), .ZN(_04197_ ) );
OAI21_X1 _11941_ ( .A(_04197_ ), .B1(_02592_ ), .B2(_02835_ ), .ZN(_04198_ ) );
AND2_X1 _11942_ ( .A1(_04198_ ), .A2(_02838_ ), .ZN(_04199_ ) );
AOI221_X1 _11943_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04186_ ), .C1(_04196_ ), .C2(_04199_ ), .ZN(_00122_ ) );
BUF_X4 _11944_ ( .A(_04140_ ), .Z(_04200_ ) );
NAND4_X1 _11945_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][19] ), .A4(_02688_ ), .ZN(_04201_ ) );
NAND3_X1 _11946_ ( .A1(_04111_ ), .A2(\mepc [19] ), .A3(_02688_ ), .ZN(_04202_ ) );
BUF_X4 _11947_ ( .A(_02677_ ), .Z(_04203_ ) );
BUF_X2 _11948_ ( .A(_02681_ ), .Z(_04204_ ) );
BUF_X4 _11949_ ( .A(_02687_ ), .Z(_04205_ ) );
NAND4_X1 _11950_ ( .A1(_04203_ ), .A2(_04204_ ), .A3(\mtvec [19] ), .A4(_04205_ ), .ZN(_04206_ ) );
NAND4_X1 _11951_ ( .A1(_04168_ ), .A2(_04201_ ), .A3(_04202_ ), .A4(_04206_ ), .ZN(_04207_ ) );
AND4_X1 _11952_ ( .A1(\mycsreg.CSReg[0][19] ), .A2(_04204_ ), .A3(_02688_ ), .A4(_04117_ ), .ZN(_04208_ ) );
OAI21_X1 _11953_ ( .A(_02665_ ), .B1(_04207_ ), .B2(_04208_ ), .ZN(_04209_ ) );
NAND3_X1 _11954_ ( .A1(_02715_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_02717_ ), .ZN(_04210_ ) );
AND2_X1 _11955_ ( .A1(_04209_ ), .A2(_04210_ ), .ZN(_04211_ ) );
BUF_X4 _11956_ ( .A(_01653_ ), .Z(_04212_ ) );
NAND3_X1 _11957_ ( .A1(_02847_ ), .A2(\ID_EX_pc [18] ), .A3(_04147_ ), .ZN(_04213_ ) );
XNOR2_X1 _11958_ ( .A(_04213_ ), .B(\ID_EX_pc [19] ), .ZN(_04214_ ) );
AOI21_X1 _11959_ ( .A(_04214_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04215_ ) );
INV_X1 _11960_ ( .A(_02778_ ), .ZN(_04216_ ) );
OAI21_X1 _11961_ ( .A(_02782_ ), .B1(_02768_ ), .B2(_02775_ ), .ZN(_04217_ ) );
AOI21_X1 _11962_ ( .A(_04216_ ), .B1(_04217_ ), .B2(_02789_ ), .ZN(_04218_ ) );
OR2_X1 _11963_ ( .A1(_04218_ ), .A2(_02784_ ), .ZN(_04219_ ) );
XNOR2_X1 _11964_ ( .A(_04219_ ), .B(_02777_ ), .ZN(_04220_ ) );
AOI211_X1 _11965_ ( .A(fanout_net_10 ), .B(_04215_ ), .C1(_04192_ ), .C2(_04220_ ), .ZN(_04221_ ) );
NAND2_X1 _11966_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_04222_ ) );
AOI21_X1 _11967_ ( .A(_04159_ ), .B1(_04209_ ), .B2(_04222_ ), .ZN(_04223_ ) );
OAI21_X1 _11968_ ( .A(_04212_ ), .B1(_04221_ ), .B2(_04223_ ), .ZN(_04224_ ) );
BUF_X4 _11969_ ( .A(_02578_ ), .Z(_04225_ ) );
NAND2_X1 _11970_ ( .A1(_02599_ ), .A2(fanout_net_8 ), .ZN(_04226_ ) );
BUF_X2 _11971_ ( .A(_02832_ ), .Z(_04227_ ) );
AOI21_X1 _11972_ ( .A(_01653_ ), .B1(_04220_ ), .B2(_04227_ ), .ZN(_04228_ ) );
AOI21_X1 _11973_ ( .A(_04225_ ), .B1(_04226_ ), .B2(_04228_ ), .ZN(_04229_ ) );
AOI221_X1 _11974_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04211_ ), .C1(_04224_ ), .C2(_04229_ ), .ZN(_00123_ ) );
AND4_X1 _11975_ ( .A1(\mtvec [18] ), .A2(_02678_ ), .A3(_04204_ ), .A4(_02688_ ), .ZN(_04230_ ) );
BUF_X4 _11976_ ( .A(_04138_ ), .Z(_04231_ ) );
NAND4_X1 _11977_ ( .A1(_02691_ ), .A2(_04231_ ), .A3(\mepc [18] ), .A4(_02688_ ), .ZN(_04232_ ) );
BUF_X4 _11978_ ( .A(_02680_ ), .Z(_04233_ ) );
NAND4_X1 _11979_ ( .A1(_04233_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_04174_ ), .A4(_04136_ ), .ZN(_04234_ ) );
NAND4_X1 _11980_ ( .A1(_04172_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][18] ), .A4(_04174_ ), .ZN(_04235_ ) );
AND2_X1 _11981_ ( .A1(_04234_ ), .A2(_04235_ ), .ZN(_04236_ ) );
NAND3_X1 _11982_ ( .A1(_04168_ ), .A2(_04232_ ), .A3(_04236_ ), .ZN(_04237_ ) );
OAI21_X1 _11983_ ( .A(_02665_ ), .B1(_04230_ ), .B2(_04237_ ), .ZN(_04238_ ) );
NAND3_X1 _11984_ ( .A1(_02715_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_02717_ ), .ZN(_04239_ ) );
AND2_X1 _11985_ ( .A1(_04238_ ), .A2(_04239_ ), .ZN(_04240_ ) );
INV_X1 _11986_ ( .A(\ID_EX_pc [18] ), .ZN(_04241_ ) );
XNOR2_X1 _11987_ ( .A(_04148_ ), .B(_04241_ ), .ZN(_04242_ ) );
AOI21_X1 _11988_ ( .A(_04242_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04243_ ) );
NAND2_X1 _11989_ ( .A1(_04217_ ), .A2(_02789_ ), .ZN(_04244_ ) );
XNOR2_X1 _11990_ ( .A(_04244_ ), .B(_04216_ ), .ZN(_04245_ ) );
INV_X1 _11991_ ( .A(_04245_ ), .ZN(_04246_ ) );
AOI211_X1 _11992_ ( .A(fanout_net_10 ), .B(_04243_ ), .C1(_04192_ ), .C2(_04246_ ), .ZN(_04247_ ) );
NAND2_X1 _11993_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_04248_ ) );
AOI21_X1 _11994_ ( .A(_04159_ ), .B1(_04238_ ), .B2(_04248_ ), .ZN(_04249_ ) );
OAI21_X1 _11995_ ( .A(_04212_ ), .B1(_04247_ ), .B2(_04249_ ), .ZN(_04250_ ) );
AOI21_X1 _11996_ ( .A(_02720_ ), .B1(_04246_ ), .B2(_02833_ ), .ZN(_04251_ ) );
OAI21_X1 _11997_ ( .A(_04251_ ), .B1(_02601_ ), .B2(_02835_ ), .ZN(_04252_ ) );
AND2_X1 _11998_ ( .A1(_04252_ ), .A2(_02838_ ), .ZN(_04253_ ) );
AOI221_X1 _11999_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04240_ ), .C1(_04250_ ), .C2(_04253_ ), .ZN(_00124_ ) );
NAND4_X1 _12000_ ( .A1(_04169_ ), .A2(_04233_ ), .A3(\mtvec [17] ), .A4(_02701_ ), .ZN(_04254_ ) );
NAND4_X1 _12001_ ( .A1(_04233_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_02709_ ), .A4(_02703_ ), .ZN(_04255_ ) );
BUF_X4 _12002_ ( .A(_02690_ ), .Z(_04256_ ) );
NAND4_X1 _12003_ ( .A1(_04256_ ), .A2(_02697_ ), .A3(\mepc [17] ), .A4(_04170_ ), .ZN(_04257_ ) );
NAND4_X1 _12004_ ( .A1(_04172_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][17] ), .A4(_04174_ ), .ZN(_04258_ ) );
AND4_X1 _12005_ ( .A1(_04254_ ), .A2(_04255_ ), .A3(_04257_ ), .A4(_04258_ ), .ZN(_04259_ ) );
NAND3_X1 _12006_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04259_ ), .ZN(_04260_ ) );
NAND3_X1 _12007_ ( .A1(_04180_ ), .A2(_04088_ ), .A3(_04090_ ), .ZN(_04261_ ) );
CLKBUF_X2 _12008_ ( .A(_04261_ ), .Z(_04262_ ) );
NAND3_X1 _12009_ ( .A1(_04093_ ), .A2(_04094_ ), .A3(_04100_ ), .ZN(_04263_ ) );
CLKBUF_X2 _12010_ ( .A(_04263_ ), .Z(_04264_ ) );
OR3_X1 _12011_ ( .A1(_04262_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_04264_ ), .ZN(_04265_ ) );
AND2_X1 _12012_ ( .A1(_04260_ ), .A2(_04265_ ), .ZN(_04266_ ) );
INV_X1 _12013_ ( .A(_04266_ ), .ZN(_04267_ ) );
INV_X4 _12014_ ( .A(_04083_ ), .ZN(_04268_ ) );
AND3_X1 _12015_ ( .A1(_04146_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_04269_ ) );
AND2_X1 _12016_ ( .A1(_02847_ ), .A2(_04269_ ), .ZN(_04270_ ) );
NAND3_X1 _12017_ ( .A1(_04270_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_04271_ ) );
INV_X1 _12018_ ( .A(\ID_EX_pc [16] ), .ZN(_04272_ ) );
NOR2_X1 _12019_ ( .A1(_04271_ ), .A2(_04272_ ), .ZN(_04273_ ) );
XNOR2_X1 _12020_ ( .A(_04273_ ), .B(\ID_EX_pc [17] ), .ZN(_04274_ ) );
AND2_X2 _12021_ ( .A1(_04268_ ), .A2(_04274_ ), .ZN(_04275_ ) );
AND2_X1 _12022_ ( .A1(_02776_ ), .A2(_02780_ ), .ZN(_04276_ ) );
OR2_X1 _12023_ ( .A1(_04276_ ), .A2(_02787_ ), .ZN(_04277_ ) );
XNOR2_X1 _12024_ ( .A(_04277_ ), .B(_02781_ ), .ZN(_04278_ ) );
AOI211_X2 _12025_ ( .A(fanout_net_10 ), .B(_04275_ ), .C1(_04192_ ), .C2(_04278_ ), .ZN(_04279_ ) );
NAND3_X1 _12026_ ( .A1(_04260_ ), .A2(fanout_net_10 ), .A3(_04265_ ), .ZN(_04280_ ) );
INV_X1 _12027_ ( .A(_04280_ ), .ZN(_04281_ ) );
OAI21_X1 _12028_ ( .A(_04212_ ), .B1(_04279_ ), .B2(_04281_ ), .ZN(_04282_ ) );
BUF_X4 _12029_ ( .A(_02578_ ), .Z(_04283_ ) );
NAND2_X1 _12030_ ( .A1(_02603_ ), .A2(fanout_net_8 ), .ZN(_04284_ ) );
AOI21_X1 _12031_ ( .A(_01653_ ), .B1(_04278_ ), .B2(_04227_ ), .ZN(_04285_ ) );
AOI21_X1 _12032_ ( .A(_04283_ ), .B1(_04284_ ), .B2(_04285_ ), .ZN(_04286_ ) );
AOI221_X1 _12033_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04267_ ), .C1(_04282_ ), .C2(_04286_ ), .ZN(_00125_ ) );
NAND4_X1 _12034_ ( .A1(_04169_ ), .A2(_04233_ ), .A3(\mtvec [16] ), .A4(_02709_ ), .ZN(_04287_ ) );
NAND4_X1 _12035_ ( .A1(_04233_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_02709_ ), .A4(_04136_ ), .ZN(_04288_ ) );
NAND4_X1 _12036_ ( .A1(_04256_ ), .A2(_02697_ ), .A3(\mepc [16] ), .A4(_04170_ ), .ZN(_04289_ ) );
NAND4_X1 _12037_ ( .A1(_04172_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][16] ), .A4(_04174_ ), .ZN(_04290_ ) );
AND4_X1 _12038_ ( .A1(_04287_ ), .A2(_04288_ ), .A3(_04289_ ), .A4(_04290_ ), .ZN(_04291_ ) );
NAND3_X1 _12039_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04291_ ), .ZN(_04292_ ) );
OR3_X1 _12040_ ( .A1(_04262_ ), .A2(\EX_LS_result_csreg_mem [16] ), .A3(_04264_ ), .ZN(_04293_ ) );
AND2_X1 _12041_ ( .A1(_04292_ ), .A2(_04293_ ), .ZN(_04294_ ) );
INV_X1 _12042_ ( .A(_04294_ ), .ZN(_04295_ ) );
XNOR2_X1 _12043_ ( .A(_04271_ ), .B(\ID_EX_pc [16] ), .ZN(_04296_ ) );
AOI21_X1 _12044_ ( .A(_04296_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04297_ ) );
XOR2_X1 _12045_ ( .A(_02776_ ), .B(_02780_ ), .Z(_04298_ ) );
INV_X1 _12046_ ( .A(_04298_ ), .ZN(_04299_ ) );
AOI211_X1 _12047_ ( .A(fanout_net_10 ), .B(_04297_ ), .C1(_04192_ ), .C2(_04299_ ), .ZN(_04300_ ) );
NAND3_X1 _12048_ ( .A1(_04292_ ), .A2(fanout_net_10 ), .A3(_04293_ ), .ZN(_04301_ ) );
INV_X1 _12049_ ( .A(_04301_ ), .ZN(_04302_ ) );
OAI21_X1 _12050_ ( .A(_04212_ ), .B1(_04300_ ), .B2(_04302_ ), .ZN(_04303_ ) );
OAI21_X1 _12051_ ( .A(fanout_net_8 ), .B1(_02604_ ), .B2(_02594_ ), .ZN(_04304_ ) );
AOI21_X1 _12052_ ( .A(_01653_ ), .B1(_04299_ ), .B2(_04227_ ), .ZN(_04305_ ) );
AOI21_X1 _12053_ ( .A(_04283_ ), .B1(_04304_ ), .B2(_04305_ ), .ZN(_04306_ ) );
AOI221_X1 _12054_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04295_ ), .C1(_04303_ ), .C2(_04306_ ), .ZN(_00126_ ) );
AND4_X1 _12055_ ( .A1(\mtvec [15] ), .A2(_02678_ ), .A3(_04204_ ), .A4(_02688_ ), .ZN(_04307_ ) );
NAND4_X1 _12056_ ( .A1(_04204_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_02688_ ), .A4(_04117_ ), .ZN(_04308_ ) );
NAND4_X1 _12057_ ( .A1(_04256_ ), .A2(_02697_ ), .A3(\mepc [15] ), .A4(_04174_ ), .ZN(_04309_ ) );
NAND4_X1 _12058_ ( .A1(_04172_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][15] ), .A4(_04134_ ), .ZN(_04310_ ) );
AND2_X1 _12059_ ( .A1(_04309_ ), .A2(_04310_ ), .ZN(_04311_ ) );
NAND3_X1 _12060_ ( .A1(_04168_ ), .A2(_04308_ ), .A3(_04311_ ), .ZN(_04312_ ) );
OAI21_X1 _12061_ ( .A(_02665_ ), .B1(_04307_ ), .B2(_04312_ ), .ZN(_04313_ ) );
NAND3_X1 _12062_ ( .A1(_02715_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_02717_ ), .ZN(_04314_ ) );
AND2_X1 _12063_ ( .A1(_04313_ ), .A2(_04314_ ), .ZN(_04315_ ) );
NAND3_X1 _12064_ ( .A1(_02847_ ), .A2(\ID_EX_pc [14] ), .A3(_04269_ ), .ZN(_04316_ ) );
XNOR2_X1 _12065_ ( .A(_04316_ ), .B(\ID_EX_pc [15] ), .ZN(_04317_ ) );
AOI21_X1 _12066_ ( .A(_04317_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04318_ ) );
INV_X1 _12067_ ( .A(_02763_ ), .ZN(_04319_ ) );
OAI21_X1 _12068_ ( .A(_02767_ ), .B1(_02752_ ), .B2(_02760_ ), .ZN(_04320_ ) );
AOI21_X1 _12069_ ( .A(_04319_ ), .B1(_04320_ ), .B2(_02773_ ), .ZN(_04321_ ) );
OR2_X1 _12070_ ( .A1(_04321_ ), .A2(_02769_ ), .ZN(_04322_ ) );
XNOR2_X1 _12071_ ( .A(_04322_ ), .B(_02762_ ), .ZN(_04323_ ) );
AOI211_X1 _12072_ ( .A(fanout_net_10 ), .B(_04318_ ), .C1(_04192_ ), .C2(_04323_ ), .ZN(_04324_ ) );
NAND2_X1 _12073_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [15] ), .ZN(_04325_ ) );
AOI21_X1 _12074_ ( .A(_04159_ ), .B1(_04313_ ), .B2(_04325_ ), .ZN(_04326_ ) );
OAI21_X1 _12075_ ( .A(_04212_ ), .B1(_04324_ ), .B2(_04326_ ), .ZN(_04327_ ) );
NAND2_X1 _12076_ ( .A1(_02611_ ), .A2(fanout_net_8 ), .ZN(_04328_ ) );
AOI21_X1 _12077_ ( .A(_01653_ ), .B1(_04323_ ), .B2(_04227_ ), .ZN(_04329_ ) );
AOI21_X1 _12078_ ( .A(_04283_ ), .B1(_04328_ ), .B2(_04329_ ), .ZN(_04330_ ) );
AOI221_X1 _12079_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04315_ ), .C1(_04327_ ), .C2(_04330_ ), .ZN(_00127_ ) );
AND4_X2 _12080_ ( .A1(_02642_ ), .A2(_02668_ ), .A3(_02670_ ), .A4(_02679_ ), .ZN(_04331_ ) );
AND3_X2 _12081_ ( .A1(_02666_ ), .A2(_02684_ ), .A3(_02672_ ), .ZN(_04332_ ) );
NAND3_X1 _12082_ ( .A1(_04331_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_04332_ ), .ZN(_04333_ ) );
NAND3_X1 _12083_ ( .A1(_04111_ ), .A2(\mepc [14] ), .A3(_04107_ ), .ZN(_04334_ ) );
NAND2_X1 _12084_ ( .A1(_04333_ ), .A2(_04334_ ), .ZN(_04335_ ) );
AOI21_X1 _12085_ ( .A(_04335_ ), .B1(_04181_ ), .B2(_04183_ ), .ZN(_04336_ ) );
AND4_X1 _12086_ ( .A1(\mycsreg.CSReg[3][14] ), .A2(_02697_ ), .A3(_04173_ ), .A4(_04134_ ), .ZN(_04337_ ) );
NOR3_X1 _12087_ ( .A1(_02675_ ), .A2(_04166_ ), .A3(_04337_ ), .ZN(_04338_ ) );
NAND4_X1 _12088_ ( .A1(_02668_ ), .A2(_02671_ ), .A3(_02679_ ), .A4(_02658_ ), .ZN(_04339_ ) );
NAND3_X1 _12089_ ( .A1(_02666_ ), .A2(_02684_ ), .A3(\ID_EX_csr [2] ), .ZN(_04340_ ) );
NOR2_X1 _12090_ ( .A1(_04339_ ), .A2(_04340_ ), .ZN(_04341_ ) );
NAND2_X1 _12091_ ( .A1(_04341_ ), .A2(\mtvec [14] ), .ZN(_04342_ ) );
NAND3_X1 _12092_ ( .A1(_04336_ ), .A2(_04338_ ), .A3(_04342_ ), .ZN(_04343_ ) );
OR3_X1 _12093_ ( .A1(_04262_ ), .A2(\EX_LS_result_csreg_mem [14] ), .A3(_04264_ ), .ZN(_04344_ ) );
AND2_X1 _12094_ ( .A1(_04343_ ), .A2(_04344_ ), .ZN(_04345_ ) );
INV_X1 _12095_ ( .A(_04345_ ), .ZN(_04346_ ) );
INV_X1 _12096_ ( .A(\ID_EX_pc [14] ), .ZN(_04347_ ) );
XNOR2_X1 _12097_ ( .A(_04270_ ), .B(_04347_ ), .ZN(_04348_ ) );
AOI21_X1 _12098_ ( .A(_04348_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04349_ ) );
NAND2_X1 _12099_ ( .A1(_04320_ ), .A2(_02773_ ), .ZN(_04350_ ) );
XNOR2_X1 _12100_ ( .A(_04350_ ), .B(_04319_ ), .ZN(_04351_ ) );
INV_X1 _12101_ ( .A(_04351_ ), .ZN(_04352_ ) );
AOI211_X1 _12102_ ( .A(fanout_net_10 ), .B(_04349_ ), .C1(_04192_ ), .C2(_04352_ ), .ZN(_04353_ ) );
AND3_X1 _12103_ ( .A1(_04343_ ), .A2(fanout_net_10 ), .A3(_04344_ ), .ZN(_04354_ ) );
OAI21_X1 _12104_ ( .A(_04212_ ), .B1(_04353_ ), .B2(_04354_ ), .ZN(_04355_ ) );
AOI21_X1 _12105_ ( .A(_02833_ ), .B1(_02612_ ), .B2(_02608_ ), .ZN(_04356_ ) );
OAI21_X1 _12106_ ( .A(_01649_ ), .B1(_04351_ ), .B2(fanout_net_8 ), .ZN(_04357_ ) );
NOR2_X1 _12107_ ( .A1(_04356_ ), .A2(_04357_ ), .ZN(_04358_ ) );
NOR2_X1 _12108_ ( .A1(_04358_ ), .A2(_04225_ ), .ZN(_04359_ ) );
AOI221_X1 _12109_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04346_ ), .C1(_04355_ ), .C2(_04359_ ), .ZN(_00128_ ) );
NAND4_X1 _12110_ ( .A1(_04203_ ), .A2(_02682_ ), .A3(\mtvec [13] ), .A4(_04107_ ), .ZN(_04360_ ) );
NAND4_X1 _12111_ ( .A1(_02682_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_04107_ ), .A4(_02703_ ), .ZN(_04361_ ) );
NAND4_X1 _12112_ ( .A1(_04256_ ), .A2(_02705_ ), .A3(\mepc [13] ), .A4(_02701_ ), .ZN(_04362_ ) );
NAND4_X1 _12113_ ( .A1(_02705_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][13] ), .A4(_02701_ ), .ZN(_04363_ ) );
NAND4_X1 _12114_ ( .A1(_04360_ ), .A2(_04361_ ), .A3(_04362_ ), .A4(_04363_ ), .ZN(_04364_ ) );
BUF_X2 _12115_ ( .A(_02652_ ), .Z(_04365_ ) );
BUF_X2 _12116_ ( .A(_02663_ ), .Z(_04366_ ) );
AOI211_X1 _12117_ ( .A(_02675_ ), .B(_04364_ ), .C1(_04365_ ), .C2(_04366_ ), .ZN(_04367_ ) );
INV_X1 _12118_ ( .A(\EX_LS_result_csreg_mem [13] ), .ZN(_04368_ ) );
AND3_X1 _12119_ ( .A1(_02714_ ), .A2(_04368_ ), .A3(_02716_ ), .ZN(_04369_ ) );
OR2_X1 _12120_ ( .A1(_04367_ ), .A2(_04369_ ), .ZN(_04370_ ) );
NAND3_X1 _12121_ ( .A1(_02846_ ), .A2(\ID_EX_pc [9] ), .A3(_04146_ ), .ZN(_04371_ ) );
INV_X1 _12122_ ( .A(\ID_EX_pc [12] ), .ZN(_04372_ ) );
NOR2_X1 _12123_ ( .A1(_04371_ ), .A2(_04372_ ), .ZN(_04373_ ) );
INV_X1 _12124_ ( .A(\ID_EX_pc [13] ), .ZN(_04374_ ) );
XNOR2_X1 _12125_ ( .A(_04373_ ), .B(_04374_ ), .ZN(_04375_ ) );
AOI21_X1 _12126_ ( .A(_04375_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04376_ ) );
OAI21_X1 _12127_ ( .A(_02766_ ), .B1(_02752_ ), .B2(_02760_ ), .ZN(_04377_ ) );
NAND2_X1 _12128_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_04378_ ) );
NAND2_X1 _12129_ ( .A1(_04377_ ), .A2(_04378_ ), .ZN(_04379_ ) );
XNOR2_X1 _12130_ ( .A(_04379_ ), .B(_02765_ ), .ZN(_04380_ ) );
AOI211_X1 _12131_ ( .A(fanout_net_10 ), .B(_04376_ ), .C1(_04192_ ), .C2(_04380_ ), .ZN(_04381_ ) );
OR3_X1 _12132_ ( .A1(_04120_ ), .A2(_04368_ ), .A3(_04121_ ), .ZN(_04382_ ) );
BUF_X4 _12133_ ( .A(_04140_ ), .Z(_04383_ ) );
BUF_X4 _12134_ ( .A(_02686_ ), .Z(_04384_ ) );
BUF_X4 _12135_ ( .A(_04384_ ), .Z(_04385_ ) );
NAND4_X1 _12136_ ( .A1(_04231_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][13] ), .A4(_04385_ ), .ZN(_04386_ ) );
AND2_X1 _12137_ ( .A1(_04105_ ), .A2(_04386_ ), .ZN(_04387_ ) );
BUF_X4 _12138_ ( .A(_04111_ ), .Z(_04388_ ) );
BUF_X4 _12139_ ( .A(_04384_ ), .Z(_04389_ ) );
BUF_X4 _12140_ ( .A(_04389_ ), .Z(_04390_ ) );
NAND3_X1 _12141_ ( .A1(_04388_ ), .A2(\mepc [13] ), .A3(_04390_ ), .ZN(_04391_ ) );
BUF_X4 _12142_ ( .A(_04203_ ), .Z(_04392_ ) );
BUF_X4 _12143_ ( .A(_02682_ ), .Z(_04393_ ) );
BUF_X4 _12144_ ( .A(_04112_ ), .Z(_04394_ ) );
NAND4_X1 _12145_ ( .A1(_04392_ ), .A2(_04393_ ), .A3(\mtvec [13] ), .A4(_04394_ ), .ZN(_04395_ ) );
BUF_X4 _12146_ ( .A(_02681_ ), .Z(_04396_ ) );
BUF_X4 _12147_ ( .A(_04396_ ), .Z(_04397_ ) );
BUF_X4 _12148_ ( .A(_02703_ ), .Z(_04398_ ) );
NAND4_X1 _12149_ ( .A1(_04397_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_04113_ ), .A4(_04398_ ), .ZN(_04399_ ) );
NAND4_X1 _12150_ ( .A1(_04387_ ), .A2(_04391_ ), .A3(_04395_ ), .A4(_04399_ ), .ZN(_04400_ ) );
BUF_X4 _12151_ ( .A(_04101_ ), .Z(_04401_ ) );
BUF_X4 _12152_ ( .A(_01677_ ), .Z(_04402_ ) );
OAI21_X1 _12153_ ( .A(_04400_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04403_ ) );
AOI21_X1 _12154_ ( .A(_04159_ ), .B1(_04382_ ), .B2(_04403_ ), .ZN(_04404_ ) );
OAI21_X1 _12155_ ( .A(_04212_ ), .B1(_04381_ ), .B2(_04404_ ), .ZN(_04405_ ) );
NAND2_X1 _12156_ ( .A1(_02615_ ), .A2(fanout_net_8 ), .ZN(_04406_ ) );
AOI21_X1 _12157_ ( .A(_01653_ ), .B1(_04380_ ), .B2(_02835_ ), .ZN(_04407_ ) );
AOI21_X1 _12158_ ( .A(_04283_ ), .B1(_04406_ ), .B2(_04407_ ), .ZN(_04408_ ) );
AOI221_X1 _12159_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04370_ ), .C1(_04405_ ), .C2(_04408_ ), .ZN(_00129_ ) );
NAND4_X1 _12160_ ( .A1(_04169_ ), .A2(_02682_ ), .A3(\mtvec [12] ), .A4(_02701_ ), .ZN(_04409_ ) );
NAND4_X1 _12161_ ( .A1(_04256_ ), .A2(_04172_ ), .A3(\mepc [12] ), .A4(_02709_ ), .ZN(_04410_ ) );
NAND4_X1 _12162_ ( .A1(_04233_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_02709_ ), .A4(_02703_ ), .ZN(_04411_ ) );
NAND4_X1 _12163_ ( .A1(_02705_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][12] ), .A4(_04170_ ), .ZN(_04412_ ) );
AND4_X1 _12164_ ( .A1(_04409_ ), .A2(_04410_ ), .A3(_04411_ ), .A4(_04412_ ), .ZN(_04413_ ) );
NAND3_X1 _12165_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04413_ ), .ZN(_04414_ ) );
INV_X1 _12166_ ( .A(\EX_LS_result_csreg_mem [12] ), .ZN(_04415_ ) );
NAND3_X1 _12167_ ( .A1(_04181_ ), .A2(_04415_ ), .A3(_04183_ ), .ZN(_04416_ ) );
AND2_X1 _12168_ ( .A1(_04414_ ), .A2(_04416_ ), .ZN(_04417_ ) );
INV_X1 _12169_ ( .A(_04417_ ), .ZN(_04418_ ) );
XNOR2_X1 _12170_ ( .A(_04371_ ), .B(\ID_EX_pc [12] ), .ZN(_04419_ ) );
AOI21_X1 _12171_ ( .A(_04419_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04420_ ) );
XOR2_X1 _12172_ ( .A(_02761_ ), .B(_02766_ ), .Z(_04421_ ) );
INV_X1 _12173_ ( .A(_04421_ ), .ZN(_04422_ ) );
AOI211_X1 _12174_ ( .A(fanout_net_10 ), .B(_04420_ ), .C1(_04192_ ), .C2(_04422_ ), .ZN(_04423_ ) );
AND3_X1 _12175_ ( .A1(_04414_ ), .A2(fanout_net_10 ), .A3(_04416_ ), .ZN(_04424_ ) );
OAI21_X1 _12176_ ( .A(_04212_ ), .B1(_04423_ ), .B2(_04424_ ), .ZN(_04425_ ) );
AOI21_X1 _12177_ ( .A(_02720_ ), .B1(_04422_ ), .B2(_02833_ ), .ZN(_04426_ ) );
BUF_X4 _12178_ ( .A(_02832_ ), .Z(_04427_ ) );
OAI21_X1 _12179_ ( .A(_04426_ ), .B1(_02616_ ), .B2(_04427_ ), .ZN(_04428_ ) );
AND2_X1 _12180_ ( .A1(_04428_ ), .A2(_02838_ ), .ZN(_04429_ ) );
AOI221_X1 _12181_ ( .A(fanout_net_2 ), .B1(_02638_ ), .B2(_04418_ ), .C1(_04425_ ), .C2(_04429_ ), .ZN(_00130_ ) );
BUF_X4 _12182_ ( .A(_02578_ ), .Z(_04430_ ) );
NAND4_X1 _12183_ ( .A1(_04169_ ), .A2(_04133_ ), .A3(\mtvec [11] ), .A4(_04170_ ), .ZN(_04431_ ) );
NAND4_X1 _12184_ ( .A1(_04256_ ), .A2(_02697_ ), .A3(\mepc [11] ), .A4(_04174_ ), .ZN(_04432_ ) );
NAND4_X1 _12185_ ( .A1(_04133_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_04134_ ), .A4(_04136_ ), .ZN(_04433_ ) );
NAND4_X1 _12186_ ( .A1(_02697_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][11] ), .A4(_04134_ ), .ZN(_04434_ ) );
AND4_X1 _12187_ ( .A1(_04431_ ), .A2(_04432_ ), .A3(_04433_ ), .A4(_04434_ ), .ZN(_04435_ ) );
NAND3_X1 _12188_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04435_ ), .ZN(_04436_ ) );
INV_X1 _12189_ ( .A(\EX_LS_result_csreg_mem [11] ), .ZN(_04437_ ) );
NAND3_X1 _12190_ ( .A1(_04181_ ), .A2(_04437_ ), .A3(_04183_ ), .ZN(_04438_ ) );
AND2_X1 _12191_ ( .A1(_04436_ ), .A2(_04438_ ), .ZN(_04439_ ) );
INV_X1 _12192_ ( .A(_04439_ ), .ZN(_04440_ ) );
AND2_X1 _12193_ ( .A1(_02847_ ), .A2(\ID_EX_pc [10] ), .ZN(_04441_ ) );
INV_X1 _12194_ ( .A(\ID_EX_pc [11] ), .ZN(_04442_ ) );
XNOR2_X1 _12195_ ( .A(_04441_ ), .B(_04442_ ), .ZN(_04443_ ) );
AOI21_X1 _12196_ ( .A(_04443_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04444_ ) );
INV_X1 _12197_ ( .A(_02747_ ), .ZN(_04445_ ) );
OAI21_X1 _12198_ ( .A(_02751_ ), .B1(_02743_ ), .B2(_02744_ ), .ZN(_04446_ ) );
AOI21_X1 _12199_ ( .A(_04445_ ), .B1(_04446_ ), .B2(_02758_ ), .ZN(_04447_ ) );
OR2_X1 _12200_ ( .A1(_04447_ ), .A2(_02753_ ), .ZN(_04448_ ) );
XNOR2_X1 _12201_ ( .A(_04448_ ), .B(_02746_ ), .ZN(_04449_ ) );
AOI211_X1 _12202_ ( .A(fanout_net_10 ), .B(_04444_ ), .C1(_04192_ ), .C2(_04449_ ), .ZN(_04450_ ) );
AND3_X1 _12203_ ( .A1(_04436_ ), .A2(fanout_net_10 ), .A3(_04438_ ), .ZN(_04451_ ) );
OAI21_X1 _12204_ ( .A(_04212_ ), .B1(_04450_ ), .B2(_04451_ ), .ZN(_04452_ ) );
AOI21_X1 _12205_ ( .A(_02720_ ), .B1(_04449_ ), .B2(_02833_ ), .ZN(_04453_ ) );
OAI21_X1 _12206_ ( .A(_02228_ ), .B1(_02174_ ), .B2(_02180_ ), .ZN(_04454_ ) );
AOI21_X1 _12207_ ( .A(_02284_ ), .B1(\ID_EX_imm [9] ), .B2(_02225_ ), .ZN(_04455_ ) );
AND2_X1 _12208_ ( .A1(_04454_ ), .A2(_04455_ ), .ZN(_04456_ ) );
AND3_X1 _12209_ ( .A1(_02247_ ), .A2(_02250_ ), .A3(_02248_ ), .ZN(_04457_ ) );
NOR3_X1 _12210_ ( .A1(_04456_ ), .A2(_02279_ ), .A3(_04457_ ), .ZN(_04458_ ) );
NOR2_X1 _12211_ ( .A1(_04458_ ), .A2(_02279_ ), .ZN(_04459_ ) );
XNOR2_X1 _12212_ ( .A(_04459_ ), .B(_02274_ ), .ZN(_04460_ ) );
OAI21_X1 _12213_ ( .A(_04453_ ), .B1(_04460_ ), .B2(_04427_ ), .ZN(_04461_ ) );
AND2_X1 _12214_ ( .A1(_04461_ ), .A2(_02838_ ), .ZN(_04462_ ) );
AOI221_X1 _12215_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04440_ ), .C1(_04452_ ), .C2(_04462_ ), .ZN(_00131_ ) );
NAND4_X1 _12216_ ( .A1(_04203_ ), .A2(_02682_ ), .A3(\mtvec [28] ), .A4(_04107_ ), .ZN(_04463_ ) );
NAND4_X1 _12217_ ( .A1(_02682_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_04107_ ), .A4(_02703_ ), .ZN(_04464_ ) );
NAND4_X1 _12218_ ( .A1(_04256_ ), .A2(_02705_ ), .A3(\mepc [28] ), .A4(_02701_ ), .ZN(_04465_ ) );
NAND4_X1 _12219_ ( .A1(_02705_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][28] ), .A4(_02701_ ), .ZN(_04466_ ) );
NAND4_X1 _12220_ ( .A1(_04463_ ), .A2(_04464_ ), .A3(_04465_ ), .A4(_04466_ ), .ZN(_04467_ ) );
AOI211_X1 _12221_ ( .A(_02675_ ), .B(_04467_ ), .C1(_04365_ ), .C2(_02716_ ), .ZN(_04468_ ) );
INV_X1 _12222_ ( .A(\EX_LS_result_csreg_mem [28] ), .ZN(_04469_ ) );
AND3_X1 _12223_ ( .A1(_02714_ ), .A2(_04469_ ), .A3(_02716_ ), .ZN(_04470_ ) );
OR2_X1 _12224_ ( .A1(_04468_ ), .A2(_04470_ ), .ZN(_04471_ ) );
INV_X1 _12225_ ( .A(\ID_EX_pc [28] ), .ZN(_04472_ ) );
XNOR2_X1 _12226_ ( .A(_04155_ ), .B(_04472_ ), .ZN(_04473_ ) );
AOI21_X1 _12227_ ( .A(_04473_ ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_04474_ ) );
BUF_X4 _12228_ ( .A(_04084_ ), .Z(_04475_ ) );
XNOR2_X1 _12229_ ( .A(_02821_ ), .B(_02822_ ), .ZN(_04476_ ) );
AOI211_X1 _12230_ ( .A(fanout_net_10 ), .B(_04474_ ), .C1(_04475_ ), .C2(_04476_ ), .ZN(_04477_ ) );
OR3_X1 _12231_ ( .A1(_04120_ ), .A2(_04469_ ), .A3(_04121_ ), .ZN(_04478_ ) );
NAND4_X1 _12232_ ( .A1(_04231_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][28] ), .A4(_04385_ ), .ZN(_04479_ ) );
AND2_X1 _12233_ ( .A1(_04105_ ), .A2(_04479_ ), .ZN(_04480_ ) );
NAND3_X1 _12234_ ( .A1(_04388_ ), .A2(\mepc [28] ), .A3(_04390_ ), .ZN(_04481_ ) );
NAND4_X1 _12235_ ( .A1(_04392_ ), .A2(_02683_ ), .A3(\mtvec [28] ), .A4(_04394_ ), .ZN(_04482_ ) );
NAND4_X1 _12236_ ( .A1(_04397_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_04113_ ), .A4(_04398_ ), .ZN(_04483_ ) );
NAND4_X1 _12237_ ( .A1(_04480_ ), .A2(_04481_ ), .A3(_04482_ ), .A4(_04483_ ), .ZN(_04484_ ) );
OAI21_X1 _12238_ ( .A(_04484_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04485_ ) );
AOI21_X1 _12239_ ( .A(_04159_ ), .B1(_04478_ ), .B2(_04485_ ), .ZN(_04486_ ) );
OAI21_X1 _12240_ ( .A(_04212_ ), .B1(_04477_ ), .B2(_04486_ ), .ZN(_04487_ ) );
OAI21_X1 _12241_ ( .A(fanout_net_8 ), .B1(_02619_ ), .B2(_02517_ ), .ZN(_04488_ ) );
AOI21_X1 _12242_ ( .A(_01653_ ), .B1(_04476_ ), .B2(_02835_ ), .ZN(_04489_ ) );
AOI21_X1 _12243_ ( .A(_04283_ ), .B1(_04488_ ), .B2(_04489_ ), .ZN(_04490_ ) );
AOI221_X1 _12244_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04471_ ), .C1(_04487_ ), .C2(_04490_ ), .ZN(_00132_ ) );
NAND4_X1 _12245_ ( .A1(_04231_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][10] ), .A4(_04389_ ), .ZN(_04491_ ) );
NAND3_X1 _12246_ ( .A1(_04111_ ), .A2(\mepc [10] ), .A3(_04205_ ), .ZN(_04492_ ) );
NAND4_X1 _12247_ ( .A1(_04203_ ), .A2(_04396_ ), .A3(\mtvec [10] ), .A4(_04385_ ), .ZN(_04493_ ) );
NAND4_X1 _12248_ ( .A1(_04167_ ), .A2(_04491_ ), .A3(_04492_ ), .A4(_04493_ ), .ZN(_04494_ ) );
AND4_X1 _12249_ ( .A1(\mycsreg.CSReg[0][10] ), .A2(_04204_ ), .A3(_04205_ ), .A4(_04117_ ), .ZN(_04495_ ) );
OAI21_X1 _12250_ ( .A(_02665_ ), .B1(_04494_ ), .B2(_04495_ ), .ZN(_04496_ ) );
NAND3_X1 _12251_ ( .A1(_04365_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_04366_ ), .ZN(_04497_ ) );
AND2_X1 _12252_ ( .A1(_04496_ ), .A2(_04497_ ), .ZN(_04498_ ) );
BUF_X4 _12253_ ( .A(_01653_ ), .Z(_04499_ ) );
INV_X1 _12254_ ( .A(\ID_EX_pc [10] ), .ZN(_04500_ ) );
XNOR2_X1 _12255_ ( .A(_02847_ ), .B(_04500_ ), .ZN(_04501_ ) );
BUF_X4 _12256_ ( .A(_04078_ ), .Z(_04502_ ) );
BUF_X4 _12257_ ( .A(_04081_ ), .Z(_04503_ ) );
AOI21_X1 _12258_ ( .A(_04501_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04504_ ) );
NAND2_X1 _12259_ ( .A1(_04446_ ), .A2(_02758_ ), .ZN(_04505_ ) );
XNOR2_X1 _12260_ ( .A(_04505_ ), .B(_04445_ ), .ZN(_04506_ ) );
INV_X1 _12261_ ( .A(_04506_ ), .ZN(_04507_ ) );
AOI211_X1 _12262_ ( .A(fanout_net_10 ), .B(_04504_ ), .C1(_04475_ ), .C2(_04507_ ), .ZN(_04508_ ) );
NAND2_X1 _12263_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [10] ), .ZN(_04509_ ) );
AOI21_X1 _12264_ ( .A(_04159_ ), .B1(_04496_ ), .B2(_04509_ ), .ZN(_04510_ ) );
OAI21_X1 _12265_ ( .A(_04499_ ), .B1(_04508_ ), .B2(_04510_ ), .ZN(_04511_ ) );
BUF_X4 _12266_ ( .A(_02832_ ), .Z(_04512_ ) );
AOI21_X1 _12267_ ( .A(_02720_ ), .B1(_04507_ ), .B2(_04512_ ), .ZN(_04513_ ) );
XNOR2_X1 _12268_ ( .A(_04456_ ), .B(_02251_ ), .ZN(_04514_ ) );
OAI21_X1 _12269_ ( .A(_04513_ ), .B1(_04514_ ), .B2(_04427_ ), .ZN(_04515_ ) );
CLKBUF_X2 _12270_ ( .A(_02837_ ), .Z(_04516_ ) );
AND2_X1 _12271_ ( .A1(_04515_ ), .A2(_04516_ ), .ZN(_04517_ ) );
AOI221_X1 _12272_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04498_ ), .C1(_04511_ ), .C2(_04517_ ), .ZN(_00133_ ) );
AND4_X1 _12273_ ( .A1(\mtvec [9] ), .A2(_02677_ ), .A3(_02681_ ), .A4(_04384_ ), .ZN(_04518_ ) );
NAND4_X1 _12274_ ( .A1(_02690_ ), .A2(_02696_ ), .A3(\mepc [9] ), .A4(_02700_ ), .ZN(_04519_ ) );
NAND4_X1 _12275_ ( .A1(_02680_ ), .A2(\mycsreg.CSReg[0][9] ), .A3(_02686_ ), .A4(_02702_ ), .ZN(_04520_ ) );
NAND4_X1 _12276_ ( .A1(_02695_ ), .A2(_02707_ ), .A3(\mycsreg.CSReg[3][9] ), .A4(_02686_ ), .ZN(_04521_ ) );
AND2_X1 _12277_ ( .A1(_04520_ ), .A2(_04521_ ), .ZN(_04522_ ) );
NAND3_X1 _12278_ ( .A1(_04167_ ), .A2(_04519_ ), .A3(_04522_ ), .ZN(_04523_ ) );
OAI21_X1 _12279_ ( .A(_02665_ ), .B1(_04518_ ), .B2(_04523_ ), .ZN(_04524_ ) );
NAND3_X1 _12280_ ( .A1(_02652_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_02663_ ), .ZN(_04525_ ) );
AND2_X1 _12281_ ( .A1(_04524_ ), .A2(_04525_ ), .ZN(_04526_ ) );
OR2_X1 _12282_ ( .A1(_04526_ ), .A2(_04086_ ), .ZN(_04527_ ) );
XNOR2_X1 _12283_ ( .A(_02846_ ), .B(\ID_EX_pc [9] ), .ZN(_04528_ ) );
AND2_X1 _12284_ ( .A1(_02745_ ), .A2(_02749_ ), .ZN(_04529_ ) );
OR2_X1 _12285_ ( .A1(_04529_ ), .A2(_02756_ ), .ZN(_04530_ ) );
XNOR2_X1 _12286_ ( .A(_04530_ ), .B(_02750_ ), .ZN(_04531_ ) );
MUX2_X1 _12287_ ( .A(_04528_ ), .B(_04531_ ), .S(_04084_ ), .Z(_04532_ ) );
OAI21_X1 _12288_ ( .A(_04527_ ), .B1(_04532_ ), .B2(fanout_net_10 ), .ZN(_04533_ ) );
NAND2_X1 _12289_ ( .A1(_04533_ ), .A2(_01654_ ), .ZN(_04534_ ) );
AND3_X1 _12290_ ( .A1(_02200_ ), .A2(_02203_ ), .A3(_02201_ ), .ZN(_04535_ ) );
NOR3_X1 _12291_ ( .A1(_02181_ ), .A2(_02283_ ), .A3(_04535_ ), .ZN(_04536_ ) );
OR2_X1 _12292_ ( .A1(_04536_ ), .A2(_02283_ ), .ZN(_04537_ ) );
XNOR2_X1 _12293_ ( .A(_04537_ ), .B(_02227_ ), .ZN(_04538_ ) );
NAND2_X1 _12294_ ( .A1(_04538_ ), .A2(fanout_net_8 ), .ZN(_04539_ ) );
AOI21_X1 _12295_ ( .A(_01653_ ), .B1(_04531_ ), .B2(_02835_ ), .ZN(_04540_ ) );
AOI21_X1 _12296_ ( .A(_04283_ ), .B1(_04539_ ), .B2(_04540_ ), .ZN(_04541_ ) );
AOI221_X1 _12297_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04526_ ), .C1(_04534_ ), .C2(_04541_ ), .ZN(_00134_ ) );
AND3_X1 _12298_ ( .A1(_04331_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_04332_ ), .ZN(_04542_ ) );
AOI21_X1 _12299_ ( .A(_04542_ ), .B1(_04181_ ), .B2(_04183_ ), .ZN(_04543_ ) );
AND3_X1 _12300_ ( .A1(_04110_ ), .A2(\mepc [8] ), .A3(_04384_ ), .ZN(_04544_ ) );
AND4_X1 _12301_ ( .A1(\mycsreg.CSReg[3][8] ), .A2(_02696_ ), .A3(_04140_ ), .A4(_02700_ ), .ZN(_04545_ ) );
NOR4_X1 _12302_ ( .A1(_02675_ ), .A2(_04166_ ), .A3(_04544_ ), .A4(_04545_ ), .ZN(_04546_ ) );
NAND4_X1 _12303_ ( .A1(_02678_ ), .A2(_02683_ ), .A3(\mtvec [8] ), .A4(_04115_ ), .ZN(_04547_ ) );
NAND3_X1 _12304_ ( .A1(_04543_ ), .A2(_04546_ ), .A3(_04547_ ), .ZN(_04548_ ) );
INV_X1 _12305_ ( .A(\EX_LS_result_csreg_mem [8] ), .ZN(_04549_ ) );
NAND3_X1 _12306_ ( .A1(_04181_ ), .A2(_04549_ ), .A3(_04183_ ), .ZN(_04550_ ) );
AND2_X1 _12307_ ( .A1(_04548_ ), .A2(_04550_ ), .ZN(_04551_ ) );
INV_X1 _12308_ ( .A(_04551_ ), .ZN(_04552_ ) );
INV_X1 _12309_ ( .A(\ID_EX_pc [8] ), .ZN(_04553_ ) );
XNOR2_X1 _12310_ ( .A(_02845_ ), .B(_04553_ ), .ZN(_04554_ ) );
AOI21_X1 _12311_ ( .A(_04554_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04555_ ) );
XOR2_X1 _12312_ ( .A(_02745_ ), .B(_02749_ ), .Z(_04556_ ) );
INV_X1 _12313_ ( .A(_04556_ ), .ZN(_04557_ ) );
AOI211_X1 _12314_ ( .A(fanout_net_10 ), .B(_04555_ ), .C1(_04475_ ), .C2(_04557_ ), .ZN(_04558_ ) );
AND3_X1 _12315_ ( .A1(_04548_ ), .A2(fanout_net_10 ), .A3(_04550_ ), .ZN(_04559_ ) );
OAI21_X1 _12316_ ( .A(_04499_ ), .B1(_04558_ ), .B2(_04559_ ), .ZN(_04560_ ) );
BUF_X4 _12317_ ( .A(_01652_ ), .Z(_04561_ ) );
AOI21_X1 _12318_ ( .A(_04561_ ), .B1(_04557_ ), .B2(_04512_ ), .ZN(_04562_ ) );
XNOR2_X1 _12319_ ( .A(_02181_ ), .B(_02204_ ), .ZN(_04563_ ) );
OAI21_X1 _12320_ ( .A(_04562_ ), .B1(_04563_ ), .B2(_04427_ ), .ZN(_04564_ ) );
AND2_X1 _12321_ ( .A1(_04564_ ), .A2(_04516_ ), .ZN(_04565_ ) );
AOI221_X1 _12322_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04552_ ), .C1(_04560_ ), .C2(_04565_ ), .ZN(_00135_ ) );
AND3_X1 _12323_ ( .A1(_04365_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_04366_ ), .ZN(_04566_ ) );
NAND4_X1 _12324_ ( .A1(_02691_ ), .A2(_04231_ ), .A3(\mepc [7] ), .A4(_04389_ ), .ZN(_04567_ ) );
NAND4_X1 _12325_ ( .A1(_04204_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_04389_ ), .A4(_04117_ ), .ZN(_04568_ ) );
NAND4_X1 _12326_ ( .A1(_04231_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][7] ), .A4(_04389_ ), .ZN(_04569_ ) );
AND3_X1 _12327_ ( .A1(_04567_ ), .A2(_04568_ ), .A3(_04569_ ), .ZN(_04570_ ) );
BUF_X4 _12328_ ( .A(_04205_ ), .Z(_04571_ ) );
NAND4_X1 _12329_ ( .A1(_04392_ ), .A2(_04397_ ), .A3(\mtvec [7] ), .A4(_04571_ ), .ZN(_04572_ ) );
AOI22_X1 _12330_ ( .A1(_02715_ ), .A2(_02717_ ), .B1(_04570_ ), .B2(_04572_ ), .ZN(_04573_ ) );
NOR2_X1 _12331_ ( .A1(_04566_ ), .A2(_04573_ ), .ZN(_04574_ ) );
INV_X1 _12332_ ( .A(\ID_EX_pc [7] ), .ZN(_04575_ ) );
XNOR2_X1 _12333_ ( .A(_02844_ ), .B(_04575_ ), .ZN(_04576_ ) );
AOI21_X1 _12334_ ( .A(_04576_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04577_ ) );
NAND2_X1 _12335_ ( .A1(_02741_ ), .A2(_02742_ ), .ZN(_04578_ ) );
NOR2_X1 _12336_ ( .A1(_02744_ ), .A2(_02721_ ), .ZN(_04579_ ) );
XNOR2_X1 _12337_ ( .A(_04578_ ), .B(_04579_ ), .ZN(_04580_ ) );
AOI211_X1 _12338_ ( .A(fanout_net_10 ), .B(_04577_ ), .C1(_04475_ ), .C2(_04580_ ), .ZN(_04581_ ) );
INV_X1 _12339_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_04582_ ) );
OR3_X1 _12340_ ( .A1(_04120_ ), .A2(_04582_ ), .A3(_04121_ ), .ZN(_04583_ ) );
NAND3_X1 _12341_ ( .A1(_04388_ ), .A2(\mepc [7] ), .A3(_04390_ ), .ZN(_04584_ ) );
NAND4_X1 _12342_ ( .A1(_04392_ ), .A2(_04393_ ), .A3(\mtvec [7] ), .A4(_04113_ ), .ZN(_04585_ ) );
NAND4_X1 _12343_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][7] ), .A4(_04394_ ), .ZN(_04586_ ) );
NAND4_X1 _12344_ ( .A1(_04397_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_04113_ ), .A4(_04398_ ), .ZN(_04587_ ) );
NAND4_X1 _12345_ ( .A1(_04584_ ), .A2(_04585_ ), .A3(_04586_ ), .A4(_04587_ ), .ZN(_04588_ ) );
OAI21_X1 _12346_ ( .A(_04588_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04589_ ) );
AOI21_X1 _12347_ ( .A(_04159_ ), .B1(_04583_ ), .B2(_04589_ ), .ZN(_04590_ ) );
OAI21_X1 _12348_ ( .A(_04499_ ), .B1(_04581_ ), .B2(_04590_ ), .ZN(_04591_ ) );
OAI21_X1 _12349_ ( .A(_02172_ ), .B1(_02122_ ), .B2(_02127_ ), .ZN(_04592_ ) );
AND2_X1 _12350_ ( .A1(_04592_ ), .A2(_02176_ ), .ZN(_04593_ ) );
XNOR2_X1 _12351_ ( .A(_04593_ ), .B(_02150_ ), .ZN(_04594_ ) );
NAND2_X1 _12352_ ( .A1(_04594_ ), .A2(fanout_net_8 ), .ZN(_04595_ ) );
AOI21_X1 _12353_ ( .A(_02720_ ), .B1(_04580_ ), .B2(_02835_ ), .ZN(_04596_ ) );
AOI21_X1 _12354_ ( .A(_04283_ ), .B1(_04595_ ), .B2(_04596_ ), .ZN(_04597_ ) );
AOI221_X1 _12355_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04574_ ), .C1(_04591_ ), .C2(_04597_ ), .ZN(_00136_ ) );
NAND4_X1 _12356_ ( .A1(_04203_ ), .A2(_04396_ ), .A3(\mtvec [6] ), .A4(_04385_ ), .ZN(_04598_ ) );
NAND4_X1 _12357_ ( .A1(_02691_ ), .A2(_04106_ ), .A3(\mepc [6] ), .A4(_04112_ ), .ZN(_04599_ ) );
NAND4_X1 _12358_ ( .A1(_04396_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_04112_ ), .A4(_02703_ ), .ZN(_04600_ ) );
NAND4_X1 _12359_ ( .A1(_04106_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][6] ), .A4(_04112_ ), .ZN(_04601_ ) );
NAND4_X1 _12360_ ( .A1(_04598_ ), .A2(_04599_ ), .A3(_04600_ ), .A4(_04601_ ), .ZN(_04602_ ) );
AOI211_X1 _12361_ ( .A(_02675_ ), .B(_04602_ ), .C1(_04365_ ), .C2(_04366_ ), .ZN(_04603_ ) );
INV_X1 _12362_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_04604_ ) );
AND3_X1 _12363_ ( .A1(_02714_ ), .A2(_04604_ ), .A3(_04366_ ), .ZN(_04605_ ) );
NOR2_X1 _12364_ ( .A1(_04603_ ), .A2(_04605_ ), .ZN(_04606_ ) );
INV_X1 _12365_ ( .A(_04606_ ), .ZN(_04607_ ) );
NAND3_X1 _12366_ ( .A1(_04181_ ), .A2(_04604_ ), .A3(_04183_ ), .ZN(_04608_ ) );
NAND3_X1 _12367_ ( .A1(_04331_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_04332_ ), .ZN(_04609_ ) );
OAI21_X1 _12368_ ( .A(_04609_ ), .B1(_04261_ ), .B2(_04263_ ), .ZN(_04610_ ) );
AND4_X1 _12369_ ( .A1(\mycsreg.CSReg[3][6] ), .A2(_02696_ ), .A3(_04140_ ), .A4(_02686_ ), .ZN(_04611_ ) );
AOI21_X1 _12370_ ( .A(_04611_ ), .B1(_02691_ ), .B2(_02669_ ), .ZN(_04612_ ) );
NAND3_X1 _12371_ ( .A1(_04111_ ), .A2(\mepc [6] ), .A3(_04389_ ), .ZN(_04613_ ) );
NAND2_X1 _12372_ ( .A1(_04341_ ), .A2(\mtvec [6] ), .ZN(_04614_ ) );
NAND3_X1 _12373_ ( .A1(_04612_ ), .A2(_04613_ ), .A3(_04614_ ), .ZN(_04615_ ) );
OAI211_X1 _12374_ ( .A(_04608_ ), .B(fanout_net_10 ), .C1(_04610_ ), .C2(_04615_ ), .ZN(_04616_ ) );
INV_X1 _12375_ ( .A(_04616_ ), .ZN(_04617_ ) );
INV_X1 _12376_ ( .A(\ID_EX_pc [6] ), .ZN(_04618_ ) );
XNOR2_X1 _12377_ ( .A(_02843_ ), .B(_04618_ ), .ZN(_04619_ ) );
OR2_X1 _12378_ ( .A1(_02739_ ), .A2(_02740_ ), .ZN(_04620_ ) );
XOR2_X1 _12379_ ( .A(_04620_ ), .B(_02722_ ), .Z(_04621_ ) );
MUX2_X1 _12380_ ( .A(_04619_ ), .B(_04621_ ), .S(_04083_ ), .Z(_04622_ ) );
AOI21_X1 _12381_ ( .A(_04617_ ), .B1(_04622_ ), .B2(_04086_ ), .ZN(_04623_ ) );
OR2_X2 _12382_ ( .A1(_04623_ ), .A2(_01649_ ), .ZN(_04624_ ) );
XNOR2_X1 _12383_ ( .A(_02128_ ), .B(_02172_ ), .ZN(_04625_ ) );
MUX2_X1 _12384_ ( .A(_04621_ ), .B(_04625_ ), .S(fanout_net_8 ), .Z(_04626_ ) );
AOI21_X1 _12385_ ( .A(_04283_ ), .B1(_04626_ ), .B2(_01649_ ), .ZN(_04627_ ) );
AOI221_X1 _12386_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04607_ ), .C1(_04624_ ), .C2(_04627_ ), .ZN(_00137_ ) );
NAND4_X1 _12387_ ( .A1(_04203_ ), .A2(_04396_ ), .A3(\mtvec [5] ), .A4(_04112_ ), .ZN(_04628_ ) );
NAND4_X1 _12388_ ( .A1(_04396_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_04112_ ), .A4(_02703_ ), .ZN(_04629_ ) );
NAND4_X1 _12389_ ( .A1(_02691_ ), .A2(_02705_ ), .A3(\mepc [5] ), .A4(_04107_ ), .ZN(_04630_ ) );
NAND4_X1 _12390_ ( .A1(_02705_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][5] ), .A4(_04107_ ), .ZN(_04631_ ) );
NAND4_X1 _12391_ ( .A1(_04628_ ), .A2(_04629_ ), .A3(_04630_ ), .A4(_04631_ ), .ZN(_04632_ ) );
AOI211_X1 _12392_ ( .A(_02675_ ), .B(_04632_ ), .C1(_04365_ ), .C2(_04366_ ), .ZN(_04633_ ) );
INV_X1 _12393_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_04634_ ) );
AND3_X1 _12394_ ( .A1(_02714_ ), .A2(_04634_ ), .A3(_02716_ ), .ZN(_04635_ ) );
NOR2_X1 _12395_ ( .A1(_04633_ ), .A2(_04635_ ), .ZN(_04636_ ) );
INV_X1 _12396_ ( .A(_04636_ ), .ZN(_04637_ ) );
XNOR2_X1 _12397_ ( .A(_02842_ ), .B(\ID_EX_pc [5] ), .ZN(_04638_ ) );
AND2_X2 _12398_ ( .A1(_04268_ ), .A2(_04638_ ), .ZN(_04639_ ) );
NAND2_X1 _12399_ ( .A1(_02737_ ), .A2(_02738_ ), .ZN(_04640_ ) );
NOR2_X1 _12400_ ( .A1(_02740_ ), .A2(_02723_ ), .ZN(_04641_ ) );
XNOR2_X1 _12401_ ( .A(_04640_ ), .B(_04641_ ), .ZN(_04642_ ) );
AOI211_X2 _12402_ ( .A(fanout_net_10 ), .B(_04639_ ), .C1(_04475_ ), .C2(_04642_ ), .ZN(_04643_ ) );
BUF_X4 _12403_ ( .A(_04086_ ), .Z(_04644_ ) );
OR3_X1 _12404_ ( .A1(_04120_ ), .A2(_04634_ ), .A3(_04121_ ), .ZN(_04645_ ) );
NAND4_X1 _12405_ ( .A1(_04106_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][5] ), .A4(_04385_ ), .ZN(_04646_ ) );
AND2_X1 _12406_ ( .A1(_04105_ ), .A2(_04646_ ), .ZN(_04647_ ) );
NAND3_X1 _12407_ ( .A1(_04388_ ), .A2(\mepc [5] ), .A3(_04390_ ), .ZN(_04648_ ) );
NAND4_X1 _12408_ ( .A1(_04392_ ), .A2(_02683_ ), .A3(\mtvec [5] ), .A4(_04394_ ), .ZN(_04649_ ) );
NAND4_X1 _12409_ ( .A1(_04397_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_04113_ ), .A4(_04398_ ), .ZN(_04650_ ) );
NAND4_X1 _12410_ ( .A1(_04647_ ), .A2(_04648_ ), .A3(_04649_ ), .A4(_04650_ ), .ZN(_04651_ ) );
OAI21_X1 _12411_ ( .A(_04651_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04652_ ) );
AOI21_X1 _12412_ ( .A(_04644_ ), .B1(_04645_ ), .B2(_04652_ ), .ZN(_04653_ ) );
OAI21_X1 _12413_ ( .A(_04499_ ), .B1(_04643_ ), .B2(_04653_ ), .ZN(_04654_ ) );
NOR2_X1 _12414_ ( .A1(_02073_ ), .A2(_02121_ ), .ZN(_04655_ ) );
AND2_X1 _12415_ ( .A1(_02118_ ), .A2(\ID_EX_imm [4] ), .ZN(_04656_ ) );
NOR2_X1 _12416_ ( .A1(_04655_ ), .A2(_04656_ ), .ZN(_04657_ ) );
XNOR2_X1 _12417_ ( .A(_04657_ ), .B(_02097_ ), .ZN(_04658_ ) );
NAND2_X1 _12418_ ( .A1(_04658_ ), .A2(fanout_net_8 ), .ZN(_04659_ ) );
AOI21_X1 _12419_ ( .A(_02720_ ), .B1(_04642_ ), .B2(_02835_ ), .ZN(_04660_ ) );
AOI21_X1 _12420_ ( .A(_04283_ ), .B1(_04659_ ), .B2(_04660_ ), .ZN(_04661_ ) );
AOI221_X1 _12421_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04637_ ), .C1(_04654_ ), .C2(_04661_ ), .ZN(_00138_ ) );
NAND4_X1 _12422_ ( .A1(_02677_ ), .A2(_02681_ ), .A3(\mtvec [4] ), .A4(_02687_ ), .ZN(_04662_ ) );
NAND4_X1 _12423_ ( .A1(_04138_ ), .A2(_04140_ ), .A3(\mycsreg.CSReg[3][4] ), .A4(_04384_ ), .ZN(_04663_ ) );
NAND4_X1 _12424_ ( .A1(_02681_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_04384_ ), .A4(_04136_ ), .ZN(_04664_ ) );
NAND4_X1 _12425_ ( .A1(_02690_ ), .A2(_04138_ ), .A3(\mepc [4] ), .A4(_04384_ ), .ZN(_04665_ ) );
NAND4_X1 _12426_ ( .A1(_04662_ ), .A2(_04663_ ), .A3(_04664_ ), .A4(_04665_ ), .ZN(_04666_ ) );
AOI211_X1 _12427_ ( .A(_02674_ ), .B(_04666_ ), .C1(_02652_ ), .C2(_02663_ ), .ZN(_04667_ ) );
INV_X1 _12428_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_04668_ ) );
AND3_X1 _12429_ ( .A1(_02652_ ), .A2(_04668_ ), .A3(_02663_ ), .ZN(_04669_ ) );
NOR2_X1 _12430_ ( .A1(_04667_ ), .A2(_04669_ ), .ZN(_04670_ ) );
INV_X1 _12431_ ( .A(_04670_ ), .ZN(_04671_ ) );
INV_X1 _12432_ ( .A(\ID_EX_pc [4] ), .ZN(_04672_ ) );
XNOR2_X1 _12433_ ( .A(_02841_ ), .B(_04672_ ), .ZN(_04673_ ) );
AOI21_X1 _12434_ ( .A(_04673_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04674_ ) );
XNOR2_X1 _12435_ ( .A(_02735_ ), .B(_02736_ ), .ZN(_04675_ ) );
AOI211_X1 _12436_ ( .A(fanout_net_10 ), .B(_04674_ ), .C1(_04475_ ), .C2(_04675_ ), .ZN(_04676_ ) );
OR3_X1 _12437_ ( .A1(_04120_ ), .A2(_04668_ ), .A3(_04121_ ), .ZN(_04677_ ) );
NAND4_X1 _12438_ ( .A1(_04106_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][4] ), .A4(_04385_ ), .ZN(_04678_ ) );
AND2_X1 _12439_ ( .A1(_04105_ ), .A2(_04678_ ), .ZN(_04679_ ) );
NAND3_X1 _12440_ ( .A1(_04388_ ), .A2(\mepc [4] ), .A3(_04390_ ), .ZN(_04680_ ) );
NAND4_X1 _12441_ ( .A1(_02678_ ), .A2(_02683_ ), .A3(\mtvec [4] ), .A4(_04115_ ), .ZN(_04681_ ) );
NAND4_X1 _12442_ ( .A1(_04397_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_04113_ ), .A4(_04398_ ), .ZN(_04682_ ) );
NAND4_X1 _12443_ ( .A1(_04679_ ), .A2(_04680_ ), .A3(_04681_ ), .A4(_04682_ ), .ZN(_04683_ ) );
OAI21_X1 _12444_ ( .A(_04683_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04684_ ) );
AOI21_X1 _12445_ ( .A(_04644_ ), .B1(_04677_ ), .B2(_04684_ ), .ZN(_04685_ ) );
OAI21_X1 _12446_ ( .A(_04499_ ), .B1(_04676_ ), .B2(_04685_ ), .ZN(_04686_ ) );
AOI21_X1 _12447_ ( .A(_04561_ ), .B1(_04675_ ), .B2(_04512_ ), .ZN(_04687_ ) );
XNOR2_X1 _12448_ ( .A(_02073_ ), .B(_02120_ ), .ZN(_04688_ ) );
OAI21_X1 _12449_ ( .A(_04687_ ), .B1(_04688_ ), .B2(_04427_ ), .ZN(_04689_ ) );
AND2_X1 _12450_ ( .A1(_04689_ ), .A2(_04516_ ), .ZN(_04690_ ) );
AOI221_X1 _12451_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04671_ ), .C1(_04686_ ), .C2(_04690_ ), .ZN(_00139_ ) );
NAND4_X1 _12452_ ( .A1(_02677_ ), .A2(_02681_ ), .A3(\mtvec [3] ), .A4(_04384_ ), .ZN(_04691_ ) );
NAND4_X1 _12453_ ( .A1(_02690_ ), .A2(_02696_ ), .A3(\mepc [3] ), .A4(_02700_ ), .ZN(_04692_ ) );
NAND4_X1 _12454_ ( .A1(_02681_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_02700_ ), .A4(_02702_ ), .ZN(_04693_ ) );
NAND4_X1 _12455_ ( .A1(_02696_ ), .A2(_04140_ ), .A3(\mycsreg.CSReg[3][3] ), .A4(_02700_ ), .ZN(_04694_ ) );
NAND4_X1 _12456_ ( .A1(_04691_ ), .A2(_04692_ ), .A3(_04693_ ), .A4(_04694_ ), .ZN(_04695_ ) );
AOI221_X4 _12457_ ( .A(_04695_ ), .B1(_02691_ ), .B2(_02669_ ), .C1(_02652_ ), .C2(_02663_ ), .ZN(_04696_ ) );
INV_X1 _12458_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_04697_ ) );
AND3_X1 _12459_ ( .A1(_02714_ ), .A2(_04697_ ), .A3(_02716_ ), .ZN(_04698_ ) );
NOR2_X1 _12460_ ( .A1(_04696_ ), .A2(_04698_ ), .ZN(_04699_ ) );
INV_X1 _12461_ ( .A(_04699_ ), .ZN(_04700_ ) );
XOR2_X1 _12462_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .Z(_04701_ ) );
AOI21_X1 _12463_ ( .A(_04701_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04702_ ) );
XOR2_X1 _12464_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_imm [3] ), .Z(_04703_ ) );
XOR2_X1 _12465_ ( .A(_02731_ ), .B(_04703_ ), .Z(_04704_ ) );
INV_X1 _12466_ ( .A(_04704_ ), .ZN(_04705_ ) );
AOI211_X1 _12467_ ( .A(fanout_net_10 ), .B(_04702_ ), .C1(_04475_ ), .C2(_04705_ ), .ZN(_04706_ ) );
OR3_X1 _12468_ ( .A1(_04120_ ), .A2(_04697_ ), .A3(_04121_ ), .ZN(_04707_ ) );
NAND4_X1 _12469_ ( .A1(_04106_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][3] ), .A4(_04385_ ), .ZN(_04708_ ) );
AND2_X1 _12470_ ( .A1(_04105_ ), .A2(_04708_ ), .ZN(_04709_ ) );
NAND3_X1 _12471_ ( .A1(_04111_ ), .A2(\mepc [3] ), .A3(_04390_ ), .ZN(_04710_ ) );
NAND4_X1 _12472_ ( .A1(_02678_ ), .A2(_02683_ ), .A3(\mtvec [3] ), .A4(_04115_ ), .ZN(_04711_ ) );
NAND4_X1 _12473_ ( .A1(_04397_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_04394_ ), .A4(_04398_ ), .ZN(_04712_ ) );
NAND4_X1 _12474_ ( .A1(_04709_ ), .A2(_04710_ ), .A3(_04711_ ), .A4(_04712_ ), .ZN(_04713_ ) );
OAI21_X1 _12475_ ( .A(_04713_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04714_ ) );
AOI21_X1 _12476_ ( .A(_04644_ ), .B1(_04707_ ), .B2(_04714_ ), .ZN(_04715_ ) );
OAI21_X1 _12477_ ( .A(_04499_ ), .B1(_04706_ ), .B2(_04715_ ), .ZN(_04716_ ) );
AOI21_X1 _12478_ ( .A(_04561_ ), .B1(_04705_ ), .B2(_04512_ ), .ZN(_04717_ ) );
XOR2_X1 _12479_ ( .A(_02047_ ), .B(_02070_ ), .Z(_04718_ ) );
OAI21_X1 _12480_ ( .A(_04717_ ), .B1(_04718_ ), .B2(_04427_ ), .ZN(_04719_ ) );
AND2_X1 _12481_ ( .A1(_04719_ ), .A2(_04516_ ), .ZN(_04720_ ) );
AOI221_X1 _12482_ ( .A(fanout_net_2 ), .B1(_04430_ ), .B2(_04700_ ), .C1(_04716_ ), .C2(_04720_ ), .ZN(_00140_ ) );
NAND4_X1 _12483_ ( .A1(_04231_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][2] ), .A4(_04389_ ), .ZN(_04721_ ) );
NAND3_X1 _12484_ ( .A1(_04111_ ), .A2(\mepc [2] ), .A3(_04205_ ), .ZN(_04722_ ) );
NAND4_X1 _12485_ ( .A1(_04203_ ), .A2(_04396_ ), .A3(\mtvec [2] ), .A4(_04385_ ), .ZN(_04723_ ) );
NAND4_X1 _12486_ ( .A1(_04167_ ), .A2(_04721_ ), .A3(_04722_ ), .A4(_04723_ ), .ZN(_04724_ ) );
AND4_X1 _12487_ ( .A1(\mycsreg.CSReg[0][2] ), .A2(_04396_ ), .A3(_04205_ ), .A4(_04117_ ), .ZN(_04725_ ) );
OAI21_X1 _12488_ ( .A(_02665_ ), .B1(_04724_ ), .B2(_04725_ ), .ZN(_04726_ ) );
NAND3_X1 _12489_ ( .A1(_04365_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_04366_ ), .ZN(_04727_ ) );
AND2_X1 _12490_ ( .A1(_04726_ ), .A2(_04727_ ), .ZN(_04728_ ) );
AOI21_X1 _12491_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04729_ ) );
NOR2_X1 _12492_ ( .A1(_02727_ ), .A2(_02728_ ), .ZN(_04730_ ) );
XNOR2_X1 _12493_ ( .A(_04730_ ), .B(_02724_ ), .ZN(_04731_ ) );
INV_X1 _12494_ ( .A(_04731_ ), .ZN(_04732_ ) );
AOI211_X1 _12495_ ( .A(fanout_net_10 ), .B(_04729_ ), .C1(_04475_ ), .C2(_04732_ ), .ZN(_04733_ ) );
INV_X1 _12496_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_04734_ ) );
OR3_X1 _12497_ ( .A1(_04101_ ), .A2(_04734_ ), .A3(_01677_ ), .ZN(_04735_ ) );
AOI21_X1 _12498_ ( .A(_04644_ ), .B1(_04726_ ), .B2(_04735_ ), .ZN(_04736_ ) );
OAI21_X1 _12499_ ( .A(_04499_ ), .B1(_04733_ ), .B2(_04736_ ), .ZN(_04737_ ) );
AOI21_X1 _12500_ ( .A(_04561_ ), .B1(_04732_ ), .B2(_04512_ ), .ZN(_04738_ ) );
XNOR2_X1 _12501_ ( .A(_02043_ ), .B(_02046_ ), .ZN(_04739_ ) );
OAI21_X1 _12502_ ( .A(_04738_ ), .B1(_04739_ ), .B2(_04427_ ), .ZN(_04740_ ) );
AND2_X1 _12503_ ( .A1(_04740_ ), .A2(_04516_ ), .ZN(_04741_ ) );
AOI221_X1 _12504_ ( .A(fanout_net_2 ), .B1(_04225_ ), .B2(_04728_ ), .C1(_04737_ ), .C2(_04741_ ), .ZN(_00141_ ) );
NAND4_X1 _12505_ ( .A1(_04169_ ), .A2(_04233_ ), .A3(\mtvec [1] ), .A4(_02709_ ), .ZN(_04742_ ) );
NAND4_X1 _12506_ ( .A1(_04256_ ), .A2(_02697_ ), .A3(\mepc [1] ), .A4(_04170_ ), .ZN(_04743_ ) );
NAND4_X1 _12507_ ( .A1(_04133_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_04174_ ), .A4(_04136_ ), .ZN(_04744_ ) );
NAND4_X1 _12508_ ( .A1(_02697_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][1] ), .A4(_04134_ ), .ZN(_04745_ ) );
AND4_X1 _12509_ ( .A1(_04742_ ), .A2(_04743_ ), .A3(_04744_ ), .A4(_04745_ ), .ZN(_04746_ ) );
OR2_X1 _12510_ ( .A1(_02664_ ), .A2(_04746_ ), .ZN(_04747_ ) );
NAND3_X1 _12511_ ( .A1(_04365_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_04366_ ), .ZN(_04748_ ) );
AND2_X1 _12512_ ( .A1(_04747_ ), .A2(_04748_ ), .ZN(_04749_ ) );
AOI21_X1 _12513_ ( .A(\ID_EX_pc [1] ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04750_ ) );
XOR2_X1 _12514_ ( .A(_02725_ ), .B(_02726_ ), .Z(_04751_ ) );
INV_X1 _12515_ ( .A(_04751_ ), .ZN(_04752_ ) );
AOI211_X1 _12516_ ( .A(fanout_net_10 ), .B(_04750_ ), .C1(_04475_ ), .C2(_04752_ ), .ZN(_04753_ ) );
INV_X1 _12517_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_04754_ ) );
OR3_X1 _12518_ ( .A1(_04120_ ), .A2(_04754_ ), .A3(_04121_ ), .ZN(_04755_ ) );
NAND3_X1 _12519_ ( .A1(_04388_ ), .A2(\mepc [1] ), .A3(_04390_ ), .ZN(_04756_ ) );
NAND4_X1 _12520_ ( .A1(_04392_ ), .A2(_04393_ ), .A3(\mtvec [1] ), .A4(_04113_ ), .ZN(_04757_ ) );
NAND4_X1 _12521_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][1] ), .A4(_04115_ ), .ZN(_04758_ ) );
NAND4_X1 _12522_ ( .A1(_04393_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_04394_ ), .A4(_04398_ ), .ZN(_04759_ ) );
NAND4_X1 _12523_ ( .A1(_04756_ ), .A2(_04757_ ), .A3(_04758_ ), .A4(_04759_ ), .ZN(_04760_ ) );
OAI21_X1 _12524_ ( .A(_04760_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04761_ ) );
AOI21_X1 _12525_ ( .A(_04644_ ), .B1(_04755_ ), .B2(_04761_ ), .ZN(_04762_ ) );
OAI21_X1 _12526_ ( .A(_04499_ ), .B1(_04753_ ), .B2(_04762_ ), .ZN(_04763_ ) );
AOI21_X1 _12527_ ( .A(_04561_ ), .B1(_04752_ ), .B2(_04512_ ), .ZN(_04764_ ) );
XOR2_X1 _12528_ ( .A(_02016_ ), .B(_02039_ ), .Z(_04765_ ) );
OAI21_X1 _12529_ ( .A(_04764_ ), .B1(_04765_ ), .B2(_04427_ ), .ZN(_04766_ ) );
AND2_X1 _12530_ ( .A1(_04766_ ), .A2(_04516_ ), .ZN(_04767_ ) );
AOI221_X1 _12531_ ( .A(fanout_net_2 ), .B1(_04225_ ), .B2(_04749_ ), .C1(_04763_ ), .C2(_04767_ ), .ZN(_00142_ ) );
NAND3_X1 _12532_ ( .A1(_04331_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_04332_ ), .ZN(_04768_ ) );
NAND3_X1 _12533_ ( .A1(_04111_ ), .A2(\mepc [27] ), .A3(_04389_ ), .ZN(_04769_ ) );
NAND2_X1 _12534_ ( .A1(_04768_ ), .A2(_04769_ ), .ZN(_04770_ ) );
AND4_X1 _12535_ ( .A1(\mycsreg.CSReg[3][27] ), .A2(_04106_ ), .A3(_02708_ ), .A4(_04112_ ), .ZN(_04771_ ) );
NOR3_X1 _12536_ ( .A1(_02675_ ), .A2(_04770_ ), .A3(_04771_ ), .ZN(_04772_ ) );
NAND2_X1 _12537_ ( .A1(_04341_ ), .A2(\mtvec [27] ), .ZN(_04773_ ) );
OAI211_X1 _12538_ ( .A(_04772_ ), .B(_04773_ ), .C1(_04262_ ), .C2(_04264_ ), .ZN(_04774_ ) );
INV_X1 _12539_ ( .A(\EX_LS_result_csreg_mem [27] ), .ZN(_04775_ ) );
NAND3_X1 _12540_ ( .A1(_04181_ ), .A2(_04775_ ), .A3(_04183_ ), .ZN(_04776_ ) );
NAND2_X1 _12541_ ( .A1(_04774_ ), .A2(_04776_ ), .ZN(_04777_ ) );
NAND3_X1 _12542_ ( .A1(_04148_ ), .A2(\ID_EX_pc [26] ), .A3(_04151_ ), .ZN(_04778_ ) );
XNOR2_X1 _12543_ ( .A(_04778_ ), .B(\ID_EX_pc [27] ), .ZN(_04779_ ) );
AOI21_X1 _12544_ ( .A(_04779_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04780_ ) );
NAND2_X1 _12545_ ( .A1(_02815_ ), .A2(_02817_ ), .ZN(_04781_ ) );
NAND2_X1 _12546_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_04782_ ) );
NAND2_X1 _12547_ ( .A1(_04781_ ), .A2(_04782_ ), .ZN(_04783_ ) );
XNOR2_X1 _12548_ ( .A(_04783_ ), .B(_02816_ ), .ZN(_04784_ ) );
AOI211_X1 _12549_ ( .A(\ID_EX_typ [3] ), .B(_04780_ ), .C1(_04475_ ), .C2(_04784_ ), .ZN(_04785_ ) );
OR3_X1 _12550_ ( .A1(_04101_ ), .A2(_04775_ ), .A3(_01677_ ), .ZN(_04786_ ) );
NAND4_X1 _12551_ ( .A1(_04106_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][27] ), .A4(_04385_ ), .ZN(_04787_ ) );
AND2_X1 _12552_ ( .A1(_04105_ ), .A2(_04787_ ), .ZN(_04788_ ) );
NAND4_X1 _12553_ ( .A1(_02678_ ), .A2(_02683_ ), .A3(\mtvec [27] ), .A4(_04115_ ), .ZN(_04789_ ) );
NAND4_X1 _12554_ ( .A1(_04393_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_04394_ ), .A4(_04398_ ), .ZN(_04790_ ) );
NAND4_X1 _12555_ ( .A1(_04788_ ), .A2(_04769_ ), .A3(_04789_ ), .A4(_04790_ ), .ZN(_04791_ ) );
OAI21_X1 _12556_ ( .A(_04791_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04792_ ) );
AOI21_X1 _12557_ ( .A(_04644_ ), .B1(_04786_ ), .B2(_04792_ ), .ZN(_04793_ ) );
OAI21_X1 _12558_ ( .A(_04499_ ), .B1(_04785_ ), .B2(_04793_ ), .ZN(_04794_ ) );
NAND2_X1 _12559_ ( .A1(_02623_ ), .A2(fanout_net_8 ), .ZN(_04795_ ) );
AOI21_X1 _12560_ ( .A(_02720_ ), .B1(_04784_ ), .B2(_02835_ ), .ZN(_04796_ ) );
AOI21_X1 _12561_ ( .A(_04283_ ), .B1(_04795_ ), .B2(_04796_ ), .ZN(_04797_ ) );
AOI221_X1 _12562_ ( .A(fanout_net_2 ), .B1(_04225_ ), .B2(_04777_ ), .C1(_04794_ ), .C2(_04797_ ), .ZN(_00143_ ) );
XOR2_X1 _12563_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_04798_ ) );
OAI21_X1 _12564_ ( .A(_04086_ ), .B1(_04268_ ), .B2(_04798_ ), .ZN(_04799_ ) );
INV_X1 _12565_ ( .A(\ID_EX_pc [0] ), .ZN(_04800_ ) );
AOI21_X1 _12566_ ( .A(_04799_ ), .B1(_04800_ ), .B2(_04268_ ), .ZN(_04801_ ) );
AND4_X1 _12567_ ( .A1(\mtvec [0] ), .A2(_04169_ ), .A3(_04133_ ), .A4(_04170_ ), .ZN(_04802_ ) );
NAND4_X1 _12568_ ( .A1(_02690_ ), .A2(_04138_ ), .A3(\mepc [0] ), .A4(_02687_ ), .ZN(_04803_ ) );
NAND4_X1 _12569_ ( .A1(_04138_ ), .A2(_04140_ ), .A3(\mycsreg.CSReg[3][0] ), .A4(_02687_ ), .ZN(_04804_ ) );
NAND4_X1 _12570_ ( .A1(_02681_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_02687_ ), .A4(_04136_ ), .ZN(_04805_ ) );
NAND4_X1 _12571_ ( .A1(_04167_ ), .A2(_04803_ ), .A3(_04804_ ), .A4(_04805_ ), .ZN(_04806_ ) );
OAI21_X1 _12572_ ( .A(_02665_ ), .B1(_04802_ ), .B2(_04806_ ), .ZN(_04807_ ) );
INV_X1 _12573_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_04808_ ) );
OR3_X1 _12574_ ( .A1(_04101_ ), .A2(_04808_ ), .A3(_01677_ ), .ZN(_04809_ ) );
AOI21_X1 _12575_ ( .A(_04644_ ), .B1(_04807_ ), .B2(_04809_ ), .ZN(_04810_ ) );
OAI21_X1 _12576_ ( .A(_02840_ ), .B1(_04801_ ), .B2(_04810_ ), .ZN(_04811_ ) );
BUF_X4 _12577_ ( .A(_02837_ ), .Z(_04812_ ) );
NAND4_X1 _12578_ ( .A1(_04798_ ), .A2(\ID_EX_typ [7] ), .A3(\myexu.pc_jump_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_A ), .A4(_01648_ ), .ZN(_04813_ ) );
AND3_X2 _12579_ ( .A1(_04811_ ), .A2(_04812_ ), .A3(_04813_ ), .ZN(_04814_ ) );
NAND3_X1 _12580_ ( .A1(_02714_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_02716_ ), .ZN(_04815_ ) );
AND2_X1 _12581_ ( .A1(_04807_ ), .A2(_04815_ ), .ZN(_04816_ ) );
AOI211_X1 _12582_ ( .A(fanout_net_2 ), .B(_04814_ ), .C1(_04163_ ), .C2(_04816_ ), .ZN(_00144_ ) );
NAND4_X1 _12583_ ( .A1(_04169_ ), .A2(_04233_ ), .A3(\mtvec [26] ), .A4(_02709_ ), .ZN(_04817_ ) );
NAND4_X1 _12584_ ( .A1(_04256_ ), .A2(_04172_ ), .A3(\mepc [26] ), .A4(_04170_ ), .ZN(_04818_ ) );
NAND4_X1 _12585_ ( .A1(_04233_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_04170_ ), .A4(_04136_ ), .ZN(_04819_ ) );
NAND4_X1 _12586_ ( .A1(_04172_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][26] ), .A4(_04174_ ), .ZN(_04820_ ) );
AND4_X1 _12587_ ( .A1(_04817_ ), .A2(_04818_ ), .A3(_04819_ ), .A4(_04820_ ), .ZN(_04821_ ) );
OR2_X1 _12588_ ( .A1(_02664_ ), .A2(_04821_ ), .ZN(_04822_ ) );
NAND3_X1 _12589_ ( .A1(_02715_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_02717_ ), .ZN(_04823_ ) );
AND2_X1 _12590_ ( .A1(_04822_ ), .A2(_04823_ ), .ZN(_04824_ ) );
XNOR2_X1 _12591_ ( .A(_04152_ ), .B(_04154_ ), .ZN(_04825_ ) );
AND2_X2 _12592_ ( .A1(_04268_ ), .A2(_04825_ ), .ZN(_04826_ ) );
XNOR2_X1 _12593_ ( .A(_02815_ ), .B(_02817_ ), .ZN(_04827_ ) );
AOI211_X2 _12594_ ( .A(\ID_EX_typ [3] ), .B(_04826_ ), .C1(_04084_ ), .C2(_04827_ ), .ZN(_04828_ ) );
NAND2_X1 _12595_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [26] ), .ZN(_04829_ ) );
NAND3_X1 _12596_ ( .A1(_04388_ ), .A2(\mepc [26] ), .A3(_04390_ ), .ZN(_04830_ ) );
NAND4_X1 _12597_ ( .A1(_04392_ ), .A2(_04393_ ), .A3(\mtvec [26] ), .A4(_04113_ ), .ZN(_04831_ ) );
NAND4_X1 _12598_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][26] ), .A4(_04115_ ), .ZN(_04832_ ) );
NAND4_X1 _12599_ ( .A1(_04393_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_04394_ ), .A4(_04398_ ), .ZN(_04833_ ) );
NAND4_X1 _12600_ ( .A1(_04830_ ), .A2(_04831_ ), .A3(_04832_ ), .A4(_04833_ ), .ZN(_04834_ ) );
OAI21_X1 _12601_ ( .A(_04834_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04835_ ) );
AOI21_X1 _12602_ ( .A(_04644_ ), .B1(_04829_ ), .B2(_04835_ ), .ZN(_04836_ ) );
OAI21_X1 _12603_ ( .A(_04499_ ), .B1(_04828_ ), .B2(_04836_ ), .ZN(_04837_ ) );
AOI21_X1 _12604_ ( .A(_04561_ ), .B1(_04827_ ), .B2(_04512_ ), .ZN(_04838_ ) );
OAI21_X1 _12605_ ( .A(_04838_ ), .B1(_02624_ ), .B2(_04427_ ), .ZN(_04839_ ) );
AND2_X1 _12606_ ( .A1(_04839_ ), .A2(_04516_ ), .ZN(_04840_ ) );
AOI221_X1 _12607_ ( .A(fanout_net_3 ), .B1(_04225_ ), .B2(_04824_ ), .C1(_04837_ ), .C2(_04840_ ), .ZN(_00145_ ) );
AND3_X1 _12608_ ( .A1(_04365_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_04366_ ), .ZN(_04841_ ) );
NAND4_X1 _12609_ ( .A1(_04204_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_04205_ ), .A4(_04117_ ), .ZN(_04842_ ) );
NAND4_X1 _12610_ ( .A1(_04231_ ), .A2(_04383_ ), .A3(\mycsreg.CSReg[3][25] ), .A4(_04389_ ), .ZN(_04843_ ) );
NAND4_X1 _12611_ ( .A1(_02691_ ), .A2(_04106_ ), .A3(\mepc [25] ), .A4(_04389_ ), .ZN(_04844_ ) );
AND3_X1 _12612_ ( .A1(_04842_ ), .A2(_04843_ ), .A3(_04844_ ), .ZN(_04845_ ) );
NAND4_X1 _12613_ ( .A1(_04392_ ), .A2(_04397_ ), .A3(\mtvec [25] ), .A4(_04571_ ), .ZN(_04846_ ) );
AOI22_X1 _12614_ ( .A1(_02715_ ), .A2(_02717_ ), .B1(_04845_ ), .B2(_04846_ ), .ZN(_04847_ ) );
NOR2_X1 _12615_ ( .A1(_04841_ ), .A2(_04847_ ), .ZN(_04848_ ) );
AND3_X1 _12616_ ( .A1(_04150_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_04849_ ) );
AND2_X1 _12617_ ( .A1(_04148_ ), .A2(_04849_ ), .ZN(_04850_ ) );
NAND3_X1 _12618_ ( .A1(_04850_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_04851_ ) );
INV_X1 _12619_ ( .A(\ID_EX_pc [24] ), .ZN(_04852_ ) );
NOR2_X1 _12620_ ( .A1(_04851_ ), .A2(_04852_ ), .ZN(_04853_ ) );
INV_X1 _12621_ ( .A(\ID_EX_pc [25] ), .ZN(_04854_ ) );
XNOR2_X1 _12622_ ( .A(_04853_ ), .B(_04854_ ), .ZN(_04855_ ) );
AOI21_X1 _12623_ ( .A(_04855_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04856_ ) );
AND2_X1 _12624_ ( .A1(_02808_ ), .A2(_02810_ ), .ZN(_04857_ ) );
OR2_X1 _12625_ ( .A1(_04857_ ), .A2(_02812_ ), .ZN(_04858_ ) );
XNOR2_X1 _12626_ ( .A(_04858_ ), .B(_02809_ ), .ZN(_04859_ ) );
AOI211_X1 _12627_ ( .A(\ID_EX_typ [3] ), .B(_04856_ ), .C1(_04084_ ), .C2(_04859_ ), .ZN(_04860_ ) );
NAND2_X1 _12628_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [25] ), .ZN(_04861_ ) );
NAND3_X1 _12629_ ( .A1(_04388_ ), .A2(\mepc [25] ), .A3(_04390_ ), .ZN(_04862_ ) );
NAND4_X1 _12630_ ( .A1(_04392_ ), .A2(_04393_ ), .A3(\mtvec [25] ), .A4(_04113_ ), .ZN(_04863_ ) );
NAND4_X1 _12631_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][25] ), .A4(_04115_ ), .ZN(_04864_ ) );
NAND4_X1 _12632_ ( .A1(_04393_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_04394_ ), .A4(_04117_ ), .ZN(_04865_ ) );
NAND4_X1 _12633_ ( .A1(_04862_ ), .A2(_04863_ ), .A3(_04864_ ), .A4(_04865_ ), .ZN(_04866_ ) );
OAI21_X1 _12634_ ( .A(_04866_ ), .B1(_04120_ ), .B2(_04121_ ), .ZN(_04867_ ) );
AOI21_X1 _12635_ ( .A(_04644_ ), .B1(_04861_ ), .B2(_04867_ ), .ZN(_04868_ ) );
OAI21_X1 _12636_ ( .A(_02840_ ), .B1(_04860_ ), .B2(_04868_ ), .ZN(_04869_ ) );
AOI21_X1 _12637_ ( .A(_04561_ ), .B1(_04859_ ), .B2(_04512_ ), .ZN(_04870_ ) );
OAI21_X1 _12638_ ( .A(_04870_ ), .B1(_02627_ ), .B2(_04427_ ), .ZN(_04871_ ) );
AND2_X1 _12639_ ( .A1(_04871_ ), .A2(_04516_ ), .ZN(_04872_ ) );
AOI221_X1 _12640_ ( .A(fanout_net_3 ), .B1(_04225_ ), .B2(_04848_ ), .C1(_04869_ ), .C2(_04872_ ), .ZN(_00146_ ) );
NAND4_X1 _12641_ ( .A1(_04169_ ), .A2(_02682_ ), .A3(\mtvec [24] ), .A4(_02701_ ), .ZN(_04873_ ) );
NAND4_X1 _12642_ ( .A1(_04256_ ), .A2(_04172_ ), .A3(\mepc [24] ), .A4(_02709_ ), .ZN(_04874_ ) );
NAND4_X1 _12643_ ( .A1(_04233_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_02709_ ), .A4(_02703_ ), .ZN(_04875_ ) );
NAND4_X1 _12644_ ( .A1(_04172_ ), .A2(_04173_ ), .A3(\mycsreg.CSReg[3][24] ), .A4(_04170_ ), .ZN(_04876_ ) );
AND4_X1 _12645_ ( .A1(_04873_ ), .A2(_04874_ ), .A3(_04875_ ), .A4(_04876_ ), .ZN(_04877_ ) );
NAND3_X1 _12646_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04877_ ), .ZN(_04878_ ) );
OR3_X1 _12647_ ( .A1(_04262_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_04264_ ), .ZN(_04879_ ) );
AND2_X1 _12648_ ( .A1(_04878_ ), .A2(_04879_ ), .ZN(_04880_ ) );
INV_X1 _12649_ ( .A(_04880_ ), .ZN(_04881_ ) );
XNOR2_X1 _12650_ ( .A(_04851_ ), .B(\ID_EX_pc [24] ), .ZN(_04882_ ) );
AOI21_X1 _12651_ ( .A(_04882_ ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_04883_ ) );
XNOR2_X1 _12652_ ( .A(_02808_ ), .B(_02810_ ), .ZN(_04884_ ) );
AOI211_X1 _12653_ ( .A(\ID_EX_typ [3] ), .B(_04883_ ), .C1(_04084_ ), .C2(_04884_ ), .ZN(_04885_ ) );
AND3_X1 _12654_ ( .A1(_04878_ ), .A2(\ID_EX_typ [3] ), .A3(_04879_ ), .ZN(_04886_ ) );
OAI21_X1 _12655_ ( .A(_02840_ ), .B1(_04885_ ), .B2(_04886_ ), .ZN(_04887_ ) );
AOI21_X1 _12656_ ( .A(_04561_ ), .B1(_04884_ ), .B2(_04512_ ), .ZN(_04888_ ) );
OAI21_X1 _12657_ ( .A(_04888_ ), .B1(_02628_ ), .B2(_02833_ ), .ZN(_04889_ ) );
AND2_X1 _12658_ ( .A1(_04889_ ), .A2(_04516_ ), .ZN(_04890_ ) );
AOI221_X1 _12659_ ( .A(fanout_net_3 ), .B1(_04225_ ), .B2(_04881_ ), .C1(_04887_ ), .C2(_04890_ ), .ZN(_00147_ ) );
INV_X1 _12660_ ( .A(_02794_ ), .ZN(_04891_ ) );
OAI21_X1 _12661_ ( .A(_02797_ ), .B1(_02783_ ), .B2(_02791_ ), .ZN(_04892_ ) );
AOI21_X1 _12662_ ( .A(_04891_ ), .B1(_04892_ ), .B2(_02801_ ), .ZN(_04893_ ) );
NOR2_X1 _12663_ ( .A1(_04893_ ), .A2(_02805_ ), .ZN(_04894_ ) );
XNOR2_X1 _12664_ ( .A(_04894_ ), .B(_02793_ ), .ZN(_04895_ ) );
OAI21_X1 _12665_ ( .A(_01649_ ), .B1(_04895_ ), .B2(fanout_net_8 ), .ZN(_04896_ ) );
AOI21_X1 _12666_ ( .A(_04896_ ), .B1(_02635_ ), .B2(fanout_net_8 ), .ZN(_04897_ ) );
AND3_X1 _12667_ ( .A1(_02652_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_02663_ ), .ZN(_04898_ ) );
NAND4_X1 _12668_ ( .A1(_02690_ ), .A2(_04138_ ), .A3(\mepc [23] ), .A4(_04384_ ), .ZN(_04899_ ) );
NAND4_X1 _12669_ ( .A1(_02681_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_04384_ ), .A4(_02702_ ), .ZN(_04900_ ) );
NAND4_X1 _12670_ ( .A1(_02696_ ), .A2(_04140_ ), .A3(\mycsreg.CSReg[3][23] ), .A4(_02700_ ), .ZN(_04901_ ) );
AND3_X1 _12671_ ( .A1(_04899_ ), .A2(_04900_ ), .A3(_04901_ ), .ZN(_04902_ ) );
NAND4_X1 _12672_ ( .A1(_04203_ ), .A2(_04396_ ), .A3(\mtvec [23] ), .A4(_04385_ ), .ZN(_04903_ ) );
AOI22_X1 _12673_ ( .A1(_02714_ ), .A2(_02716_ ), .B1(_04902_ ), .B2(_04903_ ), .ZN(_04904_ ) );
NOR2_X1 _12674_ ( .A1(_04898_ ), .A2(_04904_ ), .ZN(_04905_ ) );
INV_X1 _12675_ ( .A(_04905_ ), .ZN(_04906_ ) );
NAND3_X1 _12676_ ( .A1(_04148_ ), .A2(\ID_EX_pc [22] ), .A3(_04849_ ), .ZN(_04907_ ) );
XNOR2_X1 _12677_ ( .A(_04907_ ), .B(\ID_EX_pc [23] ), .ZN(_04908_ ) );
MUX2_X1 _12678_ ( .A(_04908_ ), .B(_04895_ ), .S(_04083_ ), .Z(_04909_ ) );
MUX2_X2 _12679_ ( .A(_04906_ ), .B(_04909_ ), .S(_04159_ ), .Z(_04910_ ) );
AOI211_X1 _12680_ ( .A(_04125_ ), .B(_04897_ ), .C1(_04910_ ), .C2(_04161_ ), .ZN(_04911_ ) );
AOI211_X1 _12681_ ( .A(fanout_net_3 ), .B(_04911_ ), .C1(_04163_ ), .C2(_04905_ ), .ZN(_00148_ ) );
NAND4_X1 _12682_ ( .A1(_04169_ ), .A2(_04133_ ), .A3(\mtvec [22] ), .A4(_04174_ ), .ZN(_04912_ ) );
NAND4_X1 _12683_ ( .A1(_04133_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_04134_ ), .A4(_04136_ ), .ZN(_04913_ ) );
NAND4_X1 _12684_ ( .A1(_02697_ ), .A2(_04140_ ), .A3(\mycsreg.CSReg[3][22] ), .A4(_04134_ ), .ZN(_04914_ ) );
NAND4_X1 _12685_ ( .A1(_02690_ ), .A2(_04138_ ), .A3(\mepc [22] ), .A4(_02687_ ), .ZN(_04915_ ) );
AND4_X1 _12686_ ( .A1(_04912_ ), .A2(_04913_ ), .A3(_04914_ ), .A4(_04915_ ), .ZN(_04916_ ) );
NAND3_X1 _12687_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04916_ ), .ZN(_04917_ ) );
OR3_X1 _12688_ ( .A1(_04261_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_04263_ ), .ZN(_04918_ ) );
AND2_X1 _12689_ ( .A1(_04917_ ), .A2(_04918_ ), .ZN(_04919_ ) );
INV_X1 _12690_ ( .A(_04919_ ), .ZN(_04920_ ) );
XNOR2_X1 _12691_ ( .A(_04850_ ), .B(\ID_EX_pc [22] ), .ZN(_04921_ ) );
AND2_X2 _12692_ ( .A1(_04268_ ), .A2(_04921_ ), .ZN(_04922_ ) );
NAND2_X1 _12693_ ( .A1(_04892_ ), .A2(_02801_ ), .ZN(_04923_ ) );
XNOR2_X1 _12694_ ( .A(_04923_ ), .B(_04891_ ), .ZN(_04924_ ) );
INV_X1 _12695_ ( .A(_04924_ ), .ZN(_04925_ ) );
AOI211_X2 _12696_ ( .A(\ID_EX_typ [3] ), .B(_04922_ ), .C1(_04084_ ), .C2(_04925_ ), .ZN(_04926_ ) );
NAND3_X1 _12697_ ( .A1(_04917_ ), .A2(\ID_EX_typ [3] ), .A3(_04918_ ), .ZN(_04927_ ) );
INV_X1 _12698_ ( .A(_04927_ ), .ZN(_04928_ ) );
OAI21_X1 _12699_ ( .A(_02840_ ), .B1(_04926_ ), .B2(_04928_ ), .ZN(_04929_ ) );
AOI21_X1 _12700_ ( .A(_04561_ ), .B1(_04925_ ), .B2(_04512_ ), .ZN(_04930_ ) );
AND2_X1 _12701_ ( .A1(_02636_ ), .A2(_02631_ ), .ZN(_04931_ ) );
OAI21_X1 _12702_ ( .A(_04930_ ), .B1(_04931_ ), .B2(_02833_ ), .ZN(_04932_ ) );
AND2_X1 _12703_ ( .A1(_04932_ ), .A2(_04516_ ), .ZN(_04933_ ) );
AOI221_X1 _12704_ ( .A(fanout_net_3 ), .B1(_04225_ ), .B2(_04920_ ), .C1(_04929_ ), .C2(_04933_ ), .ZN(_00149_ ) );
NAND4_X1 _12705_ ( .A1(_04203_ ), .A2(_04396_ ), .A3(\mtvec [21] ), .A4(_04112_ ), .ZN(_04934_ ) );
NAND4_X1 _12706_ ( .A1(_02691_ ), .A2(_02705_ ), .A3(\mepc [21] ), .A4(_04107_ ), .ZN(_04935_ ) );
NAND4_X1 _12707_ ( .A1(_02682_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_04107_ ), .A4(_02703_ ), .ZN(_04936_ ) );
NAND4_X1 _12708_ ( .A1(_02705_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][21] ), .A4(_02701_ ), .ZN(_04937_ ) );
NAND4_X1 _12709_ ( .A1(_04934_ ), .A2(_04935_ ), .A3(_04936_ ), .A4(_04937_ ), .ZN(_04938_ ) );
AOI211_X1 _12710_ ( .A(_02675_ ), .B(_04938_ ), .C1(_04365_ ), .C2(_04366_ ), .ZN(_04939_ ) );
INV_X1 _12711_ ( .A(\EX_LS_result_csreg_mem [21] ), .ZN(_04940_ ) );
AND3_X1 _12712_ ( .A1(_02714_ ), .A2(_04940_ ), .A3(_02716_ ), .ZN(_04941_ ) );
NOR2_X1 _12713_ ( .A1(_04939_ ), .A2(_04941_ ), .ZN(_04942_ ) );
INV_X1 _12714_ ( .A(_04942_ ), .ZN(_04943_ ) );
INV_X1 _12715_ ( .A(\ID_EX_pc [20] ), .ZN(_04944_ ) );
NOR2_X1 _12716_ ( .A1(_04187_ ), .A2(_04944_ ), .ZN(_04945_ ) );
INV_X1 _12717_ ( .A(\ID_EX_pc [21] ), .ZN(_04946_ ) );
XNOR2_X1 _12718_ ( .A(_04945_ ), .B(_04946_ ), .ZN(_04947_ ) );
AOI21_X1 _12719_ ( .A(_04947_ ), .B1(_04078_ ), .B2(_04081_ ), .ZN(_04948_ ) );
AND2_X1 _12720_ ( .A1(_02792_ ), .A2(_02795_ ), .ZN(_04949_ ) );
OR2_X1 _12721_ ( .A1(_04949_ ), .A2(_02799_ ), .ZN(_04950_ ) );
XNOR2_X1 _12722_ ( .A(_04950_ ), .B(_02796_ ), .ZN(_04951_ ) );
AOI211_X1 _12723_ ( .A(\ID_EX_typ [3] ), .B(_04948_ ), .C1(_04084_ ), .C2(_04951_ ), .ZN(_04952_ ) );
OR3_X1 _12724_ ( .A1(_04101_ ), .A2(_04940_ ), .A3(_01677_ ), .ZN(_04953_ ) );
NAND4_X1 _12725_ ( .A1(_04106_ ), .A2(_02708_ ), .A3(\mycsreg.CSReg[3][21] ), .A4(_04112_ ), .ZN(_04954_ ) );
AND2_X1 _12726_ ( .A1(_04105_ ), .A2(_04954_ ), .ZN(_04955_ ) );
NAND3_X1 _12727_ ( .A1(_04111_ ), .A2(\mepc [21] ), .A3(_04390_ ), .ZN(_04956_ ) );
NAND4_X1 _12728_ ( .A1(_02678_ ), .A2(_02683_ ), .A3(\mtvec [21] ), .A4(_04115_ ), .ZN(_04957_ ) );
NAND4_X1 _12729_ ( .A1(_04393_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_04394_ ), .A4(_04117_ ), .ZN(_04958_ ) );
NAND4_X1 _12730_ ( .A1(_04955_ ), .A2(_04956_ ), .A3(_04957_ ), .A4(_04958_ ), .ZN(_04959_ ) );
OAI21_X1 _12731_ ( .A(_04959_ ), .B1(_04120_ ), .B2(_04121_ ), .ZN(_04960_ ) );
AOI21_X1 _12732_ ( .A(_04644_ ), .B1(_04953_ ), .B2(_04960_ ), .ZN(_04961_ ) );
OAI21_X1 _12733_ ( .A(_02840_ ), .B1(_04952_ ), .B2(_04961_ ), .ZN(_04962_ ) );
AOI21_X1 _12734_ ( .A(_04561_ ), .B1(_04951_ ), .B2(_02832_ ), .ZN(_04963_ ) );
OAI21_X1 _12735_ ( .A(_04963_ ), .B1(_02590_ ), .B2(_02833_ ), .ZN(_04964_ ) );
AND2_X1 _12736_ ( .A1(_04964_ ), .A2(_02837_ ), .ZN(_04965_ ) );
AOI221_X1 _12737_ ( .A(fanout_net_3 ), .B1(_04225_ ), .B2(_04943_ ), .C1(_04962_ ), .C2(_04965_ ), .ZN(_00150_ ) );
NAND2_X1 _12738_ ( .A1(_04102_ ), .A2(\EX_LS_result_csreg_mem [31] ), .ZN(_04966_ ) );
NAND3_X1 _12739_ ( .A1(_04388_ ), .A2(\mepc [31] ), .A3(_04571_ ), .ZN(_04967_ ) );
NAND4_X1 _12740_ ( .A1(_04392_ ), .A2(_04397_ ), .A3(\mtvec [31] ), .A4(_04571_ ), .ZN(_04968_ ) );
NAND4_X1 _12741_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][31] ), .A4(_04571_ ), .ZN(_04969_ ) );
NAND4_X1 _12742_ ( .A1(_04397_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04571_ ), .A4(_04398_ ), .ZN(_04970_ ) );
NAND4_X1 _12743_ ( .A1(_04967_ ), .A2(_04968_ ), .A3(_04969_ ), .A4(_04970_ ), .ZN(_04971_ ) );
OAI21_X1 _12744_ ( .A(_04971_ ), .B1(_04401_ ), .B2(_04402_ ), .ZN(_04972_ ) );
NAND2_X1 _12745_ ( .A1(_04966_ ), .A2(_04972_ ), .ZN(_04973_ ) );
NAND2_X1 _12746_ ( .A1(_04973_ ), .A2(_04163_ ), .ZN(_04974_ ) );
AND2_X2 _12747_ ( .A1(_02573_ ), .A2(fanout_net_8 ), .ZN(_04975_ ) );
BUF_X2 _12748_ ( .A(_02833_ ), .Z(_04976_ ) );
OAI21_X1 _12749_ ( .A(_02829_ ), .B1(_02826_ ), .B2(_02827_ ), .ZN(_04977_ ) );
NAND2_X1 _12750_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_04978_ ) );
NAND2_X1 _12751_ ( .A1(_04977_ ), .A2(_04978_ ), .ZN(_04979_ ) );
XNOR2_X1 _12752_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_04980_ ) );
XOR2_X1 _12753_ ( .A(_04979_ ), .B(_04980_ ), .Z(_04981_ ) );
AOI211_X1 _12754_ ( .A(_02840_ ), .B(_04975_ ), .C1(_04976_ ), .C2(_04981_ ), .ZN(_04982_ ) );
NAND2_X1 _12755_ ( .A1(_04973_ ), .A2(\ID_EX_typ [3] ), .ZN(_04983_ ) );
INV_X1 _12756_ ( .A(\ID_EX_pc [30] ), .ZN(_04984_ ) );
NOR2_X1 _12757_ ( .A1(_02857_ ), .A2(_04984_ ), .ZN(_04985_ ) );
XNOR2_X1 _12758_ ( .A(_04985_ ), .B(\ID_EX_pc [31] ), .ZN(_04986_ ) );
MUX2_X1 _12759_ ( .A(_04986_ ), .B(_04981_ ), .S(_04084_ ), .Z(_04987_ ) );
OAI21_X1 _12760_ ( .A(_04983_ ), .B1(_04987_ ), .B2(\ID_EX_typ [3] ), .ZN(_04988_ ) );
AOI21_X1 _12761_ ( .A(_04982_ ), .B1(_04988_ ), .B2(_01655_ ), .ZN(_04989_ ) );
OAI211_X1 _12762_ ( .A(_01329_ ), .B(_04974_ ), .C1(_04989_ ), .C2(_04163_ ), .ZN(_00151_ ) );
INV_X1 _12763_ ( .A(\ID_EX_pc [31] ), .ZN(_04990_ ) );
NOR2_X1 _12764_ ( .A1(_04990_ ), .A2(fanout_net_3 ), .ZN(_00152_ ) );
NOR2_X1 _12765_ ( .A1(_04984_ ), .A2(fanout_net_3 ), .ZN(_00153_ ) );
NOR2_X1 _12766_ ( .A1(_04946_ ), .A2(fanout_net_3 ), .ZN(_00154_ ) );
NOR2_X1 _12767_ ( .A1(_04944_ ), .A2(fanout_net_3 ), .ZN(_00155_ ) );
AND2_X1 _12768_ ( .A1(_01329_ ), .A2(\ID_EX_pc [19] ), .ZN(_00156_ ) );
NOR2_X1 _12769_ ( .A1(_04241_ ), .A2(fanout_net_3 ), .ZN(_00157_ ) );
AND2_X1 _12770_ ( .A1(_01246_ ), .A2(\ID_EX_pc [17] ), .ZN(_00158_ ) );
NOR2_X1 _12771_ ( .A1(_04272_ ), .A2(fanout_net_3 ), .ZN(_00159_ ) );
INV_X1 _12772_ ( .A(\ID_EX_pc [15] ), .ZN(_04991_ ) );
NOR2_X1 _12773_ ( .A1(_04991_ ), .A2(fanout_net_3 ), .ZN(_00160_ ) );
NOR2_X1 _12774_ ( .A1(_04347_ ), .A2(fanout_net_3 ), .ZN(_00161_ ) );
NOR2_X1 _12775_ ( .A1(_04374_ ), .A2(fanout_net_3 ), .ZN(_00162_ ) );
NOR2_X1 _12776_ ( .A1(_04372_ ), .A2(fanout_net_3 ), .ZN(_00163_ ) );
NOR2_X1 _12777_ ( .A1(_02825_ ), .A2(fanout_net_3 ), .ZN(_00164_ ) );
NOR2_X1 _12778_ ( .A1(_04442_ ), .A2(fanout_net_3 ), .ZN(_00165_ ) );
NOR2_X1 _12779_ ( .A1(_04500_ ), .A2(fanout_net_3 ), .ZN(_00166_ ) );
AND2_X1 _12780_ ( .A1(_01246_ ), .A2(\ID_EX_pc [9] ), .ZN(_00167_ ) );
NOR2_X1 _12781_ ( .A1(_04553_ ), .A2(fanout_net_3 ), .ZN(_00168_ ) );
NOR2_X1 _12782_ ( .A1(_04575_ ), .A2(fanout_net_3 ), .ZN(_00169_ ) );
NOR2_X1 _12783_ ( .A1(_04618_ ), .A2(fanout_net_3 ), .ZN(_00170_ ) );
AND2_X1 _12784_ ( .A1(_01246_ ), .A2(\ID_EX_pc [5] ), .ZN(_00171_ ) );
NOR2_X1 _12785_ ( .A1(_04672_ ), .A2(fanout_net_3 ), .ZN(_00172_ ) );
AND2_X1 _12786_ ( .A1(_01246_ ), .A2(\ID_EX_pc [3] ), .ZN(_00173_ ) );
INV_X1 _12787_ ( .A(\ID_EX_pc [2] ), .ZN(_04992_ ) );
NOR2_X1 _12788_ ( .A1(_04992_ ), .A2(fanout_net_3 ), .ZN(_00174_ ) );
NOR2_X1 _12789_ ( .A1(_04472_ ), .A2(fanout_net_3 ), .ZN(_00175_ ) );
INV_X1 _12790_ ( .A(\ID_EX_pc [1] ), .ZN(_04993_ ) );
NOR2_X1 _12791_ ( .A1(_04993_ ), .A2(fanout_net_3 ), .ZN(_00176_ ) );
NOR2_X1 _12792_ ( .A1(_04800_ ), .A2(fanout_net_3 ), .ZN(_00177_ ) );
NOR2_X1 _12793_ ( .A1(_04153_ ), .A2(fanout_net_3 ), .ZN(_00178_ ) );
NOR2_X1 _12794_ ( .A1(_04154_ ), .A2(fanout_net_3 ), .ZN(_00179_ ) );
NOR2_X1 _12795_ ( .A1(_04854_ ), .A2(fanout_net_3 ), .ZN(_00180_ ) );
NOR2_X1 _12796_ ( .A1(_04852_ ), .A2(fanout_net_4 ), .ZN(_00181_ ) );
AND2_X1 _12797_ ( .A1(_01246_ ), .A2(\ID_EX_pc [23] ), .ZN(_00182_ ) );
AND2_X1 _12798_ ( .A1(_01246_ ), .A2(\ID_EX_pc [22] ), .ZN(_00183_ ) );
NOR2_X1 _12799_ ( .A1(_01656_ ), .A2(fanout_net_4 ), .ZN(_00184_ ) );
AND2_X1 _12800_ ( .A1(_01586_ ), .A2(_01620_ ), .ZN(_04994_ ) );
MUX2_X1 _12801_ ( .A(io_master_arready ), .B(_01630_ ), .S(_04994_ ), .Z(_04995_ ) );
AND2_X2 _12802_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_04996_ ) );
AND2_X1 _12803_ ( .A1(_04996_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_04997_ ) );
AND3_X1 _12804_ ( .A1(_04995_ ), .A2(_04997_ ), .A3(_01623_ ), .ZN(_04998_ ) );
NOR2_X1 _12805_ ( .A1(_01674_ ), .A2(\EX_LS_flag [2] ), .ZN(_04999_ ) );
INV_X1 _12806_ ( .A(io_master_awready ), .ZN(_05000_ ) );
AOI22_X1 _12807_ ( .A1(_04999_ ), .A2(_05000_ ), .B1(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .B2(_04996_ ), .ZN(_05001_ ) );
NOR2_X1 _12808_ ( .A1(_04998_ ), .A2(_05001_ ), .ZN(_05002_ ) );
INV_X1 _12809_ ( .A(\mylsu.state [0] ), .ZN(_05003_ ) );
INV_X1 _12810_ ( .A(\mylsu.state [4] ), .ZN(_05004_ ) );
AOI21_X1 _12811_ ( .A(_05002_ ), .B1(_05003_ ), .B2(_05004_ ), .ZN(_05005_ ) );
NOR2_X1 _12812_ ( .A1(_01543_ ), .A2(fanout_net_4 ), .ZN(_05006_ ) );
INV_X1 _12813_ ( .A(_05006_ ), .ZN(_05007_ ) );
OAI22_X1 _12814_ ( .A1(_05005_ ), .A2(_05007_ ), .B1(fanout_net_4 ), .B2(_01645_ ), .ZN(_00185_ ) );
NOR2_X1 _12815_ ( .A1(_01659_ ), .A2(fanout_net_4 ), .ZN(_00186_ ) );
NOR2_X1 _12816_ ( .A1(_01647_ ), .A2(fanout_net_4 ), .ZN(_00187_ ) );
NOR2_X1 _12817_ ( .A1(_03728_ ), .A2(fanout_net_4 ), .ZN(_00188_ ) );
NOR2_X1 _12818_ ( .A1(_04159_ ), .A2(fanout_net_4 ), .ZN(_00189_ ) );
BUF_X4 _12819_ ( .A(_03982_ ), .Z(_05008_ ) );
NOR2_X1 _12820_ ( .A1(_05008_ ), .A2(fanout_net_4 ), .ZN(_00190_ ) );
NOR2_X1 _12821_ ( .A1(_04073_ ), .A2(fanout_net_4 ), .ZN(_00191_ ) );
BUF_X2 _12822_ ( .A(_04227_ ), .Z(_05009_ ) );
NOR2_X1 _12823_ ( .A1(_05009_ ), .A2(fanout_net_4 ), .ZN(_00192_ ) );
INV_X32 _12824_ ( .A(\IF_ID_inst [3] ), .ZN(_05010_ ) );
NAND3_X1 _12825_ ( .A1(_05010_ ), .A2(\IF_ID_inst [1] ), .A3(\IF_ID_inst [0] ), .ZN(_05011_ ) );
NOR2_X1 _12826_ ( .A1(_05011_ ), .A2(\IF_ID_inst [2] ), .ZN(_05012_ ) );
INV_X1 _12827_ ( .A(\IF_ID_inst [12] ), .ZN(_05013_ ) );
AND4_X1 _12828_ ( .A1(\IF_ID_inst [4] ), .A2(_05013_ ), .A3(\IF_ID_inst [5] ), .A4(\IF_ID_inst [6] ), .ZN(_05014_ ) );
AND2_X1 _12829_ ( .A1(_05012_ ), .A2(_05014_ ), .ZN(_05015_ ) );
NAND2_X2 _12830_ ( .A1(_05015_ ), .A2(\IF_ID_inst [13] ), .ZN(_05016_ ) );
AND4_X1 _12831_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [6] ), .A4(\IF_ID_inst [12] ), .ZN(_05017_ ) );
AND2_X1 _12832_ ( .A1(_05012_ ), .A2(_05017_ ), .ZN(_05018_ ) );
INV_X1 _12833_ ( .A(_05018_ ), .ZN(_05019_ ) );
AOI211_X1 _12834_ ( .A(fanout_net_4 ), .B(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .C1(_05016_ ), .C2(_05019_ ), .ZN(_00193_ ) );
AOI211_X1 _12835_ ( .A(fanout_net_4 ), .B(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .C1(_05016_ ), .C2(_05019_ ), .ZN(_00194_ ) );
INV_X1 _12836_ ( .A(\IF_ID_inst [21] ), .ZN(_05020_ ) );
AOI211_X1 _12837_ ( .A(fanout_net_4 ), .B(_05020_ ), .C1(_05016_ ), .C2(_05019_ ), .ZN(_00195_ ) );
AND2_X1 _12838_ ( .A1(_05016_ ), .A2(_05019_ ), .ZN(_05021_ ) );
INV_X1 _12839_ ( .A(_05021_ ), .ZN(_05022_ ) );
BUF_X2 _12840_ ( .A(_05022_ ), .Z(_05023_ ) );
INV_X1 _12841_ ( .A(\IF_ID_inst [20] ), .ZN(_05024_ ) );
AOI21_X1 _12842_ ( .A(fanout_net_4 ), .B1(_05023_ ), .B2(_05024_ ), .ZN(_00196_ ) );
INV_X1 _12843_ ( .A(\IF_ID_inst [29] ), .ZN(_05025_ ) );
AOI21_X1 _12844_ ( .A(fanout_net_4 ), .B1(_05023_ ), .B2(_05025_ ), .ZN(_00197_ ) );
INV_X1 _12845_ ( .A(\IF_ID_inst [28] ), .ZN(_05026_ ) );
AOI21_X1 _12846_ ( .A(fanout_net_4 ), .B1(_05023_ ), .B2(_05026_ ), .ZN(_00198_ ) );
AOI211_X1 _12847_ ( .A(fanout_net_4 ), .B(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C1(_05016_ ), .C2(_05019_ ), .ZN(_00199_ ) );
NAND3_X1 _12848_ ( .A1(_05023_ ), .A2(_01052_ ), .A3(\IF_ID_inst [26] ), .ZN(_05027_ ) );
NOR4_X1 _12849_ ( .A1(\IF_ID_inst [10] ), .A2(\IF_ID_inst [9] ), .A3(\IF_ID_inst [8] ), .A4(\IF_ID_inst [7] ), .ZN(_05028_ ) );
INV_X1 _12850_ ( .A(\IF_ID_inst [11] ), .ZN(_05029_ ) );
INV_X1 _12851_ ( .A(\IF_ID_inst [15] ), .ZN(_05030_ ) );
NAND3_X1 _12852_ ( .A1(_05028_ ), .A2(_05029_ ), .A3(_05030_ ), .ZN(_05031_ ) );
NOR2_X1 _12853_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_05032_ ) );
CLKBUF_X2 _12854_ ( .A(_05032_ ), .Z(_05033_ ) );
INV_X1 _12855_ ( .A(_05033_ ), .ZN(_05034_ ) );
NOR2_X1 _12856_ ( .A1(_05031_ ), .A2(_05034_ ), .ZN(_05035_ ) );
NOR4_X1 _12857_ ( .A1(\IF_ID_inst [31] ), .A2(\IF_ID_inst [30] ), .A3(\IF_ID_inst [29] ), .A4(\IF_ID_inst [28] ), .ZN(_05036_ ) );
NOR2_X1 _12858_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_05037_ ) );
NOR2_X1 _12859_ ( .A1(\IF_ID_inst [24] ), .A2(\IF_ID_inst [27] ), .ZN(_05038_ ) );
AND2_X1 _12860_ ( .A1(_05037_ ), .A2(_05038_ ), .ZN(_05039_ ) );
AND2_X1 _12861_ ( .A1(_05036_ ), .A2(_05039_ ), .ZN(_05040_ ) );
AND3_X1 _12862_ ( .A1(_05035_ ), .A2(_05015_ ), .A3(_05040_ ), .ZN(_05041_ ) );
NOR2_X1 _12863_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_05042_ ) );
NOR2_X1 _12864_ ( .A1(\IF_ID_inst [18] ), .A2(\IF_ID_inst [19] ), .ZN(_05043_ ) );
NOR2_X1 _12865_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_05044_ ) );
AND3_X1 _12866_ ( .A1(_05042_ ), .A2(_05043_ ), .A3(_05044_ ), .ZN(_05045_ ) );
AND3_X1 _12867_ ( .A1(_05045_ ), .A2(_05020_ ), .A3(_05024_ ), .ZN(_05046_ ) );
AND2_X1 _12868_ ( .A1(_05041_ ), .A2(_05046_ ), .ZN(_05047_ ) );
OR2_X1 _12869_ ( .A1(_05047_ ), .A2(_05023_ ), .ZN(_05048_ ) );
OAI21_X1 _12870_ ( .A(_05027_ ), .B1(_05048_ ), .B2(fanout_net_4 ), .ZN(_00200_ ) );
AOI211_X1 _12871_ ( .A(fanout_net_4 ), .B(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .C1(_05016_ ), .C2(_05019_ ), .ZN(_00201_ ) );
INV_X1 _12872_ ( .A(\IF_ID_inst [24] ), .ZN(_05049_ ) );
AOI211_X1 _12873_ ( .A(fanout_net_4 ), .B(_05049_ ), .C1(_05016_ ), .C2(_05019_ ), .ZN(_00202_ ) );
INV_X1 _12874_ ( .A(\IF_ID_inst [23] ), .ZN(_05050_ ) );
AOI211_X1 _12875_ ( .A(fanout_net_4 ), .B(_05050_ ), .C1(_05016_ ), .C2(_05019_ ), .ZN(_00203_ ) );
AOI22_X1 _12876_ ( .A1(_05023_ ), .A2(\IF_ID_inst [22] ), .B1(_05046_ ), .B2(_05041_ ), .ZN(_05051_ ) );
NOR2_X1 _12877_ ( .A1(_05051_ ), .A2(fanout_net_4 ), .ZN(_00204_ ) );
AND2_X1 _12878_ ( .A1(_01246_ ), .A2(\myidu.state [2] ), .ZN(_00205_ ) );
CLKBUF_X2 _12879_ ( .A(_05012_ ), .Z(_05052_ ) );
AND2_X2 _12880_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05053_ ) );
INV_X1 _12881_ ( .A(\IF_ID_inst [6] ), .ZN(_05054_ ) );
NOR2_X1 _12882_ ( .A1(_05054_ ), .A2(\IF_ID_inst [12] ), .ZN(_05055_ ) );
AND3_X1 _12883_ ( .A1(_05052_ ), .A2(_05053_ ), .A3(_05055_ ), .ZN(_05056_ ) );
NOR2_X1 _12884_ ( .A1(_05024_ ), .A2(\IF_ID_inst [21] ), .ZN(_05057_ ) );
AND4_X1 _12885_ ( .A1(_05056_ ), .A2(_05035_ ), .A3(_05040_ ), .A4(_05057_ ), .ZN(_05058_ ) );
AND2_X1 _12886_ ( .A1(_05058_ ), .A2(_05045_ ), .ZN(_05059_ ) );
AND3_X1 _12887_ ( .A1(_05035_ ), .A2(_05056_ ), .A3(_05046_ ), .ZN(_05060_ ) );
AND2_X1 _12888_ ( .A1(_05060_ ), .A2(_05040_ ), .ZN(_05061_ ) );
NOR2_X1 _12889_ ( .A1(\IF_ID_inst [31] ), .A2(\IF_ID_inst [30] ), .ZN(_05062_ ) );
AND2_X1 _12890_ ( .A1(_05042_ ), .A2(_05043_ ), .ZN(_05063_ ) );
AND4_X1 _12891_ ( .A1(\IF_ID_inst [21] ), .A2(_05024_ ), .A3(\IF_ID_inst [29] ), .A4(\IF_ID_inst [28] ), .ZN(_05064_ ) );
AND4_X1 _12892_ ( .A1(_05062_ ), .A2(_05063_ ), .A3(_05064_ ), .A4(_05044_ ), .ZN(_05065_ ) );
AND3_X1 _12893_ ( .A1(_05035_ ), .A2(_05056_ ), .A3(_05065_ ), .ZN(_05066_ ) );
AND2_X1 _12894_ ( .A1(_05066_ ), .A2(_05039_ ), .ZN(_05067_ ) );
NOR3_X1 _12895_ ( .A1(_05059_ ), .A2(_05061_ ), .A3(_05067_ ), .ZN(_05068_ ) );
INV_X1 _12896_ ( .A(\IF_ID_inst [4] ), .ZN(_05069_ ) );
AND2_X1 _12897_ ( .A1(_05069_ ), .A2(\IF_ID_inst [5] ), .ZN(_05070_ ) );
NOR2_X1 _12898_ ( .A1(\IF_ID_inst [6] ), .A2(\IF_ID_inst [12] ), .ZN(_05071_ ) );
AND3_X1 _12899_ ( .A1(_05052_ ), .A2(_05070_ ), .A3(_05071_ ), .ZN(_05072_ ) );
INV_X1 _12900_ ( .A(\IF_ID_inst [13] ), .ZN(_05073_ ) );
NOR2_X1 _12901_ ( .A1(_05073_ ), .A2(\IF_ID_inst [14] ), .ZN(_05074_ ) );
AND2_X1 _12902_ ( .A1(_05072_ ), .A2(_05074_ ), .ZN(_05075_ ) );
INV_X1 _12903_ ( .A(_05075_ ), .ZN(_05076_ ) );
AND2_X2 _12904_ ( .A1(_05070_ ), .A2(\IF_ID_inst [6] ), .ZN(_05077_ ) );
AND2_X4 _12905_ ( .A1(_05077_ ), .A2(_05012_ ), .ZN(_05078_ ) );
INV_X1 _12906_ ( .A(_05074_ ), .ZN(_05079_ ) );
AND2_X1 _12907_ ( .A1(_05078_ ), .A2(_05079_ ), .ZN(_05080_ ) );
INV_X1 _12908_ ( .A(_05080_ ), .ZN(_05081_ ) );
AND3_X1 _12909_ ( .A1(\IF_ID_inst [1] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [2] ), .ZN(_05082_ ) );
AND3_X1 _12910_ ( .A1(_05082_ ), .A2(\IF_ID_inst [3] ), .A3(_05033_ ), .ZN(_05083_ ) );
NOR2_X1 _12911_ ( .A1(_05013_ ), .A2(\IF_ID_inst [6] ), .ZN(_05084_ ) );
NOR2_X1 _12912_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05085_ ) );
AND2_X1 _12913_ ( .A1(_05084_ ), .A2(_05085_ ), .ZN(_05086_ ) );
AND2_X1 _12914_ ( .A1(_05083_ ), .A2(_05086_ ), .ZN(_05087_ ) );
INV_X1 _12915_ ( .A(_05087_ ), .ZN(_05088_ ) );
NAND4_X1 _12916_ ( .A1(_05084_ ), .A2(_05069_ ), .A3(\IF_ID_inst [5] ), .A4(_05033_ ), .ZN(_05089_ ) );
NOR3_X1 _12917_ ( .A1(_05089_ ), .A2(\IF_ID_inst [2] ), .A3(_05011_ ), .ZN(_05090_ ) );
AOI21_X1 _12918_ ( .A(_05090_ ), .B1(_05033_ ), .B2(_05072_ ), .ZN(_05091_ ) );
AND4_X1 _12919_ ( .A1(_05076_ ), .A2(_05081_ ), .A3(_05088_ ), .A4(_05091_ ), .ZN(_05092_ ) );
AND4_X1 _12920_ ( .A1(_01242_ ), .A2(_05068_ ), .A3(\IF_ID_inst [11] ), .A4(_05092_ ), .ZN(_00206_ ) );
AND4_X1 _12921_ ( .A1(_01242_ ), .A2(_05068_ ), .A3(\IF_ID_inst [10] ), .A4(_05092_ ), .ZN(_00207_ ) );
AND4_X1 _12922_ ( .A1(_01052_ ), .A2(_05068_ ), .A3(\IF_ID_inst [9] ), .A4(_05092_ ), .ZN(_00208_ ) );
AND4_X1 _12923_ ( .A1(_01052_ ), .A2(_05068_ ), .A3(\IF_ID_inst [8] ), .A4(_05092_ ), .ZN(_00209_ ) );
AND4_X1 _12924_ ( .A1(_01052_ ), .A2(_05068_ ), .A3(\IF_ID_inst [7] ), .A4(_05092_ ), .ZN(_00210_ ) );
INV_X1 _12925_ ( .A(\IF_ID_inst [7] ), .ZN(_05093_ ) );
AND4_X1 _12926_ ( .A1(_05093_ ), .A2(_05052_ ), .A3(\IF_ID_inst [6] ), .A4(_05053_ ), .ZN(_05094_ ) );
NOR4_X1 _12927_ ( .A1(\IF_ID_inst [15] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [14] ), .A4(\IF_ID_inst [12] ), .ZN(_05095_ ) );
NOR4_X1 _12928_ ( .A1(\IF_ID_inst [10] ), .A2(\IF_ID_inst [9] ), .A3(\IF_ID_inst [8] ), .A4(\IF_ID_inst [11] ), .ZN(_05096_ ) );
AND3_X1 _12929_ ( .A1(_05094_ ), .A2(_05095_ ), .A3(_05096_ ), .ZN(_05097_ ) );
AND4_X1 _12930_ ( .A1(_05040_ ), .A2(_05063_ ), .A3(_05044_ ), .A4(_05057_ ), .ZN(_05098_ ) );
NAND4_X1 _12931_ ( .A1(_05039_ ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .A4(_05062_ ), .ZN(_05099_ ) );
NAND4_X1 _12932_ ( .A1(_05063_ ), .A2(\IF_ID_inst [21] ), .A3(_05024_ ), .A4(_05044_ ), .ZN(_05100_ ) );
NOR2_X1 _12933_ ( .A1(_05099_ ), .A2(_05100_ ), .ZN(_05101_ ) );
OAI21_X1 _12934_ ( .A(_05097_ ), .B1(_05098_ ), .B2(_05101_ ), .ZN(_05102_ ) );
AND2_X1 _12935_ ( .A1(_05046_ ), .A2(_05040_ ), .ZN(_05103_ ) );
NAND2_X1 _12936_ ( .A1(_05097_ ), .A2(_05103_ ), .ZN(_05104_ ) );
NAND2_X1 _12937_ ( .A1(_05102_ ), .A2(_05104_ ), .ZN(_05105_ ) );
INV_X1 _12938_ ( .A(\IF_ID_inst [19] ), .ZN(_05106_ ) );
AND2_X1 _12939_ ( .A1(_05082_ ), .A2(\IF_ID_inst [3] ), .ZN(_05107_ ) );
AND2_X1 _12940_ ( .A1(_05077_ ), .A2(_05107_ ), .ZN(_05108_ ) );
BUF_X2 _12941_ ( .A(_05108_ ), .Z(_05109_ ) );
INV_X1 _12942_ ( .A(_05109_ ), .ZN(_05110_ ) );
AND4_X1 _12943_ ( .A1(_05054_ ), .A2(_05033_ ), .A3(_05085_ ), .A4(\IF_ID_inst [12] ), .ZN(_05111_ ) );
BUF_X2 _12944_ ( .A(_05107_ ), .Z(_05112_ ) );
AND2_X1 _12945_ ( .A1(_05111_ ), .A2(_05112_ ), .ZN(_05113_ ) );
INV_X1 _12946_ ( .A(_05113_ ), .ZN(_05114_ ) );
AND2_X1 _12947_ ( .A1(_05082_ ), .A2(_05010_ ), .ZN(_05115_ ) );
NOR2_X1 _12948_ ( .A1(_05069_ ), .A2(\IF_ID_inst [6] ), .ZN(_05116_ ) );
AND2_X1 _12949_ ( .A1(_05115_ ), .A2(_05116_ ), .ZN(_05117_ ) );
INV_X1 _12950_ ( .A(_05117_ ), .ZN(_05118_ ) );
NAND3_X1 _12951_ ( .A1(_05110_ ), .A2(_05114_ ), .A3(_05118_ ), .ZN(_05119_ ) );
NOR4_X1 _12952_ ( .A1(_05105_ ), .A2(fanout_net_4 ), .A3(_05106_ ), .A4(_05119_ ), .ZN(_00211_ ) );
INV_X1 _12953_ ( .A(\IF_ID_inst [18] ), .ZN(_05120_ ) );
NOR4_X1 _12954_ ( .A1(_05105_ ), .A2(fanout_net_4 ), .A3(_05120_ ), .A4(_05119_ ), .ZN(_00212_ ) );
INV_X1 _12955_ ( .A(\IF_ID_inst [17] ), .ZN(_05121_ ) );
NOR4_X1 _12956_ ( .A1(_05105_ ), .A2(fanout_net_4 ), .A3(_05121_ ), .A4(_05119_ ), .ZN(_00213_ ) );
NOR2_X1 _12957_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .ZN(_05122_ ) );
NOR2_X1 _12958_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_05123_ ) );
AND3_X1 _12959_ ( .A1(_05122_ ), .A2(_05123_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05124_ ) );
AND2_X1 _12960_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_05125_ ) );
AND3_X1 _12961_ ( .A1(_05124_ ), .A2(_05125_ ), .A3(_05037_ ), .ZN(_05126_ ) );
AND2_X2 _12962_ ( .A1(_05012_ ), .A2(_05071_ ), .ZN(_05127_ ) );
AND3_X1 _12963_ ( .A1(_05126_ ), .A2(_05053_ ), .A3(_05127_ ), .ZN(_05128_ ) );
INV_X1 _12964_ ( .A(_05128_ ), .ZN(_05129_ ) );
INV_X1 _12965_ ( .A(\IF_ID_inst [14] ), .ZN(_05130_ ) );
NOR2_X1 _12966_ ( .A1(_05130_ ), .A2(\IF_ID_inst [13] ), .ZN(_05131_ ) );
AND2_X1 _12967_ ( .A1(_05131_ ), .A2(_05037_ ), .ZN(_05132_ ) );
AND2_X1 _12968_ ( .A1(_05132_ ), .A2(_05124_ ), .ZN(_05133_ ) );
AND2_X1 _12969_ ( .A1(_05032_ ), .A2(_05037_ ), .ZN(_05134_ ) );
AND2_X1 _12970_ ( .A1(_05124_ ), .A2(_05134_ ), .ZN(_05135_ ) );
OAI211_X1 _12971_ ( .A(_05053_ ), .B(_05127_ ), .C1(_05133_ ), .C2(_05135_ ), .ZN(_05136_ ) );
AND2_X1 _12972_ ( .A1(_05012_ ), .A2(_05084_ ), .ZN(_05137_ ) );
AND2_X1 _12973_ ( .A1(_05137_ ), .A2(_05053_ ), .ZN(_05138_ ) );
INV_X1 _12974_ ( .A(_05138_ ), .ZN(_05139_ ) );
OAI211_X1 _12975_ ( .A(_05124_ ), .B(_05037_ ), .C1(_05073_ ), .C2(_05130_ ), .ZN(_05140_ ) );
OAI211_X1 _12976_ ( .A(_05129_ ), .B(_05136_ ), .C1(_05139_ ), .C2(_05140_ ), .ZN(_05141_ ) );
NOR3_X1 _12977_ ( .A1(\IF_ID_inst [29] ), .A2(\IF_ID_inst [28] ), .A3(\IF_ID_inst [27] ), .ZN(_05142_ ) );
AND3_X1 _12978_ ( .A1(_05142_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\IF_ID_inst [30] ), .ZN(_05143_ ) );
AND2_X1 _12979_ ( .A1(_05143_ ), .A2(_05132_ ), .ZN(_05144_ ) );
AND2_X1 _12980_ ( .A1(_05138_ ), .A2(_05144_ ), .ZN(_05145_ ) );
AND2_X1 _12981_ ( .A1(_05138_ ), .A2(_05126_ ), .ZN(_05146_ ) );
NOR3_X1 _12982_ ( .A1(_05141_ ), .A2(_05145_ ), .A3(_05146_ ), .ZN(_05147_ ) );
NOR2_X1 _12983_ ( .A1(_05069_ ), .A2(\IF_ID_inst [5] ), .ZN(_05148_ ) );
AND2_X1 _12984_ ( .A1(_05127_ ), .A2(_05148_ ), .ZN(_05149_ ) );
AND2_X1 _12985_ ( .A1(_05149_ ), .A2(_05074_ ), .ZN(_05150_ ) );
AND2_X1 _12986_ ( .A1(_05127_ ), .A2(_05085_ ), .ZN(_05151_ ) );
AND2_X1 _12987_ ( .A1(_05151_ ), .A2(_05074_ ), .ZN(_05152_ ) );
INV_X1 _12988_ ( .A(_05152_ ), .ZN(_05153_ ) );
AND2_X1 _12989_ ( .A1(_05137_ ), .A2(_05148_ ), .ZN(_05154_ ) );
BUF_X2 _12990_ ( .A(_05154_ ), .Z(_05155_ ) );
NAND2_X1 _12991_ ( .A1(_05155_ ), .A2(_05074_ ), .ZN(_05156_ ) );
NAND2_X1 _12992_ ( .A1(_05153_ ), .A2(_05156_ ), .ZN(_05157_ ) );
AND3_X1 _12993_ ( .A1(_05070_ ), .A2(_05055_ ), .A3(_05033_ ), .ZN(_05158_ ) );
AOI211_X1 _12994_ ( .A(_05150_ ), .B(_05157_ ), .C1(_05052_ ), .C2(_05158_ ), .ZN(_05159_ ) );
AND2_X1 _12995_ ( .A1(_05149_ ), .A2(_05079_ ), .ZN(_05160_ ) );
INV_X1 _12996_ ( .A(_05160_ ), .ZN(_05161_ ) );
NAND3_X1 _12997_ ( .A1(_05144_ ), .A2(_05137_ ), .A3(_05148_ ), .ZN(_05162_ ) );
NAND4_X1 _12998_ ( .A1(_05137_ ), .A2(_05148_ ), .A3(_05124_ ), .A4(_05132_ ), .ZN(_05163_ ) );
AND3_X1 _12999_ ( .A1(_05037_ ), .A2(_05122_ ), .A3(_05123_ ), .ZN(_05164_ ) );
AND3_X1 _13000_ ( .A1(_05164_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_05074_ ), .ZN(_05165_ ) );
NAND3_X1 _13001_ ( .A1(_05165_ ), .A2(_05053_ ), .A3(_05127_ ), .ZN(_05166_ ) );
NAND4_X1 _13002_ ( .A1(_05127_ ), .A2(_05053_ ), .A3(_05134_ ), .A4(_05143_ ), .ZN(_05167_ ) );
AND4_X1 _13003_ ( .A1(_05162_ ), .A2(_05163_ ), .A3(_05166_ ), .A4(_05167_ ), .ZN(_05168_ ) );
AND2_X1 _13004_ ( .A1(_05158_ ), .A2(_05115_ ), .ZN(_05169_ ) );
CLKBUF_X2 _13005_ ( .A(_05077_ ), .Z(_05170_ ) );
AND3_X1 _13006_ ( .A1(_05170_ ), .A2(\IF_ID_inst [12] ), .A3(_05052_ ), .ZN(_05171_ ) );
AOI21_X1 _13007_ ( .A(_05169_ ), .B1(_05171_ ), .B2(_05125_ ), .ZN(_05172_ ) );
NAND2_X1 _13008_ ( .A1(_05155_ ), .A2(_05125_ ), .ZN(_05173_ ) );
AND4_X1 _13009_ ( .A1(_05161_ ), .A2(_05168_ ), .A3(_05172_ ), .A4(_05173_ ), .ZN(_05174_ ) );
AND2_X1 _13010_ ( .A1(_05078_ ), .A2(_05013_ ), .ZN(_05175_ ) );
AOI221_X4 _13011_ ( .A(_05022_ ), .B1(_05073_ ), .B2(_05171_ ), .C1(\IF_ID_inst [14] ), .C2(_05175_ ), .ZN(_05176_ ) );
AND4_X1 _13012_ ( .A1(_05147_ ), .A2(_05159_ ), .A3(_05174_ ), .A4(_05176_ ), .ZN(_05177_ ) );
NOR2_X1 _13013_ ( .A1(_05105_ ), .A2(_05119_ ), .ZN(_05178_ ) );
AND2_X1 _13014_ ( .A1(_05076_ ), .A2(_05091_ ), .ZN(_05179_ ) );
AND2_X1 _13015_ ( .A1(_05155_ ), .A2(_05135_ ), .ZN(_05180_ ) );
INV_X1 _13016_ ( .A(_05180_ ), .ZN(_05181_ ) );
NAND3_X1 _13017_ ( .A1(_05086_ ), .A2(_05073_ ), .A3(_05052_ ), .ZN(_05182_ ) );
NAND3_X1 _13018_ ( .A1(_05127_ ), .A2(_05073_ ), .A3(_05085_ ), .ZN(_05183_ ) );
AND4_X1 _13019_ ( .A1(_05179_ ), .A2(_05181_ ), .A3(_05182_ ), .A4(_05183_ ), .ZN(_05184_ ) );
AND3_X1 _13020_ ( .A1(_05177_ ), .A2(_05178_ ), .A3(_05184_ ), .ZN(_05185_ ) );
BUF_X4 _13021_ ( .A(_05185_ ), .Z(_05186_ ) );
AND2_X1 _13022_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
INV_X1 _13023_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_05187_ ) );
XNOR2_X1 _13024_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_05188_ ) );
XNOR2_X1 _13025_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_05189_ ) );
XNOR2_X1 _13026_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_05190_ ) );
XNOR2_X1 _13027_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_05191_ ) );
AND4_X1 _13028_ ( .A1(_05188_ ), .A2(_05189_ ), .A3(_05190_ ), .A4(_05191_ ), .ZN(_05192_ ) );
XNOR2_X1 _13029_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_05193_ ) );
XNOR2_X1 _13030_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_05194_ ) );
XNOR2_X1 _13031_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_05195_ ) );
XNOR2_X1 _13032_ ( .A(\IF_ID_pc [4] ), .B(\myexu.pc_jump [4] ), .ZN(_05196_ ) );
AND4_X1 _13033_ ( .A1(_05193_ ), .A2(_05194_ ), .A3(_05195_ ), .A4(_05196_ ), .ZN(_05197_ ) );
XNOR2_X1 _13034_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_05198_ ) );
XNOR2_X1 _13035_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_05199_ ) );
XNOR2_X1 _13036_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_05200_ ) );
XNOR2_X1 _13037_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_05201_ ) );
AND4_X1 _13038_ ( .A1(_05198_ ), .A2(_05199_ ), .A3(_05200_ ), .A4(_05201_ ), .ZN(_05202_ ) );
XNOR2_X1 _13039_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_05203_ ) );
XNOR2_X1 _13040_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_05204_ ) );
XNOR2_X1 _13041_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_05205_ ) );
XNOR2_X1 _13042_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_05206_ ) );
AND4_X1 _13043_ ( .A1(_05203_ ), .A2(_05204_ ), .A3(_05205_ ), .A4(_05206_ ), .ZN(_05207_ ) );
AND4_X1 _13044_ ( .A1(_05192_ ), .A2(_05197_ ), .A3(_05202_ ), .A4(_05207_ ), .ZN(_05208_ ) );
NOR2_X1 _13045_ ( .A1(_01487_ ), .A2(\myexu.pc_jump [17] ), .ZN(_05209_ ) );
AOI21_X1 _13046_ ( .A(_05209_ ), .B1(_01402_ ), .B2(\myexu.pc_jump [23] ), .ZN(_05210_ ) );
XNOR2_X1 _13047_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_05211_ ) );
INV_X1 _13048_ ( .A(\IF_ID_pc [8] ), .ZN(_05212_ ) );
AOI22_X1 _13049_ ( .A1(_01420_ ), .A2(\myexu.pc_jump [21] ), .B1(_05212_ ), .B2(\myexu.pc_jump [8] ), .ZN(_05213_ ) );
INV_X1 _13050_ ( .A(\myexu.pc_jump [21] ), .ZN(_05214_ ) );
AOI22_X1 _13051_ ( .A1(\IF_ID_pc [21] ), .A2(_05214_ ), .B1(_01487_ ), .B2(\myexu.pc_jump [17] ), .ZN(_05215_ ) );
NAND4_X1 _13052_ ( .A1(_05210_ ), .A2(_05211_ ), .A3(_05213_ ), .A4(_05215_ ), .ZN(_05216_ ) );
XNOR2_X1 _13053_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_05217_ ) );
NAND2_X1 _13054_ ( .A1(_01379_ ), .A2(\myexu.pc_jump [24] ), .ZN(_05218_ ) );
OAI211_X1 _13055_ ( .A(_05217_ ), .B(_05218_ ), .C1(_05212_ ), .C2(\myexu.pc_jump [8] ), .ZN(_05219_ ) );
INV_X1 _13056_ ( .A(\IF_ID_pc [2] ), .ZN(_05220_ ) );
NAND2_X1 _13057_ ( .A1(_05220_ ), .A2(\myexu.pc_jump [2] ), .ZN(_05221_ ) );
OAI21_X1 _13058_ ( .A(_05221_ ), .B1(_01478_ ), .B2(\myexu.pc_jump [22] ), .ZN(_05222_ ) );
NAND2_X1 _13059_ ( .A1(_01478_ ), .A2(\myexu.pc_jump [22] ), .ZN(_05223_ ) );
OAI21_X1 _13060_ ( .A(_05223_ ), .B1(_01402_ ), .B2(\myexu.pc_jump [23] ), .ZN(_05224_ ) );
NOR4_X1 _13061_ ( .A1(_05216_ ), .A2(_05219_ ), .A3(_05222_ ), .A4(_05224_ ), .ZN(_05225_ ) );
XNOR2_X1 _13062_ ( .A(\IF_ID_pc [3] ), .B(\myexu.pc_jump [3] ), .ZN(_05226_ ) );
OAI221_X1 _13063_ ( .A(_05226_ ), .B1(_01379_ ), .B2(\myexu.pc_jump [24] ), .C1(_01388_ ), .C2(\myexu.pc_jump [25] ), .ZN(_05227_ ) );
XNOR2_X1 _13064_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_05228_ ) );
XNOR2_X1 _13065_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_05229_ ) );
XNOR2_X1 _13066_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_05230_ ) );
XNOR2_X1 _13067_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_05231_ ) );
NAND4_X1 _13068_ ( .A1(_05228_ ), .A2(_05229_ ), .A3(_05230_ ), .A4(_05231_ ), .ZN(_05232_ ) );
XNOR2_X1 _13069_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_05233_ ) );
NAND2_X1 _13070_ ( .A1(_01388_ ), .A2(\myexu.pc_jump [25] ), .ZN(_05234_ ) );
OAI211_X1 _13071_ ( .A(_05233_ ), .B(_05234_ ), .C1(\myexu.pc_jump [2] ), .C2(_05220_ ), .ZN(_05235_ ) );
NOR3_X1 _13072_ ( .A1(_05227_ ), .A2(_05232_ ), .A3(_05235_ ), .ZN(_05236_ ) );
AND3_X1 _13073_ ( .A1(_05208_ ), .A2(_05225_ ), .A3(_05236_ ), .ZN(_05237_ ) );
INV_X1 _13074_ ( .A(_05237_ ), .ZN(_05238_ ) );
AOI21_X1 _13075_ ( .A(_05187_ ), .B1(_05238_ ), .B2(check_quest ), .ZN(_05239_ ) );
INV_X1 _13076_ ( .A(_05239_ ), .ZN(_05240_ ) );
BUF_X4 _13077_ ( .A(_05240_ ), .Z(_05241_ ) );
OAI21_X1 _13078_ ( .A(\ID_EX_rs1 [3] ), .B1(_05186_ ), .B2(_05241_ ), .ZN(_05242_ ) );
NAND2_X1 _13079_ ( .A1(_05177_ ), .A2(_05184_ ), .ZN(_05243_ ) );
NAND4_X1 _13080_ ( .A1(_05243_ ), .A2(\IF_ID_inst [18] ), .A3(_05178_ ), .A4(_05239_ ), .ZN(_05244_ ) );
AOI21_X1 _13081_ ( .A(fanout_net_4 ), .B1(_05242_ ), .B2(_05244_ ), .ZN(_00214_ ) );
INV_X1 _13082_ ( .A(\IF_ID_inst [16] ), .ZN(_05245_ ) );
NOR4_X1 _13083_ ( .A1(_05105_ ), .A2(fanout_net_4 ), .A3(_05245_ ), .A4(_05119_ ), .ZN(_00215_ ) );
OAI21_X1 _13084_ ( .A(\ID_EX_rs1 [2] ), .B1(_05186_ ), .B2(_05241_ ), .ZN(_05246_ ) );
NAND4_X1 _13085_ ( .A1(_05243_ ), .A2(\IF_ID_inst [17] ), .A3(_05178_ ), .A4(_05239_ ), .ZN(_05247_ ) );
AOI21_X1 _13086_ ( .A(fanout_net_4 ), .B1(_05246_ ), .B2(_05247_ ), .ZN(_00216_ ) );
NOR4_X1 _13087_ ( .A1(_05105_ ), .A2(fanout_net_4 ), .A3(_05030_ ), .A4(_05119_ ), .ZN(_00217_ ) );
OAI21_X1 _13088_ ( .A(\ID_EX_rs1 [1] ), .B1(_05186_ ), .B2(_05241_ ), .ZN(_05248_ ) );
NAND4_X1 _13089_ ( .A1(_05243_ ), .A2(\IF_ID_inst [16] ), .A3(_05178_ ), .A4(_05239_ ), .ZN(_05249_ ) );
AOI21_X1 _13090_ ( .A(fanout_net_5 ), .B1(_05248_ ), .B2(_05249_ ), .ZN(_00218_ ) );
NAND3_X1 _13091_ ( .A1(_05041_ ), .A2(_05045_ ), .A3(_05057_ ), .ZN(_05250_ ) );
NAND2_X1 _13092_ ( .A1(_05250_ ), .A2(_05088_ ), .ZN(_05251_ ) );
AND3_X1 _13093_ ( .A1(_05064_ ), .A2(_05062_ ), .A3(_05044_ ), .ZN(_05252_ ) );
AND3_X1 _13094_ ( .A1(_05252_ ), .A2(_05039_ ), .A3(_05063_ ), .ZN(_05253_ ) );
AND3_X1 _13095_ ( .A1(_05253_ ), .A2(_05015_ ), .A3(_05035_ ), .ZN(_05254_ ) );
NOR3_X1 _13096_ ( .A1(_05251_ ), .A2(_05047_ ), .A3(_05254_ ), .ZN(_05255_ ) );
AOI211_X1 _13097_ ( .A(_05018_ ), .B(_05109_ ), .C1(_05155_ ), .C2(\IF_ID_inst [13] ), .ZN(_05256_ ) );
NAND4_X1 _13098_ ( .A1(_05255_ ), .A2(_05016_ ), .A3(_05161_ ), .A4(_05256_ ), .ZN(_05257_ ) );
AOI21_X1 _13099_ ( .A(_05169_ ), .B1(_05151_ ), .B2(_05074_ ), .ZN(_05258_ ) );
AND2_X1 _13100_ ( .A1(_05086_ ), .A2(_05052_ ), .ZN(_05259_ ) );
AOI21_X1 _13101_ ( .A(_05259_ ), .B1(_05127_ ), .B2(_05085_ ), .ZN(_05260_ ) );
OAI21_X1 _13102_ ( .A(_05258_ ), .B1(\IF_ID_inst [13] ), .B2(_05260_ ), .ZN(_05261_ ) );
INV_X1 _13103_ ( .A(_05155_ ), .ZN(_05262_ ) );
NOR2_X1 _13104_ ( .A1(_05133_ ), .A2(_05135_ ), .ZN(_05263_ ) );
INV_X1 _13105_ ( .A(_05144_ ), .ZN(_05264_ ) );
AOI21_X1 _13106_ ( .A(_05262_ ), .B1(_05263_ ), .B2(_05264_ ), .ZN(_05265_ ) );
OR4_X2 _13107_ ( .A1(_05117_ ), .A2(_05261_ ), .A3(_05265_ ), .A4(_05150_ ), .ZN(_05266_ ) );
NOR4_X1 _13108_ ( .A1(_05257_ ), .A2(_05266_ ), .A3(fanout_net_5 ), .A4(_05049_ ), .ZN(_00219_ ) );
OAI21_X1 _13109_ ( .A(\ID_EX_rs1 [0] ), .B1(_05186_ ), .B2(_05241_ ), .ZN(_05267_ ) );
NAND4_X1 _13110_ ( .A1(_05243_ ), .A2(\IF_ID_inst [15] ), .A3(_05178_ ), .A4(_05239_ ), .ZN(_05268_ ) );
AOI21_X1 _13111_ ( .A(fanout_net_5 ), .B1(_05267_ ), .B2(_05268_ ), .ZN(_00220_ ) );
NOR4_X1 _13112_ ( .A1(_05257_ ), .A2(_05266_ ), .A3(fanout_net_5 ), .A4(_05050_ ), .ZN(_00221_ ) );
INV_X1 _13113_ ( .A(\IF_ID_inst [22] ), .ZN(_05269_ ) );
NOR4_X1 _13114_ ( .A1(_05257_ ), .A2(_05266_ ), .A3(fanout_net_5 ), .A4(_05269_ ), .ZN(_00222_ ) );
NOR2_X1 _13115_ ( .A1(_05185_ ), .A2(_05240_ ), .ZN(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _13116_ ( .A(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_05270_ ) );
OR4_X1 _13117_ ( .A1(_05050_ ), .A2(_05270_ ), .A3(_05257_ ), .A4(_05266_ ), .ZN(_05271_ ) );
OAI21_X1 _13118_ ( .A(\ID_EX_rs2 [3] ), .B1(_05186_ ), .B2(_05241_ ), .ZN(_05272_ ) );
AOI21_X1 _13119_ ( .A(fanout_net_5 ), .B1(_05271_ ), .B2(_05272_ ), .ZN(_00223_ ) );
NOR4_X1 _13120_ ( .A1(_05257_ ), .A2(_05266_ ), .A3(fanout_net_5 ), .A4(_05020_ ), .ZN(_00224_ ) );
NOR2_X1 _13121_ ( .A1(_05257_ ), .A2(_05266_ ), .ZN(_05273_ ) );
AOI211_X1 _13122_ ( .A(_05241_ ), .B(_05186_ ), .C1(\IF_ID_inst [22] ), .C2(_05273_ ), .ZN(_05274_ ) );
AOI211_X1 _13123_ ( .A(fanout_net_5 ), .B(_05274_ ), .C1(_02914_ ), .C2(_05270_ ), .ZN(_00225_ ) );
NOR4_X1 _13124_ ( .A1(_05257_ ), .A2(_05266_ ), .A3(fanout_net_5 ), .A4(_05024_ ), .ZN(_00226_ ) );
AOI211_X1 _13125_ ( .A(_05241_ ), .B(_05185_ ), .C1(\IF_ID_inst [21] ), .C2(_05273_ ), .ZN(_05275_ ) );
AOI211_X1 _13126_ ( .A(fanout_net_5 ), .B(_05275_ ), .C1(_03346_ ), .C2(_05270_ ), .ZN(_00227_ ) );
AND4_X1 _13127_ ( .A1(_01052_ ), .A2(_05083_ ), .A3(_01643_ ), .A4(_05086_ ), .ZN(_00228_ ) );
NOR2_X1 _13128_ ( .A1(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .A2(\ID_EX_rs2 [0] ), .ZN(_05276_ ) );
OR3_X1 _13129_ ( .A1(_05257_ ), .A2(_05266_ ), .A3(_05024_ ), .ZN(_05277_ ) );
AOI211_X1 _13130_ ( .A(fanout_net_5 ), .B(_05276_ ), .C1(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .C2(_05277_ ), .ZN(_00229_ ) );
XNOR2_X1 _13131_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_05278_ ) );
XNOR2_X1 _13132_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_05279_ ) );
XNOR2_X1 _13133_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_05280_ ) );
XNOR2_X1 _13134_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_05281_ ) );
AND4_X1 _13135_ ( .A1(_05278_ ), .A2(_05279_ ), .A3(_05280_ ), .A4(_05281_ ), .ZN(_05282_ ) );
XNOR2_X1 _13136_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_05283_ ) );
AND2_X1 _13137_ ( .A1(_05282_ ), .A2(_05283_ ), .ZN(_05284_ ) );
AND2_X1 _13138_ ( .A1(_01646_ ), .A2(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A ), .ZN(_05285_ ) );
AND2_X1 _13139_ ( .A1(_05284_ ), .A2(_05285_ ), .ZN(_05286_ ) );
XNOR2_X1 _13140_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_05287_ ) );
XNOR2_X1 _13141_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_05288_ ) );
XNOR2_X1 _13142_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_05289_ ) );
AND4_X1 _13143_ ( .A1(_05285_ ), .A2(_05287_ ), .A3(_05288_ ), .A4(_05289_ ), .ZN(_05290_ ) );
XNOR2_X1 _13144_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_05291_ ) );
XNOR2_X1 _13145_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_05292_ ) );
AND3_X1 _13146_ ( .A1(_05290_ ), .A2(_05291_ ), .A3(_05292_ ), .ZN(_05293_ ) );
NOR2_X1 _13147_ ( .A1(_05286_ ), .A2(_05293_ ), .ZN(_05294_ ) );
NOR3_X1 _13148_ ( .A1(_05105_ ), .A2(_05294_ ), .A3(_05119_ ), .ZN(_05295_ ) );
INV_X1 _13149_ ( .A(_05150_ ), .ZN(_05296_ ) );
NAND3_X1 _13150_ ( .A1(_05155_ ), .A2(\IF_ID_inst [13] ), .A3(_05130_ ), .ZN(_05297_ ) );
NAND3_X1 _13151_ ( .A1(_05155_ ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [14] ), .ZN(_05298_ ) );
NAND4_X1 _13152_ ( .A1(_05296_ ), .A2(_05161_ ), .A3(_05297_ ), .A4(_05298_ ), .ZN(_05299_ ) );
NOR2_X1 _13153_ ( .A1(_05299_ ), .A2(_05261_ ), .ZN(_05300_ ) );
AND2_X1 _13154_ ( .A1(_05300_ ), .A2(_05021_ ), .ZN(_05301_ ) );
MUX2_X1 _13155_ ( .A(_05286_ ), .B(_05295_ ), .S(_05301_ ), .Z(_05302_ ) );
AND3_X1 _13156_ ( .A1(_05302_ ), .A2(_01148_ ), .A3(IDU_ready_IFU ), .ZN(_00230_ ) );
NOR3_X1 _13157_ ( .A1(_05047_ ), .A2(_05023_ ), .A3(_05254_ ), .ZN(_05303_ ) );
NOR4_X1 _13158_ ( .A1(_05080_ ), .A2(_05087_ ), .A3(_05109_ ), .A4(_05169_ ), .ZN(_05304_ ) );
AOI21_X1 _13159_ ( .A(fanout_net_5 ), .B1(_05303_ ), .B2(_05304_ ), .ZN(_00231_ ) );
NAND2_X1 _13160_ ( .A1(_05259_ ), .A2(_05033_ ), .ZN(_05305_ ) );
NAND4_X1 _13161_ ( .A1(_05153_ ), .A2(_05076_ ), .A3(_05183_ ), .A4(_05305_ ), .ZN(_05306_ ) );
AND2_X1 _13162_ ( .A1(_05072_ ), .A2(_05033_ ), .ZN(_05307_ ) );
NOR4_X1 _13163_ ( .A1(_05048_ ), .A2(_05306_ ), .A3(_05307_ ), .A4(_05090_ ), .ZN(_05308_ ) );
NAND2_X1 _13164_ ( .A1(_05259_ ), .A2(_05131_ ), .ZN(_05309_ ) );
AOI21_X1 _13165_ ( .A(fanout_net_5 ), .B1(_05308_ ), .B2(_05309_ ), .ZN(_00232_ ) );
NOR2_X1 _13166_ ( .A1(_05141_ ), .A2(_05146_ ), .ZN(_05310_ ) );
INV_X1 _13167_ ( .A(_05310_ ), .ZN(_05311_ ) );
INV_X1 _13168_ ( .A(_05061_ ), .ZN(_05312_ ) );
AND2_X1 _13169_ ( .A1(_05166_ ), .A2(_05167_ ), .ZN(_05313_ ) );
NAND4_X1 _13170_ ( .A1(_05312_ ), .A2(_05182_ ), .A3(_05313_ ), .A4(_05183_ ), .ZN(_05314_ ) );
NAND4_X1 _13171_ ( .A1(_05070_ ), .A2(_05055_ ), .A3(_05082_ ), .A4(_05010_ ), .ZN(_05315_ ) );
OAI221_X1 _13172_ ( .A(_05110_ ), .B1(_05034_ ), .B2(_05315_ ), .C1(_05139_ ), .C2(_05264_ ), .ZN(_05316_ ) );
NOR4_X1 _13173_ ( .A1(_05311_ ), .A2(_05314_ ), .A3(_05152_ ), .A4(_05316_ ), .ZN(_05317_ ) );
INV_X1 _13174_ ( .A(_05133_ ), .ZN(_05318_ ) );
AOI21_X1 _13175_ ( .A(_05262_ ), .B1(_05264_ ), .B2(_05318_ ), .ZN(_05319_ ) );
NOR2_X1 _13176_ ( .A1(_05319_ ), .A2(_05180_ ), .ZN(_05320_ ) );
NOR2_X1 _13177_ ( .A1(_05150_ ), .A2(_05117_ ), .ZN(_05321_ ) );
NAND2_X1 _13178_ ( .A1(_05320_ ), .A2(_05321_ ), .ZN(_05322_ ) );
OAI21_X1 _13179_ ( .A(_05161_ ), .B1(_05073_ ), .B2(_05262_ ), .ZN(_05323_ ) );
NOR2_X1 _13180_ ( .A1(_05322_ ), .A2(_05323_ ), .ZN(_05324_ ) );
AOI21_X1 _13181_ ( .A(fanout_net_5 ), .B1(_05317_ ), .B2(_05324_ ), .ZN(_00233_ ) );
AOI21_X1 _13182_ ( .A(fanout_net_5 ), .B1(_05324_ ), .B2(_05088_ ), .ZN(_00234_ ) );
AND2_X1 _13183_ ( .A1(_05035_ ), .A2(_05015_ ), .ZN(_05325_ ) );
AOI21_X1 _13184_ ( .A(_05075_ ), .B1(_05325_ ), .B2(_05253_ ), .ZN(_05326_ ) );
AND2_X1 _13185_ ( .A1(_05127_ ), .A2(_05053_ ), .ZN(_05327_ ) );
AND3_X1 _13186_ ( .A1(_05124_ ), .A2(_05074_ ), .A3(_05037_ ), .ZN(_05328_ ) );
AND2_X1 _13187_ ( .A1(_05143_ ), .A2(_05134_ ), .ZN(_05329_ ) );
OAI21_X1 _13188_ ( .A(_05327_ ), .B1(_05328_ ), .B2(_05329_ ), .ZN(_05330_ ) );
AND2_X1 _13189_ ( .A1(_05326_ ), .A2(_05330_ ), .ZN(_05331_ ) );
AOI21_X1 _13190_ ( .A(fanout_net_5 ), .B1(_05331_ ), .B2(_05321_ ), .ZN(_00235_ ) );
AOI21_X1 _13191_ ( .A(_05139_ ), .B1(_05264_ ), .B2(_05140_ ), .ZN(_05332_ ) );
AND4_X1 _13192_ ( .A1(\IF_ID_inst [14] ), .A2(_05170_ ), .A3(\IF_ID_inst [12] ), .A4(_05052_ ), .ZN(_05333_ ) );
NOR3_X1 _13193_ ( .A1(_05265_ ), .A2(_05332_ ), .A3(_05333_ ), .ZN(_05334_ ) );
BUF_X2 _13194_ ( .A(_05118_ ), .Z(_05335_ ) );
NAND3_X1 _13195_ ( .A1(_05052_ ), .A2(\IF_ID_inst [13] ), .A3(_05017_ ), .ZN(_05336_ ) );
AND4_X1 _13196_ ( .A1(_05076_ ), .A2(_05334_ ), .A3(_05335_ ), .A4(_05336_ ), .ZN(_05337_ ) );
OAI21_X1 _13197_ ( .A(_05074_ ), .B1(_05151_ ), .B2(_05155_ ), .ZN(_05338_ ) );
AOI21_X1 _13198_ ( .A(fanout_net_5 ), .B1(_05337_ ), .B2(_05338_ ), .ZN(_00236_ ) );
AND2_X1 _13199_ ( .A1(_05327_ ), .A2(_05133_ ), .ZN(_05339_ ) );
OR2_X1 _13200_ ( .A1(_05339_ ), .A2(_05075_ ), .ZN(_05340_ ) );
AOI211_X1 _13201_ ( .A(_05128_ ), .B(_05340_ ), .C1(\IF_ID_inst [14] ), .C2(_05149_ ), .ZN(_05341_ ) );
AOI22_X1 _13202_ ( .A1(_05262_ ), .A2(_05139_ ), .B1(_05264_ ), .B2(_05318_ ), .ZN(_05342_ ) );
AND3_X1 _13203_ ( .A1(_05137_ ), .A2(_05033_ ), .A3(_05070_ ), .ZN(_05343_ ) );
INV_X1 _13204_ ( .A(_05343_ ), .ZN(_05344_ ) );
NAND3_X1 _13205_ ( .A1(_05078_ ), .A2(\IF_ID_inst [14] ), .A3(_05013_ ), .ZN(_05345_ ) );
NAND3_X1 _13206_ ( .A1(_05344_ ), .A2(_05016_ ), .A3(_05345_ ), .ZN(_05346_ ) );
AND3_X1 _13207_ ( .A1(_05054_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_05347_ ) );
AND2_X1 _13208_ ( .A1(_05115_ ), .A2(_05347_ ), .ZN(_05348_ ) );
NAND2_X1 _13209_ ( .A1(_05309_ ), .A2(_05305_ ), .ZN(_05349_ ) );
NOR4_X1 _13210_ ( .A1(_05342_ ), .A2(_05346_ ), .A3(_05348_ ), .A4(_05349_ ), .ZN(_05350_ ) );
AOI21_X1 _13211_ ( .A(fanout_net_5 ), .B1(_05341_ ), .B2(_05350_ ), .ZN(_00237_ ) );
NAND2_X1 _13212_ ( .A1(_05175_ ), .A2(_05125_ ), .ZN(_05351_ ) );
AOI22_X1 _13213_ ( .A1(_05327_ ), .A2(_05165_ ), .B1(_05155_ ), .B2(_05135_ ), .ZN(_05352_ ) );
OAI211_X1 _13214_ ( .A(_05053_ ), .B(_05137_ ), .C1(_05144_ ), .C2(_05135_ ), .ZN(_05353_ ) );
NAND2_X1 _13215_ ( .A1(_05352_ ), .A2(_05353_ ), .ZN(_05354_ ) );
NOR2_X1 _13216_ ( .A1(_05354_ ), .A2(_05059_ ), .ZN(_05355_ ) );
AOI22_X1 _13217_ ( .A1(_05327_ ), .A2(_05133_ ), .B1(_05138_ ), .B2(_05126_ ), .ZN(_05356_ ) );
NAND4_X1 _13218_ ( .A1(_05127_ ), .A2(_05073_ ), .A3(\IF_ID_inst [14] ), .A4(_05148_ ), .ZN(_05357_ ) );
AND4_X1 _13219_ ( .A1(_05173_ ), .A2(_05355_ ), .A3(_05356_ ), .A4(_05357_ ), .ZN(_05358_ ) );
NAND2_X1 _13220_ ( .A1(_05056_ ), .A2(_05125_ ), .ZN(_05359_ ) );
OAI21_X1 _13221_ ( .A(_05131_ ), .B1(_05151_ ), .B2(_05259_ ), .ZN(_05360_ ) );
AND4_X1 _13222_ ( .A1(_05351_ ), .A2(_05358_ ), .A3(_05359_ ), .A4(_05360_ ), .ZN(_05361_ ) );
AND4_X1 _13223_ ( .A1(\IF_ID_inst [12] ), .A2(_05170_ ), .A3(_05052_ ), .A4(_05033_ ), .ZN(_05362_ ) );
AOI21_X1 _13224_ ( .A(_05362_ ), .B1(_05155_ ), .B2(_05144_ ), .ZN(_05363_ ) );
AOI22_X1 _13225_ ( .A1(_05072_ ), .A2(_05074_ ), .B1(_05018_ ), .B2(\IF_ID_inst [14] ), .ZN(_05364_ ) );
AND4_X1 _13226_ ( .A1(_05091_ ), .A2(_05363_ ), .A3(_05172_ ), .A4(_05364_ ), .ZN(_05365_ ) );
AOI21_X1 _13227_ ( .A(fanout_net_5 ), .B1(_05361_ ), .B2(_05365_ ), .ZN(_00238_ ) );
NAND4_X1 _13228_ ( .A1(_05238_ ), .A2(_01217_ ), .A3(check_quest ), .A4(\myexu.pc_jump [0] ), .ZN(_05366_ ) );
INV_X1 _13229_ ( .A(_05366_ ), .ZN(_00242_ ) );
NOR2_X2 _13230_ ( .A1(_05237_ ), .A2(_01641_ ), .ZN(_05367_ ) );
INV_X1 _13231_ ( .A(_05367_ ), .ZN(_05368_ ) );
BUF_X4 _13232_ ( .A(_05368_ ), .Z(_05369_ ) );
OAI21_X1 _13233_ ( .A(_01191_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [30] ), .ZN(_05370_ ) );
AND2_X2 _13234_ ( .A1(_05078_ ), .A2(\IF_ID_inst [31] ), .ZN(_05371_ ) );
AND2_X1 _13235_ ( .A1(_05371_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05372_ ) );
OAI211_X1 _13236_ ( .A(_05170_ ), .B(\IF_ID_inst [31] ), .C1(_05112_ ), .C2(_05012_ ), .ZN(_05373_ ) );
NOR2_X1 _13237_ ( .A1(_05372_ ), .A2(_05373_ ), .ZN(_05374_ ) );
BUF_X4 _13238_ ( .A(_05374_ ), .Z(_05375_ ) );
BUF_X4 _13239_ ( .A(_05375_ ), .Z(_05376_ ) );
INV_X1 _13240_ ( .A(\IF_ID_pc [29] ), .ZN(_05377_ ) );
XNOR2_X1 _13241_ ( .A(_05376_ ), .B(_05377_ ), .ZN(_05378_ ) );
INV_X1 _13242_ ( .A(_05378_ ), .ZN(_05379_ ) );
XNOR2_X1 _13243_ ( .A(_05375_ ), .B(_01388_ ), .ZN(_05380_ ) );
NAND2_X1 _13244_ ( .A1(_05109_ ), .A2(\IF_ID_inst [27] ), .ZN(_05381_ ) );
INV_X1 _13245_ ( .A(_05371_ ), .ZN(_05382_ ) );
OAI21_X1 _13246_ ( .A(_05381_ ), .B1(_05382_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05383_ ) );
XNOR2_X1 _13247_ ( .A(_05383_ ), .B(_01363_ ), .ZN(_05384_ ) );
AND2_X1 _13248_ ( .A1(_05109_ ), .A2(\IF_ID_inst [24] ), .ZN(_05385_ ) );
INV_X1 _13249_ ( .A(_05385_ ), .ZN(_05386_ ) );
OAI21_X1 _13250_ ( .A(_05386_ ), .B1(_05382_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05387_ ) );
NAND2_X1 _13251_ ( .A1(_05387_ ), .A2(\IF_ID_pc [4] ), .ZN(_05388_ ) );
INV_X1 _13252_ ( .A(_05078_ ), .ZN(_05389_ ) );
INV_X1 _13253_ ( .A(\IF_ID_inst [31] ), .ZN(_05390_ ) );
NOR3_X1 _13254_ ( .A1(_05389_ ), .A2(_05390_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_05391_ ) );
AND2_X1 _13255_ ( .A1(_05108_ ), .A2(\IF_ID_inst [23] ), .ZN(_05392_ ) );
NOR2_X1 _13256_ ( .A1(_05391_ ), .A2(_05392_ ), .ZN(_05393_ ) );
NOR3_X2 _13257_ ( .A1(_05389_ ), .A2(_05390_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_05394_ ) );
AND2_X1 _13258_ ( .A1(_05108_ ), .A2(\IF_ID_inst [21] ), .ZN(_05395_ ) );
NOR2_X1 _13259_ ( .A1(_05394_ ), .A2(_05395_ ), .ZN(_05396_ ) );
INV_X1 _13260_ ( .A(\IF_ID_pc [1] ), .ZN(_05397_ ) );
NOR2_X2 _13261_ ( .A1(_05396_ ), .A2(_05397_ ), .ZN(_05398_ ) );
NAND4_X1 _13262_ ( .A1(_05077_ ), .A2(\IF_ID_inst [31] ), .A3(_05012_ ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_05399_ ) );
NAND4_X1 _13263_ ( .A1(_05107_ ), .A2(_05269_ ), .A3(\IF_ID_inst [6] ), .A4(_05070_ ), .ZN(_05400_ ) );
AND3_X1 _13264_ ( .A1(_05399_ ), .A2(_05400_ ), .A3(\IF_ID_pc [2] ), .ZN(_05401_ ) );
AOI21_X1 _13265_ ( .A(\IF_ID_pc [2] ), .B1(_05399_ ), .B2(_05400_ ), .ZN(_05402_ ) );
NOR2_X1 _13266_ ( .A1(_05401_ ), .A2(_05402_ ), .ZN(_05403_ ) );
AND2_X1 _13267_ ( .A1(_05398_ ), .A2(_05403_ ), .ZN(_05404_ ) );
NOR2_X1 _13268_ ( .A1(_05404_ ), .A2(_05401_ ), .ZN(_05405_ ) );
INV_X2 _13269_ ( .A(\IF_ID_pc [3] ), .ZN(_05406_ ) );
XNOR2_X1 _13270_ ( .A(_05393_ ), .B(_05406_ ), .ZN(_05407_ ) );
OAI221_X1 _13271_ ( .A(_05388_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_05393_ ), .C1(_05405_ ), .C2(_05407_ ), .ZN(_05408_ ) );
OR2_X1 _13272_ ( .A1(_05387_ ), .A2(\IF_ID_pc [4] ), .ZN(_05409_ ) );
NAND2_X1 _13273_ ( .A1(_05408_ ), .A2(_05409_ ), .ZN(_05410_ ) );
OR3_X1 _13274_ ( .A1(_05389_ ), .A2(_05390_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_05411_ ) );
NAND3_X1 _13275_ ( .A1(_05077_ ), .A2(\IF_ID_inst [25] ), .A3(_05112_ ), .ZN(_05412_ ) );
NAND2_X1 _13276_ ( .A1(_05411_ ), .A2(_05412_ ), .ZN(_05413_ ) );
XNOR2_X1 _13277_ ( .A(_05413_ ), .B(\IF_ID_pc [5] ), .ZN(_05414_ ) );
AND3_X1 _13278_ ( .A1(_05077_ ), .A2(\IF_ID_inst [26] ), .A3(_05107_ ), .ZN(_05415_ ) );
INV_X1 _13279_ ( .A(_05415_ ), .ZN(_05416_ ) );
OAI21_X1 _13280_ ( .A(_05416_ ), .B1(_05382_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05417_ ) );
XNOR2_X1 _13281_ ( .A(_05417_ ), .B(\IF_ID_pc [6] ), .ZN(_05418_ ) );
NOR3_X2 _13282_ ( .A1(_05410_ ), .A2(_05414_ ), .A3(_05418_ ), .ZN(_05419_ ) );
NAND2_X1 _13283_ ( .A1(_05417_ ), .A2(\IF_ID_pc [6] ), .ZN(_05420_ ) );
NAND2_X1 _13284_ ( .A1(_05413_ ), .A2(_01429_ ), .ZN(_05421_ ) );
OAI21_X1 _13285_ ( .A(_05420_ ), .B1(_05418_ ), .B2(_05421_ ), .ZN(_05422_ ) );
OAI21_X1 _13286_ ( .A(_05384_ ), .B1(_05419_ ), .B2(_05422_ ), .ZN(_05423_ ) );
NAND2_X1 _13287_ ( .A1(_05383_ ), .A2(\IF_ID_pc [7] ), .ZN(_05424_ ) );
NAND2_X1 _13288_ ( .A1(_05423_ ), .A2(_05424_ ), .ZN(_05425_ ) );
NAND3_X1 _13289_ ( .A1(_05170_ ), .A2(\IF_ID_inst [28] ), .A3(_05112_ ), .ZN(_05426_ ) );
OAI21_X1 _13290_ ( .A(_05426_ ), .B1(_05382_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05427_ ) );
OAI21_X1 _13291_ ( .A(_05425_ ), .B1(\IF_ID_pc [8] ), .B2(_05427_ ), .ZN(_05428_ ) );
AND2_X1 _13292_ ( .A1(_05427_ ), .A2(\IF_ID_pc [8] ), .ZN(_05429_ ) );
INV_X1 _13293_ ( .A(_05429_ ), .ZN(_05430_ ) );
NAND2_X2 _13294_ ( .A1(_05428_ ), .A2(_05430_ ), .ZN(_05431_ ) );
NAND3_X1 _13295_ ( .A1(_05077_ ), .A2(\IF_ID_inst [12] ), .A3(_05112_ ), .ZN(_05432_ ) );
AOI21_X1 _13296_ ( .A(_05372_ ), .B1(_05382_ ), .B2(_05432_ ), .ZN(_05433_ ) );
XOR2_X1 _13297_ ( .A(_05433_ ), .B(\IF_ID_pc [12] ), .Z(_05434_ ) );
AND2_X1 _13298_ ( .A1(_05109_ ), .A2(\IF_ID_inst [20] ), .ZN(_05435_ ) );
INV_X1 _13299_ ( .A(_05435_ ), .ZN(_05436_ ) );
OAI21_X1 _13300_ ( .A(_05436_ ), .B1(_05382_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05437_ ) );
INV_X1 _13301_ ( .A(\IF_ID_pc [11] ), .ZN(_05438_ ) );
XNOR2_X1 _13302_ ( .A(_05437_ ), .B(_05438_ ), .ZN(_05439_ ) );
NAND3_X1 _13303_ ( .A1(_05170_ ), .A2(\IF_ID_inst [29] ), .A3(_05112_ ), .ZN(_05440_ ) );
OAI21_X1 _13304_ ( .A(_05440_ ), .B1(_05382_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05441_ ) );
INV_X1 _13305_ ( .A(\IF_ID_pc [9] ), .ZN(_05442_ ) );
XNOR2_X1 _13306_ ( .A(_05441_ ), .B(_05442_ ), .ZN(_05443_ ) );
AND2_X1 _13307_ ( .A1(_05109_ ), .A2(\IF_ID_inst [30] ), .ZN(_05444_ ) );
INV_X1 _13308_ ( .A(_05444_ ), .ZN(_05445_ ) );
OAI21_X1 _13309_ ( .A(_05445_ ), .B1(_05382_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05446_ ) );
XNOR2_X1 _13310_ ( .A(_05446_ ), .B(_01395_ ), .ZN(_05447_ ) );
AND2_X1 _13311_ ( .A1(_05443_ ), .A2(_05447_ ), .ZN(_05448_ ) );
NAND4_X1 _13312_ ( .A1(_05431_ ), .A2(_05434_ ), .A3(_05439_ ), .A4(_05448_ ), .ZN(_05449_ ) );
AND2_X1 _13313_ ( .A1(_05446_ ), .A2(\IF_ID_pc [10] ), .ZN(_05450_ ) );
INV_X1 _13314_ ( .A(_05450_ ), .ZN(_05451_ ) );
INV_X1 _13315_ ( .A(_05447_ ), .ZN(_05452_ ) );
NAND2_X1 _13316_ ( .A1(_05441_ ), .A2(\IF_ID_pc [9] ), .ZN(_05453_ ) );
OAI21_X1 _13317_ ( .A(_05451_ ), .B1(_05452_ ), .B2(_05453_ ), .ZN(_05454_ ) );
AND3_X1 _13318_ ( .A1(_05454_ ), .A2(_05434_ ), .A3(_05439_ ), .ZN(_05455_ ) );
AND2_X1 _13319_ ( .A1(_05433_ ), .A2(\IF_ID_pc [12] ), .ZN(_05456_ ) );
AND2_X1 _13320_ ( .A1(_05437_ ), .A2(\IF_ID_pc [11] ), .ZN(_05457_ ) );
AND2_X1 _13321_ ( .A1(_05434_ ), .A2(_05457_ ), .ZN(_05458_ ) );
NOR3_X1 _13322_ ( .A1(_05455_ ), .A2(_05456_ ), .A3(_05458_ ), .ZN(_05459_ ) );
NAND2_X2 _13323_ ( .A1(_05449_ ), .A2(_05459_ ), .ZN(_05460_ ) );
INV_X1 _13324_ ( .A(_05372_ ), .ZN(_05461_ ) );
OAI22_X1 _13325_ ( .A1(_05110_ ), .A2(_05245_ ), .B1(_05389_ ), .B2(_05390_ ), .ZN(_05462_ ) );
AND2_X1 _13326_ ( .A1(_05461_ ), .A2(_05462_ ), .ZN(_05463_ ) );
XOR2_X1 _13327_ ( .A(_05463_ ), .B(\IF_ID_pc [16] ), .Z(_05464_ ) );
AND3_X1 _13328_ ( .A1(_05170_ ), .A2(\IF_ID_inst [15] ), .A3(_05112_ ), .ZN(_05465_ ) );
INV_X1 _13329_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05466_ ) );
MUX2_X1 _13330_ ( .A(_05465_ ), .B(_05466_ ), .S(_05371_ ), .Z(_05467_ ) );
XOR2_X1 _13331_ ( .A(_05467_ ), .B(\IF_ID_pc [15] ), .Z(_05468_ ) );
AND3_X1 _13332_ ( .A1(_05170_ ), .A2(\IF_ID_inst [13] ), .A3(_05112_ ), .ZN(_05469_ ) );
MUX2_X1 _13333_ ( .A(_05469_ ), .B(_05466_ ), .S(_05371_ ), .Z(_05470_ ) );
XOR2_X1 _13334_ ( .A(_05470_ ), .B(\IF_ID_pc [13] ), .Z(_05471_ ) );
OAI22_X1 _13335_ ( .A1(_05110_ ), .A2(_05130_ ), .B1(_05389_ ), .B2(_05390_ ), .ZN(_05472_ ) );
AND3_X1 _13336_ ( .A1(_05461_ ), .A2(\IF_ID_pc [14] ), .A3(_05472_ ), .ZN(_05473_ ) );
AOI21_X1 _13337_ ( .A(\IF_ID_pc [14] ), .B1(_05461_ ), .B2(_05472_ ), .ZN(_05474_ ) );
NOR2_X1 _13338_ ( .A1(_05473_ ), .A2(_05474_ ), .ZN(_05475_ ) );
AND2_X1 _13339_ ( .A1(_05471_ ), .A2(_05475_ ), .ZN(_05476_ ) );
NAND4_X1 _13340_ ( .A1(_05460_ ), .A2(_05464_ ), .A3(_05468_ ), .A4(_05476_ ), .ZN(_05477_ ) );
AND2_X1 _13341_ ( .A1(_05467_ ), .A2(\IF_ID_pc [15] ), .ZN(_05478_ ) );
AND2_X1 _13342_ ( .A1(_05464_ ), .A2(_05478_ ), .ZN(_05479_ ) );
AOI21_X1 _13343_ ( .A(_05479_ ), .B1(\IF_ID_pc [16] ), .B2(_05463_ ), .ZN(_05480_ ) );
AND2_X1 _13344_ ( .A1(_05470_ ), .A2(\IF_ID_pc [13] ), .ZN(_05481_ ) );
AND2_X1 _13345_ ( .A1(_05475_ ), .A2(_05481_ ), .ZN(_05482_ ) );
OAI211_X1 _13346_ ( .A(_05464_ ), .B(_05468_ ), .C1(_05482_ ), .C2(_05473_ ), .ZN(_05483_ ) );
AND2_X1 _13347_ ( .A1(_05480_ ), .A2(_05483_ ), .ZN(_05484_ ) );
NAND2_X2 _13348_ ( .A1(_05477_ ), .A2(_05484_ ), .ZN(_05485_ ) );
XNOR2_X1 _13349_ ( .A(_05374_ ), .B(_01370_ ), .ZN(_05486_ ) );
AND3_X1 _13350_ ( .A1(_05170_ ), .A2(\IF_ID_inst [19] ), .A3(_05112_ ), .ZN(_05487_ ) );
MUX2_X1 _13351_ ( .A(_05487_ ), .B(_05466_ ), .S(_05371_ ), .Z(_05488_ ) );
XOR2_X1 _13352_ ( .A(_05488_ ), .B(\IF_ID_pc [19] ), .Z(_05489_ ) );
AND3_X1 _13353_ ( .A1(_05170_ ), .A2(\IF_ID_inst [18] ), .A3(_05112_ ), .ZN(_05490_ ) );
MUX2_X1 _13354_ ( .A(_05490_ ), .B(_05466_ ), .S(_05371_ ), .Z(_05491_ ) );
XNOR2_X1 _13355_ ( .A(_05491_ ), .B(_01400_ ), .ZN(_05492_ ) );
OAI22_X1 _13356_ ( .A1(_05110_ ), .A2(_05121_ ), .B1(_05389_ ), .B2(_05390_ ), .ZN(_05493_ ) );
OAI21_X1 _13357_ ( .A(_05493_ ), .B1(_05382_ ), .B2(_05466_ ), .ZN(_05494_ ) );
XNOR2_X1 _13358_ ( .A(_05494_ ), .B(\IF_ID_pc [17] ), .ZN(_05495_ ) );
AND2_X1 _13359_ ( .A1(_05492_ ), .A2(_05495_ ), .ZN(_05496_ ) );
NAND4_X1 _13360_ ( .A1(_05485_ ), .A2(_05486_ ), .A3(_05489_ ), .A4(_05496_ ), .ZN(_05497_ ) );
AND2_X1 _13361_ ( .A1(_05491_ ), .A2(\IF_ID_pc [18] ), .ZN(_05498_ ) );
INV_X1 _13362_ ( .A(_05498_ ), .ZN(_05499_ ) );
NOR2_X1 _13363_ ( .A1(_05491_ ), .A2(\IF_ID_pc [18] ), .ZN(_05500_ ) );
NAND3_X1 _13364_ ( .A1(_05461_ ), .A2(\IF_ID_pc [17] ), .A3(_05493_ ), .ZN(_05501_ ) );
OAI21_X1 _13365_ ( .A(_05499_ ), .B1(_05500_ ), .B2(_05501_ ), .ZN(_05502_ ) );
NAND3_X1 _13366_ ( .A1(_05502_ ), .A2(_05486_ ), .A3(_05489_ ), .ZN(_05503_ ) );
OR3_X1 _13367_ ( .A1(_05372_ ), .A2(_01370_ ), .A3(_05373_ ), .ZN(_05504_ ) );
NAND3_X1 _13368_ ( .A1(_05486_ ), .A2(\IF_ID_pc [19] ), .A3(_05488_ ), .ZN(_05505_ ) );
AND3_X1 _13369_ ( .A1(_05503_ ), .A2(_05504_ ), .A3(_05505_ ), .ZN(_05506_ ) );
AND2_X2 _13370_ ( .A1(_05497_ ), .A2(_05506_ ), .ZN(_05507_ ) );
INV_X1 _13371_ ( .A(_05507_ ), .ZN(_05508_ ) );
XNOR2_X1 _13372_ ( .A(_05374_ ), .B(_01379_ ), .ZN(_05509_ ) );
XNOR2_X1 _13373_ ( .A(_05374_ ), .B(_01402_ ), .ZN(_05510_ ) );
AND2_X1 _13374_ ( .A1(_05509_ ), .A2(_05510_ ), .ZN(_05511_ ) );
XNOR2_X1 _13375_ ( .A(_05375_ ), .B(_01478_ ), .ZN(_05512_ ) );
XNOR2_X1 _13376_ ( .A(_05374_ ), .B(_01420_ ), .ZN(_05513_ ) );
AND2_X1 _13377_ ( .A1(_05512_ ), .A2(_05513_ ), .ZN(_05514_ ) );
AND3_X2 _13378_ ( .A1(_05508_ ), .A2(_05511_ ), .A3(_05514_ ), .ZN(_05515_ ) );
AND2_X1 _13379_ ( .A1(_05375_ ), .A2(\IF_ID_pc [22] ), .ZN(_05516_ ) );
AND2_X1 _13380_ ( .A1(_05375_ ), .A2(\IF_ID_pc [21] ), .ZN(_05517_ ) );
OAI21_X1 _13381_ ( .A(_05511_ ), .B1(_05516_ ), .B2(_05517_ ), .ZN(_05518_ ) );
NAND2_X1 _13382_ ( .A1(_05375_ ), .A2(\IF_ID_pc [24] ), .ZN(_05519_ ) );
NAND2_X1 _13383_ ( .A1(_05375_ ), .A2(\IF_ID_pc [23] ), .ZN(_05520_ ) );
AND3_X1 _13384_ ( .A1(_05518_ ), .A2(_05519_ ), .A3(_05520_ ), .ZN(_05521_ ) );
INV_X1 _13385_ ( .A(_05521_ ), .ZN(_05522_ ) );
OAI21_X1 _13386_ ( .A(_05380_ ), .B1(_05515_ ), .B2(_05522_ ), .ZN(_05523_ ) );
XNOR2_X1 _13387_ ( .A(_05376_ ), .B(_01471_ ), .ZN(_05524_ ) );
INV_X1 _13388_ ( .A(_05524_ ), .ZN(_05525_ ) );
NOR2_X2 _13389_ ( .A1(_05523_ ), .A2(_05525_ ), .ZN(_05526_ ) );
XOR2_X1 _13390_ ( .A(_05375_ ), .B(\IF_ID_pc [28] ), .Z(_05527_ ) );
XNOR2_X1 _13391_ ( .A(_05375_ ), .B(_01345_ ), .ZN(_05528_ ) );
AND2_X1 _13392_ ( .A1(_05527_ ), .A2(_05528_ ), .ZN(_05529_ ) );
NAND2_X1 _13393_ ( .A1(_05526_ ), .A2(_05529_ ), .ZN(_05530_ ) );
AND2_X1 _13394_ ( .A1(_05375_ ), .A2(\IF_ID_pc [27] ), .ZN(_05531_ ) );
OAI21_X1 _13395_ ( .A(_05376_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_05532_ ) );
INV_X1 _13396_ ( .A(_05532_ ), .ZN(_05533_ ) );
AOI221_X4 _13397_ ( .A(_05531_ ), .B1(\IF_ID_pc [28] ), .B2(_05376_ ), .C1(_05529_ ), .C2(_05533_ ), .ZN(_05534_ ) );
AOI21_X2 _13398_ ( .A(_05379_ ), .B1(_05530_ ), .B2(_05534_ ), .ZN(_05535_ ) );
NOR3_X1 _13399_ ( .A1(_05372_ ), .A2(_05377_ ), .A3(_05373_ ), .ZN(_05536_ ) );
NOR2_X1 _13400_ ( .A1(_05535_ ), .A2(_05536_ ), .ZN(_05537_ ) );
XNOR2_X1 _13401_ ( .A(_05376_ ), .B(\IF_ID_pc [30] ), .ZN(_05538_ ) );
XNOR2_X1 _13402_ ( .A(_05537_ ), .B(_05538_ ), .ZN(_05539_ ) );
BUF_X4 _13403_ ( .A(_05368_ ), .Z(_05540_ ) );
BUF_X4 _13404_ ( .A(_05540_ ), .Z(_05541_ ) );
AOI21_X1 _13405_ ( .A(_05370_ ), .B1(_05539_ ), .B2(_05541_ ), .ZN(_00243_ ) );
XNOR2_X1 _13406_ ( .A(_05507_ ), .B(_05513_ ), .ZN(_05542_ ) );
NOR2_X1 _13407_ ( .A1(_05542_ ), .A2(_05367_ ), .ZN(_05543_ ) );
BUF_X4 _13408_ ( .A(_05367_ ), .Z(_05544_ ) );
AOI211_X1 _13409_ ( .A(fanout_net_5 ), .B(_05543_ ), .C1(_05214_ ), .C2(_05544_ ), .ZN(_00244_ ) );
OAI21_X1 _13410_ ( .A(_01191_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [20] ), .ZN(_05545_ ) );
AND2_X1 _13411_ ( .A1(_05485_ ), .A2(_05496_ ), .ZN(_05546_ ) );
OAI21_X1 _13412_ ( .A(_05489_ ), .B1(_05546_ ), .B2(_05502_ ), .ZN(_05547_ ) );
NAND2_X1 _13413_ ( .A1(_05488_ ), .A2(\IF_ID_pc [19] ), .ZN(_05548_ ) );
AND2_X1 _13414_ ( .A1(_05547_ ), .A2(_05548_ ), .ZN(_05549_ ) );
OR2_X1 _13415_ ( .A1(_05549_ ), .A2(_05486_ ), .ZN(_05550_ ) );
AOI21_X1 _13416_ ( .A(_05544_ ), .B1(_05549_ ), .B2(_05486_ ), .ZN(_05551_ ) );
AOI21_X1 _13417_ ( .A(_05545_ ), .B1(_05550_ ), .B2(_05551_ ), .ZN(_00245_ ) );
OAI21_X1 _13418_ ( .A(_01191_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [19] ), .ZN(_05552_ ) );
OR2_X1 _13419_ ( .A1(_05546_ ), .A2(_05502_ ), .ZN(_05553_ ) );
XNOR2_X1 _13420_ ( .A(_05553_ ), .B(_05489_ ), .ZN(_05554_ ) );
AOI21_X1 _13421_ ( .A(_05552_ ), .B1(_05554_ ), .B2(_05541_ ), .ZN(_00246_ ) );
OAI21_X1 _13422_ ( .A(_01191_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [18] ), .ZN(_05555_ ) );
NAND2_X1 _13423_ ( .A1(_05485_ ), .A2(_05495_ ), .ZN(_05556_ ) );
NAND2_X1 _13424_ ( .A1(_05556_ ), .A2(_05501_ ), .ZN(_05557_ ) );
XNOR2_X1 _13425_ ( .A(_05557_ ), .B(_05492_ ), .ZN(_05558_ ) );
AOI21_X1 _13426_ ( .A(_05555_ ), .B1(_05558_ ), .B2(_05541_ ), .ZN(_00247_ ) );
OAI21_X1 _13427_ ( .A(_01191_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [17] ), .ZN(_05559_ ) );
XNOR2_X1 _13428_ ( .A(_05485_ ), .B(_05495_ ), .ZN(_05560_ ) );
AOI21_X1 _13429_ ( .A(_05559_ ), .B1(_05560_ ), .B2(_05541_ ), .ZN(_00248_ ) );
OAI21_X1 _13430_ ( .A(_01191_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [16] ), .ZN(_05561_ ) );
NAND2_X1 _13431_ ( .A1(_05460_ ), .A2(_05476_ ), .ZN(_05562_ ) );
AOI21_X1 _13432_ ( .A(_05473_ ), .B1(_05475_ ), .B2(_05481_ ), .ZN(_05563_ ) );
NAND2_X1 _13433_ ( .A1(_05562_ ), .A2(_05563_ ), .ZN(_05564_ ) );
AND2_X1 _13434_ ( .A1(_05564_ ), .A2(_05468_ ), .ZN(_05565_ ) );
OR2_X1 _13435_ ( .A1(_05565_ ), .A2(_05478_ ), .ZN(_05566_ ) );
XNOR2_X1 _13436_ ( .A(_05566_ ), .B(_05464_ ), .ZN(_05567_ ) );
AOI21_X1 _13437_ ( .A(_05561_ ), .B1(_05567_ ), .B2(_05541_ ), .ZN(_00249_ ) );
OAI21_X1 _13438_ ( .A(_01191_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [15] ), .ZN(_05568_ ) );
XNOR2_X1 _13439_ ( .A(_05564_ ), .B(_05468_ ), .ZN(_05569_ ) );
AOI21_X1 _13440_ ( .A(_05568_ ), .B1(_05569_ ), .B2(_05541_ ), .ZN(_00250_ ) );
BUF_X4 _13441_ ( .A(_01147_ ), .Z(_05570_ ) );
OAI21_X1 _13442_ ( .A(_05570_ ), .B1(_05369_ ), .B2(\myexu.pc_jump [14] ), .ZN(_05571_ ) );
AND2_X1 _13443_ ( .A1(_05460_ ), .A2(_05471_ ), .ZN(_05572_ ) );
NOR2_X1 _13444_ ( .A1(_05572_ ), .A2(_05481_ ), .ZN(_05573_ ) );
OR2_X1 _13445_ ( .A1(_05573_ ), .A2(_05475_ ), .ZN(_05574_ ) );
AOI21_X1 _13446_ ( .A(_05544_ ), .B1(_05573_ ), .B2(_05475_ ), .ZN(_05575_ ) );
AOI21_X1 _13447_ ( .A(_05571_ ), .B1(_05574_ ), .B2(_05575_ ), .ZN(_00251_ ) );
BUF_X4 _13448_ ( .A(_05368_ ), .Z(_05576_ ) );
OAI21_X1 _13449_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [13] ), .ZN(_05577_ ) );
XNOR2_X1 _13450_ ( .A(_05460_ ), .B(_05471_ ), .ZN(_05578_ ) );
AOI21_X1 _13451_ ( .A(_05577_ ), .B1(_05578_ ), .B2(_05541_ ), .ZN(_00252_ ) );
OAI21_X1 _13452_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [12] ), .ZN(_05579_ ) );
NAND2_X1 _13453_ ( .A1(_05431_ ), .A2(_05448_ ), .ZN(_05580_ ) );
INV_X1 _13454_ ( .A(_05454_ ), .ZN(_05581_ ) );
NAND2_X1 _13455_ ( .A1(_05580_ ), .A2(_05581_ ), .ZN(_05582_ ) );
AND2_X1 _13456_ ( .A1(_05582_ ), .A2(_05439_ ), .ZN(_05583_ ) );
OR2_X1 _13457_ ( .A1(_05583_ ), .A2(_05457_ ), .ZN(_05584_ ) );
XNOR2_X1 _13458_ ( .A(_05584_ ), .B(_05434_ ), .ZN(_05585_ ) );
AOI21_X1 _13459_ ( .A(_05579_ ), .B1(_05585_ ), .B2(_05541_ ), .ZN(_00253_ ) );
OAI21_X1 _13460_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [29] ), .ZN(_05586_ ) );
AND2_X1 _13461_ ( .A1(_05530_ ), .A2(_05534_ ), .ZN(_05587_ ) );
XNOR2_X1 _13462_ ( .A(_05587_ ), .B(_05379_ ), .ZN(_05588_ ) );
AOI21_X1 _13463_ ( .A(_05586_ ), .B1(_05588_ ), .B2(_05541_ ), .ZN(_00254_ ) );
OAI21_X1 _13464_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [11] ), .ZN(_05589_ ) );
XNOR2_X1 _13465_ ( .A(_05582_ ), .B(_05439_ ), .ZN(_05590_ ) );
AOI21_X1 _13466_ ( .A(_05589_ ), .B1(_05590_ ), .B2(_05541_ ), .ZN(_00255_ ) );
OAI21_X1 _13467_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [10] ), .ZN(_05591_ ) );
NAND2_X1 _13468_ ( .A1(_05431_ ), .A2(_05443_ ), .ZN(_05592_ ) );
NAND2_X1 _13469_ ( .A1(_05592_ ), .A2(_05453_ ), .ZN(_05593_ ) );
XNOR2_X1 _13470_ ( .A(_05593_ ), .B(_05447_ ), .ZN(_05594_ ) );
BUF_X4 _13471_ ( .A(_05540_ ), .Z(_05595_ ) );
AOI21_X1 _13472_ ( .A(_05591_ ), .B1(_05594_ ), .B2(_05595_ ), .ZN(_00256_ ) );
OAI21_X1 _13473_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [9] ), .ZN(_05596_ ) );
XNOR2_X1 _13474_ ( .A(_05431_ ), .B(_05443_ ), .ZN(_05597_ ) );
AOI21_X1 _13475_ ( .A(_05596_ ), .B1(_05597_ ), .B2(_05595_ ), .ZN(_00257_ ) );
OAI21_X1 _13476_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [8] ), .ZN(_05598_ ) );
XNOR2_X1 _13477_ ( .A(_05427_ ), .B(_05212_ ), .ZN(_05599_ ) );
XNOR2_X1 _13478_ ( .A(_05425_ ), .B(_05599_ ), .ZN(_05600_ ) );
AOI21_X1 _13479_ ( .A(_05598_ ), .B1(_05600_ ), .B2(_05595_ ), .ZN(_00258_ ) );
OAI21_X1 _13480_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [7] ), .ZN(_05601_ ) );
OR2_X1 _13481_ ( .A1(_05419_ ), .A2(_05422_ ), .ZN(_05602_ ) );
XNOR2_X1 _13482_ ( .A(_05602_ ), .B(_05384_ ), .ZN(_05603_ ) );
AOI21_X1 _13483_ ( .A(_05601_ ), .B1(_05603_ ), .B2(_05595_ ), .ZN(_00259_ ) );
OAI21_X1 _13484_ ( .A(_05570_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [6] ), .ZN(_05604_ ) );
OR2_X1 _13485_ ( .A1(_05410_ ), .A2(_05414_ ), .ZN(_05605_ ) );
AND2_X1 _13486_ ( .A1(_05605_ ), .A2(_05421_ ), .ZN(_05606_ ) );
XNOR2_X1 _13487_ ( .A(_05606_ ), .B(_05418_ ), .ZN(_05607_ ) );
AOI21_X1 _13488_ ( .A(_05604_ ), .B1(_05607_ ), .B2(_05595_ ), .ZN(_00260_ ) );
BUF_X4 _13489_ ( .A(_01051_ ), .Z(_05608_ ) );
OAI21_X1 _13490_ ( .A(_05608_ ), .B1(_05576_ ), .B2(\myexu.pc_jump [5] ), .ZN(_05609_ ) );
XNOR2_X1 _13491_ ( .A(_05410_ ), .B(_05414_ ), .ZN(_05610_ ) );
AOI21_X1 _13492_ ( .A(_05609_ ), .B1(_05610_ ), .B2(_05595_ ), .ZN(_00261_ ) );
NOR2_X1 _13493_ ( .A1(_05405_ ), .A2(_05407_ ), .ZN(_05611_ ) );
NOR2_X1 _13494_ ( .A1(_05393_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05612_ ) );
OAI211_X1 _13495_ ( .A(_05388_ ), .B(_05409_ ), .C1(_05611_ ), .C2(_05612_ ), .ZN(_05613_ ) );
XNOR2_X1 _13496_ ( .A(_05387_ ), .B(\IF_ID_pc [4] ), .ZN(_05614_ ) );
OAI221_X1 _13497_ ( .A(_05614_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_05393_ ), .C1(_05405_ ), .C2(_05407_ ), .ZN(_05615_ ) );
AND3_X1 _13498_ ( .A1(_05613_ ), .A2(_05368_ ), .A3(_05615_ ), .ZN(_05616_ ) );
AOI21_X1 _13499_ ( .A(_05616_ ), .B1(\myexu.pc_jump [4] ), .B2(_05544_ ), .ZN(_05617_ ) );
NOR2_X1 _13500_ ( .A1(_05617_ ), .A2(fanout_net_5 ), .ZN(_00262_ ) );
AND2_X1 _13501_ ( .A1(_05405_ ), .A2(_05407_ ), .ZN(_05618_ ) );
NOR3_X1 _13502_ ( .A1(_05618_ ), .A2(_05611_ ), .A3(_05367_ ), .ZN(_05619_ ) );
AOI21_X1 _13503_ ( .A(_05619_ ), .B1(\myexu.pc_jump [3] ), .B2(_05544_ ), .ZN(_05620_ ) );
NOR2_X1 _13504_ ( .A1(_05620_ ), .A2(fanout_net_5 ), .ZN(_00263_ ) );
AOI211_X1 _13505_ ( .A(_05187_ ), .B(_05616_ ), .C1(\myexu.pc_jump [4] ), .C2(_05367_ ), .ZN(_05621_ ) );
INV_X1 _13506_ ( .A(\IF_ID_pc [4] ), .ZN(_05622_ ) );
BUF_X2 _13507_ ( .A(_05622_ ), .Z(_05623_ ) );
AOI211_X1 _13508_ ( .A(fanout_net_5 ), .B(_05621_ ), .C1(_05623_ ), .C2(_05187_ ), .ZN(_00264_ ) );
OAI21_X1 _13509_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [2] ), .ZN(_05624_ ) );
XNOR2_X1 _13510_ ( .A(_05398_ ), .B(_05403_ ), .ZN(_05625_ ) );
AOI21_X1 _13511_ ( .A(_05624_ ), .B1(_05625_ ), .B2(_05595_ ), .ZN(_00265_ ) );
AOI211_X1 _13512_ ( .A(_05187_ ), .B(_05619_ ), .C1(\myexu.pc_jump [3] ), .C2(_05367_ ), .ZN(_05626_ ) );
BUF_X2 _13513_ ( .A(_05406_ ), .Z(_05627_ ) );
AOI211_X1 _13514_ ( .A(fanout_net_5 ), .B(_05626_ ), .C1(_05627_ ), .C2(_05187_ ), .ZN(_00266_ ) );
OAI21_X1 _13515_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [28] ), .ZN(_05628_ ) );
OAI21_X1 _13516_ ( .A(_05528_ ), .B1(_05526_ ), .B2(_05533_ ), .ZN(_05629_ ) );
INV_X1 _13517_ ( .A(_05531_ ), .ZN(_05630_ ) );
AND2_X1 _13518_ ( .A1(_05629_ ), .A2(_05630_ ), .ZN(_05631_ ) );
OR2_X1 _13519_ ( .A1(_05631_ ), .A2(_05527_ ), .ZN(_05632_ ) );
AOI21_X1 _13520_ ( .A(_05544_ ), .B1(_05631_ ), .B2(_05527_ ), .ZN(_05633_ ) );
AOI21_X1 _13521_ ( .A(_05628_ ), .B1(_05632_ ), .B2(_05633_ ), .ZN(_00267_ ) );
OR3_X1 _13522_ ( .A1(_05237_ ), .A2(_01641_ ), .A3(\myexu.pc_jump [1] ), .ZN(_05634_ ) );
INV_X1 _13523_ ( .A(_05634_ ), .ZN(_05635_ ) );
XNOR2_X1 _13524_ ( .A(_05396_ ), .B(_05397_ ), .ZN(_05636_ ) );
AOI211_X1 _13525_ ( .A(fanout_net_5 ), .B(_05635_ ), .C1(_05369_ ), .C2(_05636_ ), .ZN(_00268_ ) );
OAI21_X1 _13526_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [27] ), .ZN(_05637_ ) );
NOR2_X1 _13527_ ( .A1(_05526_ ), .A2(_05533_ ), .ZN(_05638_ ) );
XOR2_X1 _13528_ ( .A(_05638_ ), .B(_05528_ ), .Z(_05639_ ) );
AOI21_X1 _13529_ ( .A(_05637_ ), .B1(_05639_ ), .B2(_05595_ ), .ZN(_00269_ ) );
OAI21_X1 _13530_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [26] ), .ZN(_05640_ ) );
NAND2_X1 _13531_ ( .A1(_05376_ ), .A2(\IF_ID_pc [25] ), .ZN(_05641_ ) );
AND2_X1 _13532_ ( .A1(_05523_ ), .A2(_05641_ ), .ZN(_05642_ ) );
OR2_X1 _13533_ ( .A1(_05642_ ), .A2(_05524_ ), .ZN(_05643_ ) );
AOI21_X1 _13534_ ( .A(_05544_ ), .B1(_05642_ ), .B2(_05524_ ), .ZN(_05644_ ) );
AOI21_X1 _13535_ ( .A(_05640_ ), .B1(_05643_ ), .B2(_05644_ ), .ZN(_00270_ ) );
OAI21_X1 _13536_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [25] ), .ZN(_05645_ ) );
NOR2_X1 _13537_ ( .A1(_05515_ ), .A2(_05522_ ), .ZN(_05646_ ) );
XOR2_X1 _13538_ ( .A(_05646_ ), .B(_05380_ ), .Z(_05647_ ) );
AOI21_X1 _13539_ ( .A(_05645_ ), .B1(_05647_ ), .B2(_05595_ ), .ZN(_00271_ ) );
OAI21_X1 _13540_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [24] ), .ZN(_05648_ ) );
NAND2_X1 _13541_ ( .A1(_05508_ ), .A2(_05514_ ), .ZN(_05649_ ) );
OAI21_X1 _13542_ ( .A(_05376_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_05650_ ) );
NAND2_X1 _13543_ ( .A1(_05649_ ), .A2(_05650_ ), .ZN(_05651_ ) );
NAND2_X1 _13544_ ( .A1(_05651_ ), .A2(_05510_ ), .ZN(_05652_ ) );
AND2_X1 _13545_ ( .A1(_05652_ ), .A2(_05520_ ), .ZN(_05653_ ) );
OR2_X1 _13546_ ( .A1(_05653_ ), .A2(_05509_ ), .ZN(_05654_ ) );
AOI21_X1 _13547_ ( .A(_05367_ ), .B1(_05653_ ), .B2(_05509_ ), .ZN(_05655_ ) );
AOI21_X1 _13548_ ( .A(_05648_ ), .B1(_05654_ ), .B2(_05655_ ), .ZN(_00272_ ) );
OAI21_X1 _13549_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [23] ), .ZN(_05656_ ) );
XNOR2_X1 _13550_ ( .A(_05651_ ), .B(_05510_ ), .ZN(_05657_ ) );
AOI21_X1 _13551_ ( .A(_05656_ ), .B1(_05657_ ), .B2(_05595_ ), .ZN(_00273_ ) );
OAI21_X1 _13552_ ( .A(_05608_ ), .B1(_05540_ ), .B2(\myexu.pc_jump [22] ), .ZN(_05658_ ) );
INV_X1 _13553_ ( .A(_05513_ ), .ZN(_05659_ ) );
AOI21_X1 _13554_ ( .A(_05659_ ), .B1(_05497_ ), .B2(_05506_ ), .ZN(_05660_ ) );
NOR2_X1 _13555_ ( .A1(_05660_ ), .A2(_05517_ ), .ZN(_05661_ ) );
OR2_X1 _13556_ ( .A1(_05661_ ), .A2(_05512_ ), .ZN(_05662_ ) );
AOI21_X1 _13557_ ( .A(_05367_ ), .B1(_05661_ ), .B2(_05512_ ), .ZN(_05663_ ) );
AOI21_X1 _13558_ ( .A(_05658_ ), .B1(_05662_ ), .B2(_05663_ ), .ZN(_00274_ ) );
AOI211_X1 _13559_ ( .A(_05536_ ), .B(_05535_ ), .C1(\IF_ID_pc [30] ), .C2(_05376_ ), .ZN(_05664_ ) );
NOR2_X1 _13560_ ( .A1(_05376_ ), .A2(\IF_ID_pc [30] ), .ZN(_05665_ ) );
XNOR2_X1 _13561_ ( .A(_05376_ ), .B(\IF_ID_pc [31] ), .ZN(_05666_ ) );
OR3_X4 _13562_ ( .A1(_05664_ ), .A2(_05665_ ), .A3(_05666_ ), .ZN(_05667_ ) );
OAI21_X1 _13563_ ( .A(_05666_ ), .B1(_05664_ ), .B2(_05665_ ), .ZN(_05668_ ) );
NAND3_X1 _13564_ ( .A1(_05667_ ), .A2(_05369_ ), .A3(_05668_ ), .ZN(_05669_ ) );
NAND3_X1 _13565_ ( .A1(_05238_ ), .A2(check_quest ), .A3(\myexu.pc_jump [31] ), .ZN(_05670_ ) );
NAND3_X1 _13566_ ( .A1(_05669_ ), .A2(_01329_ ), .A3(_05670_ ), .ZN(_00275_ ) );
AND4_X1 _13567_ ( .A1(_01590_ ), .A2(_01594_ ), .A3(_01572_ ), .A4(_01576_ ), .ZN(_05671_ ) );
AND4_X1 _13568_ ( .A1(_01580_ ), .A2(_01584_ ), .A3(_01551_ ), .A4(_01559_ ), .ZN(_05672_ ) );
NAND2_X1 _13569_ ( .A1(_05671_ ), .A2(_05672_ ), .ZN(_05673_ ) );
AND4_X1 _13570_ ( .A1(_01611_ ), .A2(_01615_ ), .A3(_01563_ ), .A4(_01567_ ), .ZN(_05674_ ) );
AND4_X1 _13571_ ( .A1(_01598_ ), .A2(_01602_ ), .A3(_01607_ ), .A4(\io_master_araddr [25] ), .ZN(_05675_ ) );
NAND2_X1 _13572_ ( .A1(_05674_ ), .A2(_05675_ ), .ZN(_05676_ ) );
NOR2_X1 _13573_ ( .A1(_05673_ ), .A2(_05676_ ), .ZN(_05677_ ) );
INV_X1 _13574_ ( .A(_05677_ ), .ZN(_05678_ ) );
NOR2_X1 _13575_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_05679_ ) );
NOR2_X1 _13576_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_05680_ ) );
INV_X1 _13577_ ( .A(\io_master_rid [1] ), .ZN(_05681_ ) );
NAND4_X1 _13578_ ( .A1(_05679_ ), .A2(_05680_ ), .A3(_05681_ ), .A4(\io_master_rid [0] ), .ZN(_05682_ ) );
AOI21_X1 _13579_ ( .A(_01618_ ), .B1(_05678_ ), .B2(_05682_ ), .ZN(_05683_ ) );
NAND4_X1 _13580_ ( .A1(_01590_ ), .A2(_01572_ ), .A3(_01580_ ), .A4(_01598_ ), .ZN(_05684_ ) );
NAND4_X1 _13581_ ( .A1(_01594_ ), .A2(_01576_ ), .A3(_01584_ ), .A4(_01602_ ), .ZN(_05685_ ) );
NOR2_X2 _13582_ ( .A1(_05684_ ), .A2(_05685_ ), .ZN(_05686_ ) );
NAND4_X4 _13583_ ( .A1(_01551_ ), .A2(_01607_ ), .A3(_01611_ ), .A4(_01563_ ), .ZN(_05687_ ) );
NAND4_X4 _13584_ ( .A1(_01559_ ), .A2(_01615_ ), .A3(_01567_ ), .A4(\io_master_araddr [25] ), .ZN(_05688_ ) );
NOR2_X4 _13585_ ( .A1(_05687_ ), .A2(_05688_ ), .ZN(_05689_ ) );
AND3_X1 _13586_ ( .A1(_05686_ ), .A2(_05689_ ), .A3(\myclint.state_r_$_NOT__A_Y ), .ZN(_05690_ ) );
AOI21_X1 _13587_ ( .A(io_master_rvalid ), .B1(_05686_ ), .B2(_05689_ ), .ZN(_05691_ ) );
NOR2_X1 _13588_ ( .A1(_05690_ ), .A2(_05691_ ), .ZN(_05692_ ) );
AND2_X1 _13589_ ( .A1(_05683_ ), .A2(_05692_ ), .ZN(_05693_ ) );
BUF_X4 _13590_ ( .A(_05693_ ), .Z(_05694_ ) );
BUF_X4 _13591_ ( .A(_05694_ ), .Z(_05695_ ) );
AND2_X4 _13592_ ( .A1(_05686_ ), .A2(_05689_ ), .ZN(_05696_ ) );
BUF_X4 _13593_ ( .A(_05696_ ), .Z(_05697_ ) );
BUF_X4 _13594_ ( .A(_05697_ ), .Z(_05698_ ) );
BUF_X4 _13595_ ( .A(_05698_ ), .Z(_05699_ ) );
OAI21_X1 _13596_ ( .A(_05695_ ), .B1(io_master_rlast ), .B2(_05699_ ), .ZN(_05700_ ) );
INV_X1 _13597_ ( .A(\myifu.tmp_offset [2] ), .ZN(_05701_ ) );
AND3_X1 _13598_ ( .A1(_05700_ ), .A2(_01148_ ), .A3(_05701_ ), .ZN(_00276_ ) );
NOR2_X1 _13599_ ( .A1(_01549_ ), .A2(fanout_net_5 ), .ZN(_00277_ ) );
AND2_X1 _13600_ ( .A1(_01246_ ), .A2(\EX_LS_pc [2] ), .ZN(_00278_ ) );
INV_X1 _13601_ ( .A(\mylsu.state [3] ), .ZN(_05702_ ) );
NOR2_X1 _13602_ ( .A1(_05702_ ), .A2(fanout_net_5 ), .ZN(_00279_ ) );
INV_X1 _13603_ ( .A(_01678_ ), .ZN(_05703_ ) );
OAI211_X1 _13604_ ( .A(_05703_ ), .B(_01674_ ), .C1(\EX_LS_flag [2] ), .C2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_05704_ ) );
CLKBUF_X2 _13605_ ( .A(_05704_ ), .Z(_05705_ ) );
AND2_X1 _13606_ ( .A1(_01678_ ), .A2(_01679_ ), .ZN(_05706_ ) );
INV_X1 _13607_ ( .A(_05706_ ), .ZN(_05707_ ) );
CLKBUF_X2 _13608_ ( .A(_05707_ ), .Z(_05708_ ) );
AND3_X1 _13609_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(\EX_LS_dest_csreg_mem [11] ), .ZN(_00280_ ) );
AND3_X1 _13610_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(\EX_LS_dest_csreg_mem [10] ), .ZN(_00281_ ) );
AND3_X1 _13611_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(\EX_LS_dest_csreg_mem [7] ), .ZN(_00282_ ) );
AND3_X1 _13612_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(\EX_LS_dest_csreg_mem [5] ), .ZN(_00283_ ) );
AND3_X1 _13613_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(\EX_LS_dest_csreg_mem [4] ), .ZN(_00284_ ) );
AND3_X1 _13614_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(\EX_LS_dest_csreg_mem [3] ), .ZN(_00285_ ) );
AND3_X1 _13615_ ( .A1(_05704_ ), .A2(_05707_ ), .A3(\EX_LS_dest_csreg_mem [2] ), .ZN(_00286_ ) );
AND3_X1 _13616_ ( .A1(_05704_ ), .A2(_05707_ ), .A3(fanout_net_7 ), .ZN(_00287_ ) );
INV_X1 _13617_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_05709_ ) );
NAND3_X1 _13618_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(_05709_ ), .ZN(_00288_ ) );
INV_X1 _13619_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_05710_ ) );
NAND3_X1 _13620_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(_05710_ ), .ZN(_00289_ ) );
INV_X1 _13621_ ( .A(\EX_LS_dest_csreg_mem [6] ), .ZN(_05711_ ) );
NAND3_X1 _13622_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(_05711_ ), .ZN(_00290_ ) );
INV_X1 _13623_ ( .A(fanout_net_6 ), .ZN(_05712_ ) );
NAND3_X1 _13624_ ( .A1(_05705_ ), .A2(_05708_ ), .A3(_05712_ ), .ZN(_00291_ ) );
NOR2_X1 _13625_ ( .A1(\mylsu.state [3] ), .A2(\mylsu.state [1] ), .ZN(_05713_ ) );
INV_X1 _13626_ ( .A(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_05714_ ) );
NAND3_X1 _13627_ ( .A1(_05713_ ), .A2(_05608_ ), .A3(_05714_ ), .ZN(_05715_ ) );
NAND3_X1 _13628_ ( .A1(_04995_ ), .A2(_04997_ ), .A3(_01623_ ), .ZN(_05716_ ) );
NAND3_X1 _13629_ ( .A1(_05716_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_flag [1] ), .ZN(_05717_ ) );
NOR2_X1 _13630_ ( .A1(_01679_ ), .A2(\EX_LS_flag [1] ), .ZN(_05718_ ) );
AND2_X1 _13631_ ( .A1(_05718_ ), .A2(_01673_ ), .ZN(_05719_ ) );
INV_X1 _13632_ ( .A(_05719_ ), .ZN(_05720_ ) );
AOI21_X1 _13633_ ( .A(_05715_ ), .B1(_05717_ ), .B2(_05720_ ), .ZN(_00292_ ) );
OR2_X1 _13634_ ( .A1(_05717_ ), .A2(_01673_ ), .ZN(_05721_ ) );
AOI21_X1 _13635_ ( .A(_05715_ ), .B1(_05721_ ), .B2(_05720_ ), .ZN(_00293_ ) );
NAND3_X1 _13636_ ( .A1(_05713_ ), .A2(_01147_ ), .A3(EXU_valid_LSU ), .ZN(_05722_ ) );
NOR3_X1 _13637_ ( .A1(_05717_ ), .A2(_01673_ ), .A3(_05722_ ), .ZN(_00294_ ) );
INV_X1 _13638_ ( .A(_00279_ ), .ZN(_05723_ ) );
NOR3_X1 _13639_ ( .A1(_01673_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_flag [1] ), .ZN(_05724_ ) );
NOR3_X1 _13640_ ( .A1(_05706_ ), .A2(_05724_ ), .A3(_01676_ ), .ZN(_05725_ ) );
OAI21_X1 _13641_ ( .A(_05723_ ), .B1(_05725_ ), .B2(_05722_ ), .ZN(_00295_ ) );
INV_X1 _13642_ ( .A(\mysc.state [2] ), .ZN(_05726_ ) );
NOR2_X1 _13643_ ( .A1(_05726_ ), .A2(fanout_net_5 ), .ZN(_00296_ ) );
AND2_X1 _13644_ ( .A1(_01624_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_05727_ ) );
CLKBUF_X2 _13645_ ( .A(_05727_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X1 _13646_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .ZN(_05728_ ) );
AND3_X1 _13647_ ( .A1(_01624_ ), .A2(_05728_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00239_ ) );
AND3_X1 _13648_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05623_ ), .A3(\IF_ID_pc [3] ), .ZN(_00240_ ) );
AND3_X1 _13649_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_05627_ ), .ZN(_00241_ ) );
CLKBUF_X2 _13650_ ( .A(_01533_ ), .Z(_05729_ ) );
CLKBUF_X2 _13651_ ( .A(_05729_ ), .Z(_05730_ ) );
CLKBUF_X2 _13652_ ( .A(_05730_ ), .Z(_05731_ ) );
BUF_X2 _13653_ ( .A(_05731_ ), .Z(\io_master_arburst [0] ) );
BUF_X2 _13654_ ( .A(_01542_ ), .Z(_05732_ ) );
BUF_X2 _13655_ ( .A(_01543_ ), .Z(_05733_ ) );
NOR3_X1 _13656_ ( .A1(_05732_ ), .A2(fanout_net_7 ), .A3(_05733_ ), .ZN(_05734_ ) );
INV_X1 _13657_ ( .A(_01540_ ), .ZN(_05735_ ) );
BUF_X2 _13658_ ( .A(_05735_ ), .Z(_05736_ ) );
BUF_X2 _13659_ ( .A(_05736_ ), .Z(_05737_ ) );
BUF_X4 _13660_ ( .A(_05737_ ), .Z(_05738_ ) );
INV_X1 _13661_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_05739_ ) );
AOI211_X1 _13662_ ( .A(_05734_ ), .B(_05738_ ), .C1(_05739_ ), .C2(_01631_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _13663_ ( .A1(_05732_ ), .A2(fanout_net_6 ), .A3(_05733_ ), .ZN(_05740_ ) );
INV_X1 _13664_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_05741_ ) );
AOI211_X1 _13665_ ( .A(_05740_ ), .B(_05738_ ), .C1(_05741_ ), .C2(_01631_ ), .ZN(\io_master_araddr [0] ) );
OAI221_X1 _13666_ ( .A(\IF_ID_pc [15] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_05742_ ) );
INV_X1 _13667_ ( .A(_01538_ ), .ZN(_05743_ ) );
OR3_X1 _13668_ ( .A1(_05732_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(_05733_ ), .ZN(_05744_ ) );
BUF_X4 _13669_ ( .A(_01546_ ), .Z(_05745_ ) );
OAI211_X1 _13670_ ( .A(_05743_ ), .B(_05744_ ), .C1(\mylsu.araddr_tmp [15] ), .C2(_05745_ ), .ZN(_05746_ ) );
OAI21_X1 _13671_ ( .A(_05742_ ), .B1(\io_master_arburst [0] ), .B2(_05746_ ), .ZN(\io_master_araddr [15] ) );
OAI221_X1 _13672_ ( .A(\IF_ID_pc [14] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_05747_ ) );
OR3_X1 _13673_ ( .A1(_05732_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(_01543_ ), .ZN(_05748_ ) );
OAI211_X1 _13674_ ( .A(_05743_ ), .B(_05748_ ), .C1(\mylsu.araddr_tmp [14] ), .C2(_05745_ ), .ZN(_05749_ ) );
OAI21_X1 _13675_ ( .A(_05747_ ), .B1(\io_master_arburst [0] ), .B2(_05749_ ), .ZN(\io_master_araddr [14] ) );
NOR2_X1 _13676_ ( .A1(_05745_ ), .A2(\mylsu.araddr_tmp [5] ), .ZN(_05750_ ) );
NOR3_X1 _13677_ ( .A1(_05732_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(_01543_ ), .ZN(_05751_ ) );
NOR3_X1 _13678_ ( .A1(_01538_ ), .A2(_05750_ ), .A3(_05751_ ), .ZN(_05752_ ) );
MUX2_X1 _13679_ ( .A(_05752_ ), .B(\IF_ID_pc [5] ), .S(\io_master_arburst [0] ), .Z(\io_master_araddr [5] ) );
NOR3_X1 _13680_ ( .A1(_05732_ ), .A2(_02639_ ), .A3(_05733_ ), .ZN(_05753_ ) );
AOI21_X1 _13681_ ( .A(_05753_ ), .B1(_01631_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_05754_ ) );
BUF_X4 _13682_ ( .A(_01618_ ), .Z(_05755_ ) );
OAI22_X1 _13683_ ( .A1(_05738_ ), .A2(_05754_ ), .B1(_05623_ ), .B2(_05755_ ), .ZN(\io_master_araddr [4] ) );
NOR3_X1 _13684_ ( .A1(_05732_ ), .A2(_02654_ ), .A3(_05733_ ), .ZN(_05756_ ) );
AOI21_X1 _13685_ ( .A(_05756_ ), .B1(_01631_ ), .B2(\mylsu.araddr_tmp [3] ), .ZN(_05757_ ) );
OAI22_X1 _13686_ ( .A1(_05738_ ), .A2(_05757_ ), .B1(_05627_ ), .B2(_05755_ ), .ZN(\io_master_araddr [3] ) );
INV_X1 _13687_ ( .A(_01551_ ), .ZN(\io_master_araddr [31] ) );
INV_X1 _13688_ ( .A(_01607_ ), .ZN(\io_master_araddr [30] ) );
INV_X1 _13689_ ( .A(_01611_ ), .ZN(\io_master_araddr [29] ) );
INV_X1 _13690_ ( .A(_01563_ ), .ZN(\io_master_araddr [28] ) );
INV_X1 _13691_ ( .A(_01615_ ), .ZN(\io_master_araddr [27] ) );
INV_X1 _13692_ ( .A(_01567_ ), .ZN(\io_master_araddr [26] ) );
INV_X1 _13693_ ( .A(_01559_ ), .ZN(\io_master_araddr [24] ) );
NOR2_X1 _13694_ ( .A1(_05745_ ), .A2(\mylsu.araddr_tmp [13] ), .ZN(_05758_ ) );
NOR3_X1 _13695_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(_01543_ ), .ZN(_05759_ ) );
NOR3_X1 _13696_ ( .A1(_01538_ ), .A2(_05758_ ), .A3(_05759_ ), .ZN(_05760_ ) );
MUX2_X1 _13697_ ( .A(_05760_ ), .B(\IF_ID_pc [13] ), .S(\io_master_arburst [0] ), .Z(\io_master_araddr [13] ) );
INV_X1 _13698_ ( .A(_01590_ ), .ZN(\io_master_araddr [23] ) );
INV_X1 _13699_ ( .A(_01572_ ), .ZN(\io_master_araddr [22] ) );
INV_X1 _13700_ ( .A(_01580_ ), .ZN(\io_master_araddr [21] ) );
INV_X1 _13701_ ( .A(_01598_ ), .ZN(\io_master_araddr [20] ) );
INV_X1 _13702_ ( .A(_01584_ ), .ZN(\io_master_araddr [19] ) );
INV_X1 _13703_ ( .A(_01602_ ), .ZN(\io_master_araddr [18] ) );
INV_X1 _13704_ ( .A(_01594_ ), .ZN(\io_master_araddr [17] ) );
INV_X1 _13705_ ( .A(_01576_ ), .ZN(\io_master_araddr [16] ) );
OAI221_X1 _13706_ ( .A(\IF_ID_pc [12] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01548_ ), .C2(_01549_ ), .ZN(_05761_ ) );
OR3_X1 _13707_ ( .A1(_05732_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(_01543_ ), .ZN(_05762_ ) );
OAI211_X1 _13708_ ( .A(_05743_ ), .B(_05762_ ), .C1(\mylsu.araddr_tmp [12] ), .C2(_05745_ ), .ZN(_05763_ ) );
OAI21_X1 _13709_ ( .A(_05761_ ), .B1(\io_master_arburst [0] ), .B2(_05763_ ), .ZN(\io_master_araddr [12] ) );
NOR3_X1 _13710_ ( .A1(_05732_ ), .A2(_02644_ ), .A3(_05733_ ), .ZN(_05764_ ) );
AOI21_X1 _13711_ ( .A(_05764_ ), .B1(_01631_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_05765_ ) );
OAI22_X1 _13712_ ( .A1(_05738_ ), .A2(_05765_ ), .B1(_05438_ ), .B2(_05755_ ), .ZN(\io_master_araddr [11] ) );
AND2_X2 _13713_ ( .A1(EXU_valid_LSU ), .A2(\mylsu.state [0] ), .ZN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _13714_ ( .A1(_04996_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_02650_ ), .A4(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_05766_ ) );
OAI21_X1 _13715_ ( .A(_05766_ ), .B1(_05745_ ), .B2(\mylsu.araddr_tmp [10] ), .ZN(_05767_ ) );
OAI22_X1 _13716_ ( .A1(_05738_ ), .A2(_05767_ ), .B1(_01395_ ), .B2(_05755_ ), .ZN(\io_master_araddr [10] ) );
NAND4_X1 _13717_ ( .A1(_04996_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_05709_ ), .A4(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_05768_ ) );
OAI21_X1 _13718_ ( .A(_05768_ ), .B1(_05745_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_05769_ ) );
OAI22_X1 _13719_ ( .A1(_05738_ ), .A2(_05769_ ), .B1(_05442_ ), .B2(_05755_ ), .ZN(\io_master_araddr [9] ) );
NAND4_X1 _13720_ ( .A1(_04996_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_05710_ ), .A4(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_05770_ ) );
OAI21_X1 _13721_ ( .A(_05770_ ), .B1(_05745_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_05771_ ) );
OAI22_X1 _13722_ ( .A1(_05738_ ), .A2(_05771_ ), .B1(_05212_ ), .B2(_05755_ ), .ZN(\io_master_araddr [8] ) );
OR3_X1 _13723_ ( .A1(_05732_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(_05733_ ), .ZN(_05772_ ) );
OAI21_X1 _13724_ ( .A(_05772_ ), .B1(_05745_ ), .B2(\mylsu.araddr_tmp [7] ), .ZN(_05773_ ) );
OAI22_X1 _13725_ ( .A1(_05738_ ), .A2(_05773_ ), .B1(_01363_ ), .B2(_05755_ ), .ZN(\io_master_araddr [7] ) );
NAND4_X1 _13726_ ( .A1(_04996_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_05711_ ), .A4(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ), .ZN(_05774_ ) );
OAI21_X1 _13727_ ( .A(_05774_ ), .B1(_05745_ ), .B2(\mylsu.araddr_tmp [6] ), .ZN(_05775_ ) );
OAI22_X1 _13728_ ( .A1(_05738_ ), .A2(_05775_ ), .B1(_01498_ ), .B2(_05755_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _13729_ ( .A1(_01542_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(_01543_ ), .ZN(_05776_ ) );
OAI211_X1 _13730_ ( .A(_05743_ ), .B(_05776_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01546_ ), .ZN(_05777_ ) );
NOR2_X1 _13731_ ( .A1(_01533_ ), .A2(_05777_ ), .ZN(_05778_ ) );
BUF_X4 _13732_ ( .A(_05778_ ), .Z(_05779_ ) );
BUF_X2 _13733_ ( .A(_05779_ ), .Z(\io_master_araddr [2] ) );
INV_X1 _13734_ ( .A(\EX_LS_typ [3] ), .ZN(_05780_ ) );
NOR3_X1 _13735_ ( .A1(\io_master_arburst [0] ), .A2(_05780_ ), .A3(_01538_ ), .ZN(\io_master_arsize [2] ) );
INV_X1 _13736_ ( .A(\EX_LS_typ [1] ), .ZN(_05781_ ) );
NOR3_X1 _13737_ ( .A1(\io_master_arburst [0] ), .A2(_05781_ ), .A3(_01538_ ), .ZN(\io_master_arsize [0] ) );
INV_X1 _13738_ ( .A(\EX_LS_typ [2] ), .ZN(_05782_ ) );
OAI22_X1 _13739_ ( .A1(_01531_ ), .A2(_01532_ ), .B1(_05782_ ), .B2(_01538_ ), .ZN(\io_master_arsize [1] ) );
INV_X1 _13740_ ( .A(_04994_ ), .ZN(_05783_ ) );
AND3_X1 _13741_ ( .A1(_05783_ ), .A2(_01632_ ), .A3(_01635_ ), .ZN(io_master_arvalid ) );
AND2_X1 _13742_ ( .A1(_04999_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_05784_ ) );
BUF_X4 _13743_ ( .A(_05784_ ), .Z(_05785_ ) );
BUF_X4 _13744_ ( .A(_05785_ ), .Z(_05786_ ) );
MUX2_X1 _13745_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_05786_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _13746_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_05786_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _13747_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_05786_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _13748_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_05786_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _13749_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_05786_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _13750_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_05786_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _13751_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_05786_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _13752_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_05786_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _13753_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_05786_ ), .Z(\io_master_awaddr [15] ) );
BUF_X4 _13754_ ( .A(_05785_ ), .Z(_05787_ ) );
MUX2_X1 _13755_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_05787_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _13756_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_05787_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _13757_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_05787_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _13758_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_05787_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _13759_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_05787_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _13760_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_05787_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _13761_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_05787_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _13762_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_05787_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _13763_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_05787_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _13764_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_05787_ ), .Z(\io_master_awaddr [6] ) );
BUF_X4 _13765_ ( .A(_05785_ ), .Z(_05788_ ) );
MUX2_X1 _13766_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_05788_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _13767_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_05788_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _13768_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_05788_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _13769_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_05788_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _13770_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_05788_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _13771_ ( .A(\mylsu.awaddr_tmp [1] ), .B(fanout_net_7 ), .S(_05788_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _13772_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_6 ), .S(_05788_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _13773_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_05788_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _13774_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_05788_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _13775_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_05788_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _13776_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_05785_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _13777_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_05785_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _13778_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_05785_ ), .Z(\io_master_awaddr [22] ) );
INV_X1 _13779_ ( .A(_05786_ ), .ZN(_05789_ ) );
INV_X1 _13780_ ( .A(io_master_wready ), .ZN(_05790_ ) );
AOI211_X1 _13781_ ( .A(fanout_net_5 ), .B(_05789_ ), .C1(_05000_ ), .C2(_05790_ ), .ZN(io_master_awready_$_NOR__A_Y_$_OR__A_Y_$_OR__B_Y_$_ANDNOT__B_Y ) );
INV_X1 _13782_ ( .A(\EX_LS_typ [0] ), .ZN(_05791_ ) );
NOR4_X1 _13783_ ( .A1(_05791_ ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .A4(\EX_LS_typ [4] ), .ZN(_05792_ ) );
AND3_X1 _13784_ ( .A1(_05792_ ), .A2(_04999_ ), .A3(\EX_LS_typ [1] ), .ZN(\io_master_awsize [0] ) );
NAND4_X1 _13785_ ( .A1(_05792_ ), .A2(_01675_ ), .A3(\EX_LS_flag [1] ), .A4(_01673_ ), .ZN(\io_master_awsize [1] ) );
INV_X1 _13786_ ( .A(_04999_ ), .ZN(_05793_ ) );
INV_X1 _13787_ ( .A(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_05794_ ) );
OAI21_X1 _13788_ ( .A(_05004_ ), .B1(_05793_ ), .B2(_05794_ ), .ZN(io_master_awvalid ) );
INV_X1 _13789_ ( .A(\mylsu.state [2] ), .ZN(_05795_ ) );
INV_X1 _13790_ ( .A(\mylsu.state [1] ), .ZN(_05796_ ) );
NAND4_X1 _13791_ ( .A1(_05789_ ), .A2(_05795_ ), .A3(_05004_ ), .A4(_05796_ ), .ZN(io_master_bready ) );
NOR2_X1 _13792_ ( .A1(_05681_ ), .A2(\io_master_rid [0] ), .ZN(_05797_ ) );
NAND4_X1 _13793_ ( .A1(_05797_ ), .A2(io_master_rlast ), .A3(_05679_ ), .A4(_05680_ ), .ZN(_05798_ ) );
AOI21_X1 _13794_ ( .A(_05736_ ), .B1(_05678_ ), .B2(_05798_ ), .ZN(_05799_ ) );
AND2_X1 _13795_ ( .A1(_05799_ ), .A2(_05692_ ), .ZN(_05800_ ) );
BUF_X4 _13796_ ( .A(_05702_ ), .Z(_05801_ ) );
NOR2_X1 _13797_ ( .A1(_05800_ ), .A2(_05801_ ), .ZN(_05802_ ) );
NOR2_X1 _13798_ ( .A1(\io_master_bid [3] ), .A2(\io_master_bid [2] ), .ZN(_05803_ ) );
NAND3_X1 _13799_ ( .A1(_05803_ ), .A2(\io_master_bid [1] ), .A3(\io_master_bid [0] ), .ZN(_05804_ ) );
NOR2_X1 _13800_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_05805_ ) );
NAND2_X1 _13801_ ( .A1(_05805_ ), .A2(io_master_bvalid ), .ZN(_05806_ ) );
NOR2_X1 _13802_ ( .A1(_05804_ ), .A2(_05806_ ), .ZN(_05807_ ) );
NOR2_X1 _13803_ ( .A1(_05807_ ), .A2(_05796_ ), .ZN(_05808_ ) );
NOR3_X1 _13804_ ( .A1(_01537_ ), .A2(\mylsu.state [0] ), .A3(\mylsu.state [1] ), .ZN(_05809_ ) );
NOR3_X1 _13805_ ( .A1(_05802_ ), .A2(_05808_ ), .A3(_05809_ ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__B_Y_$_NOR__A_Y ) );
AOI21_X1 _13806_ ( .A(_01628_ ), .B1(_01586_ ), .B2(_01620_ ), .ZN(io_master_rready ) );
MUX2_X1 _13807_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_6 ), .Z(_05810_ ) );
CLKBUF_X2 _13808_ ( .A(_02647_ ), .Z(_05811_ ) );
AND2_X1 _13809_ ( .A1(_05810_ ), .A2(_05811_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _13810_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_6 ), .Z(_05812_ ) );
AND2_X1 _13811_ ( .A1(_05812_ ), .A2(_05811_ ), .ZN(\io_master_wdata [14] ) );
NOR3_X1 _13812_ ( .A1(_04634_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _13813_ ( .A1(_04668_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [4] ) );
NOR3_X1 _13814_ ( .A1(_04697_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [3] ) );
NOR3_X1 _13815_ ( .A1(_04734_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [2] ) );
NOR3_X1 _13816_ ( .A1(_04754_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [1] ) );
NOR3_X1 _13817_ ( .A1(_04808_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _13818_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_6 ), .Z(_05813_ ) );
AND2_X1 _13819_ ( .A1(_05813_ ), .A2(_05811_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _13820_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_6 ), .Z(_05814_ ) );
AND2_X1 _13821_ ( .A1(_05814_ ), .A2(_05811_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _13822_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_6 ), .Z(_05815_ ) );
AND2_X1 _13823_ ( .A1(_05815_ ), .A2(_05811_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _13824_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_6 ), .Z(_05816_ ) );
AND2_X1 _13825_ ( .A1(_05816_ ), .A2(_05811_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _13826_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_6 ), .Z(_05817_ ) );
AND2_X1 _13827_ ( .A1(_05817_ ), .A2(_05811_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _13828_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_6 ), .Z(_05818_ ) );
AND2_X1 _13829_ ( .A1(_05818_ ), .A2(_05811_ ), .ZN(\io_master_wdata [8] ) );
NOR3_X1 _13830_ ( .A1(_04582_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [7] ) );
NOR3_X1 _13831_ ( .A1(_04604_ ), .A2(fanout_net_7 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _13832_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_6 ), .Z(_05819_ ) );
MUX2_X1 _13833_ ( .A(_05819_ ), .B(_05810_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _13834_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_6 ), .Z(_05820_ ) );
MUX2_X1 _13835_ ( .A(_05820_ ), .B(_05812_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [30] ) );
NAND3_X1 _13836_ ( .A1(_05712_ ), .A2(fanout_net_7 ), .A3(\EX_LS_result_csreg_mem [5] ), .ZN(_05821_ ) );
MUX2_X1 _13837_ ( .A(_04940_ ), .B(_04368_ ), .S(fanout_net_6 ), .Z(_05822_ ) );
OAI21_X1 _13838_ ( .A(_05821_ ), .B1(_05822_ ), .B2(fanout_net_7 ), .ZN(\io_master_wdata [21] ) );
NAND3_X1 _13839_ ( .A1(_05712_ ), .A2(fanout_net_7 ), .A3(\EX_LS_result_csreg_mem [4] ), .ZN(_05823_ ) );
MUX2_X1 _13840_ ( .A(_04182_ ), .B(_04415_ ), .S(fanout_net_6 ), .Z(_05824_ ) );
OAI21_X1 _13841_ ( .A(_05823_ ), .B1(_05824_ ), .B2(fanout_net_7 ), .ZN(\io_master_wdata [20] ) );
NOR2_X1 _13842_ ( .A1(_04697_ ), .A2(fanout_net_6 ), .ZN(_05825_ ) );
MUX2_X1 _13843_ ( .A(\EX_LS_result_csreg_mem [19] ), .B(\EX_LS_result_csreg_mem [11] ), .S(fanout_net_6 ), .Z(_05826_ ) );
MUX2_X1 _13844_ ( .A(_05825_ ), .B(_05826_ ), .S(_05811_ ), .Z(\io_master_wdata [19] ) );
NOR2_X1 _13845_ ( .A1(_04734_ ), .A2(fanout_net_6 ), .ZN(_05827_ ) );
MUX2_X1 _13846_ ( .A(\EX_LS_result_csreg_mem [18] ), .B(\EX_LS_result_csreg_mem [10] ), .S(fanout_net_6 ), .Z(_05828_ ) );
MUX2_X1 _13847_ ( .A(_05827_ ), .B(_05828_ ), .S(_02647_ ), .Z(\io_master_wdata [18] ) );
NOR2_X1 _13848_ ( .A1(_04754_ ), .A2(fanout_net_6 ), .ZN(_05829_ ) );
MUX2_X1 _13849_ ( .A(\EX_LS_result_csreg_mem [17] ), .B(\EX_LS_result_csreg_mem [9] ), .S(fanout_net_6 ), .Z(_05830_ ) );
MUX2_X1 _13850_ ( .A(_05829_ ), .B(_05830_ ), .S(_02647_ ), .Z(\io_master_wdata [17] ) );
NOR2_X1 _13851_ ( .A1(_04808_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .ZN(_05831_ ) );
MUX2_X1 _13852_ ( .A(\EX_LS_result_csreg_mem [16] ), .B(\EX_LS_result_csreg_mem [8] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05832_ ) );
MUX2_X1 _13853_ ( .A(_05831_ ), .B(_05832_ ), .S(_02647_ ), .Z(\io_master_wdata [16] ) );
MUX2_X1 _13854_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05833_ ) );
MUX2_X1 _13855_ ( .A(_05833_ ), .B(_05813_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _13856_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05834_ ) );
MUX2_X1 _13857_ ( .A(_05834_ ), .B(_05814_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _13858_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05835_ ) );
MUX2_X1 _13859_ ( .A(_05835_ ), .B(_05815_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _13860_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05836_ ) );
MUX2_X1 _13861_ ( .A(_05836_ ), .B(_05816_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _13862_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05837_ ) );
MUX2_X1 _13863_ ( .A(_05837_ ), .B(_05817_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _13864_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05838_ ) );
MUX2_X1 _13865_ ( .A(_05838_ ), .B(_05818_ ), .S(fanout_net_7 ), .Z(\io_master_wdata [24] ) );
NOR2_X1 _13866_ ( .A1(_04582_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .ZN(_05839_ ) );
MUX2_X1 _13867_ ( .A(\EX_LS_result_csreg_mem [23] ), .B(\EX_LS_result_csreg_mem [15] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05840_ ) );
MUX2_X1 _13868_ ( .A(_05839_ ), .B(_05840_ ), .S(_02647_ ), .Z(\io_master_wdata [23] ) );
NOR2_X1 _13869_ ( .A1(_04604_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .ZN(_05841_ ) );
MUX2_X1 _13870_ ( .A(\EX_LS_result_csreg_mem [22] ), .B(\EX_LS_result_csreg_mem [14] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05842_ ) );
MUX2_X1 _13871_ ( .A(_05841_ ), .B(_05842_ ), .S(_02647_ ), .Z(\io_master_wdata [22] ) );
MUX2_X1 _13872_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05843_ ) );
AND2_X1 _13873_ ( .A1(_05843_ ), .A2(_05811_ ), .ZN(\io_master_wstrb [1] ) );
NOR3_X1 _13874_ ( .A1(_05791_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _13875_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05844_ ) );
MUX2_X1 _13876_ ( .A(_05844_ ), .B(_05843_ ), .S(fanout_net_7 ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _13877_ ( .A1(_05712_ ), .A2(fanout_net_7 ), .A3(\EX_LS_typ [0] ), .ZN(_05845_ ) );
MUX2_X1 _13878_ ( .A(_05782_ ), .B(_05781_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_05846_ ) );
OAI21_X1 _13879_ ( .A(_05845_ ), .B1(_05846_ ), .B2(fanout_net_7 ), .ZN(\io_master_wstrb [2] ) );
OAI21_X1 _13880_ ( .A(_05795_ ), .B1(_05793_ ), .B2(_05794_ ), .ZN(io_master_wvalid ) );
NOR2_X1 _13881_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_05847_ ) );
AND2_X1 _13882_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_05848_ ) );
NOR2_X1 _13883_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_05849_ ) );
NOR2_X1 _13884_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_05850_ ) );
AND4_X1 _13885_ ( .A1(_05847_ ), .A2(_05848_ ), .A3(_05849_ ), .A4(_05850_ ), .ZN(_05851_ ) );
AND2_X1 _13886_ ( .A1(_01051_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(_05852_ ) );
INV_X1 _13887_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_05853_ ) );
NOR3_X1 _13888_ ( .A1(_05853_ ), .A2(\LS_WB_waddr_csreg [1] ), .A3(\LS_WB_waddr_csreg [3] ), .ZN(_05854_ ) );
AND4_X1 _13889_ ( .A1(\LS_WB_waddr_csreg [2] ), .A2(_05851_ ), .A3(_05852_ ), .A4(_05854_ ), .ZN(\mycsreg.CSReg[1]_$_DFFE_PP__Q_E ) );
INV_X1 _13890_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_05855_ ) );
AND3_X1 _13891_ ( .A1(_05852_ ), .A2(_05848_ ), .A3(_05850_ ), .ZN(_05856_ ) );
NOR3_X1 _13892_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .A3(\LS_WB_waddr_csreg [7] ), .ZN(_05857_ ) );
AND3_X1 _13893_ ( .A1(_05857_ ), .A2(\LS_WB_waddr_csreg [6] ), .A3(_05847_ ), .ZN(_05858_ ) );
AND4_X1 _13894_ ( .A1(_05855_ ), .A2(_05856_ ), .A3(\LS_WB_waddr_csreg [0] ), .A4(_05858_ ), .ZN(\mycsreg.CSReg[2]_$_DFFE_PP__Q_E ) );
OR2_X1 _13895_ ( .A1(\LS_WB_wen_csreg [1] ), .A2(\LS_WB_wdata_csreg [1] ), .ZN(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _13896_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [1] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _13897_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [1] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
NAND2_X1 _13898_ ( .A1(_04765_ ), .A2(_02579_ ), .ZN(_05859_ ) );
INV_X1 _13899_ ( .A(_02576_ ), .ZN(_05860_ ) );
BUF_X4 _13900_ ( .A(_05860_ ), .Z(_05861_ ) );
BUF_X4 _13901_ ( .A(_05861_ ), .Z(_05862_ ) );
OAI21_X1 _13902_ ( .A(_05859_ ), .B1(_02642_ ), .B2(_05862_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _13903_ ( .A(_03645_ ), .B(\ID_EX_imm [0] ), .ZN(_05863_ ) );
BUF_X4 _13904_ ( .A(_02576_ ), .Z(_05864_ ) );
BUF_X4 _13905_ ( .A(_05864_ ), .Z(_05865_ ) );
AOI22_X1 _13906_ ( .A1(_05863_ ), .A2(_02584_ ), .B1(_02670_ ), .B2(_05865_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND2_X1 _13907_ ( .A1(_04514_ ), .A2(_04812_ ), .ZN(_05866_ ) );
BUF_X4 _13908_ ( .A(_05860_ ), .Z(_05867_ ) );
MUX2_X1 _13909_ ( .A(\ID_EX_csr [10] ), .B(_05866_ ), .S(_05867_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
NOR4_X1 _13910_ ( .A1(_01656_ ), .A2(_01659_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [9] ), .ZN(_05868_ ) );
AOI21_X1 _13911_ ( .A(_05868_ ), .B1(_04538_ ), .B2(_02584_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
NOR2_X1 _13912_ ( .A1(_04563_ ), .A2(_02580_ ), .ZN(_05869_ ) );
BUF_X4 _13913_ ( .A(_02576_ ), .Z(_05870_ ) );
BUF_X4 _13914_ ( .A(_05870_ ), .Z(_05871_ ) );
AOI21_X1 _13915_ ( .A(_05869_ ), .B1(_02640_ ), .B2(_05871_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND4_X1 _13916_ ( .A1(_01647_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_csr [7] ), .ZN(_05872_ ) );
OAI21_X1 _13917_ ( .A(_05872_ ), .B1(_04594_ ), .B2(_02581_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
NOR2_X1 _13918_ ( .A1(_04625_ ), .A2(_02580_ ), .ZN(_05873_ ) );
AOI21_X1 _13919_ ( .A(_05873_ ), .B1(_02692_ ), .B2(_05871_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND4_X1 _13920_ ( .A1(_01647_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_csr [5] ), .ZN(_05874_ ) );
OAI21_X1 _13921_ ( .A(_05874_ ), .B1(_04658_ ), .B2(_02581_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _13922_ ( .A1(_04688_ ), .A2(_02579_ ), .ZN(_05875_ ) );
OAI21_X1 _13923_ ( .A(_05875_ ), .B1(_02679_ ), .B2(_05862_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _13924_ ( .A1(_04718_ ), .A2(_02579_ ), .ZN(_05876_ ) );
OAI21_X1 _13925_ ( .A(_05876_ ), .B1(_02658_ ), .B2(_05862_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _13926_ ( .A1(_04739_ ), .A2(_02579_ ), .ZN(_05877_ ) );
OAI21_X1 _13927_ ( .A(_05877_ ), .B1(_02645_ ), .B2(_05862_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
NAND2_X1 _13928_ ( .A1(_04460_ ), .A2(_02579_ ), .ZN(_05878_ ) );
OAI21_X1 _13929_ ( .A(_05878_ ), .B1(_02657_ ), .B2(_05862_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X4 _13930_ ( .A(_05864_ ), .Z(_05879_ ) );
AND3_X1 _13931_ ( .A1(_01841_ ), .A2(_04227_ ), .A3(_01842_ ), .ZN(_05880_ ) );
NOR2_X1 _13932_ ( .A1(_04976_ ), .A2(\ID_EX_imm [21] ), .ZN(_05881_ ) );
NOR2_X1 _13933_ ( .A1(_05880_ ), .A2(_05881_ ), .ZN(_05882_ ) );
NOR2_X1 _13934_ ( .A1(_04073_ ), .A2(\ID_EX_typ [2] ), .ZN(_05883_ ) );
INV_X1 _13935_ ( .A(_05883_ ), .ZN(_05884_ ) );
BUF_X4 _13936_ ( .A(_05884_ ), .Z(_05885_ ) );
NOR3_X1 _13937_ ( .A1(_04939_ ), .A2(_05885_ ), .A3(_04941_ ), .ZN(_05886_ ) );
OAI221_X1 _13938_ ( .A(_05879_ ), .B1(_04942_ ), .B2(_05008_ ), .C1(_05882_ ), .C2(_05886_ ), .ZN(_05887_ ) );
BUF_X4 _13939_ ( .A(_05861_ ), .Z(_05888_ ) );
NAND4_X1 _13940_ ( .A1(_04946_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_05889_ ) );
OAI211_X1 _13941_ ( .A(_05888_ ), .B(_05889_ ), .C1(_04063_ ), .C2(_04163_ ), .ZN(_05890_ ) );
NAND2_X1 _13942_ ( .A1(_05887_ ), .A2(_05890_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
CLKBUF_X2 _13943_ ( .A(_05860_ ), .Z(_05891_ ) );
NAND2_X1 _13944_ ( .A1(_01870_ ), .A2(fanout_net_8 ), .ZN(_05892_ ) );
OAI221_X1 _13945_ ( .A(_05892_ ), .B1(fanout_net_8 ), .B2(_01869_ ), .C1(_04185_ ), .C2(_05008_ ), .ZN(_05893_ ) );
BUF_X4 _13946_ ( .A(_05883_ ), .Z(_05894_ ) );
NAND3_X1 _13947_ ( .A1(_04179_ ), .A2(_05894_ ), .A3(_04184_ ), .ZN(_05895_ ) );
AOI21_X1 _13948_ ( .A(_05891_ ), .B1(_05893_ ), .B2(_05895_ ), .ZN(_05896_ ) );
AND3_X1 _13949_ ( .A1(_01646_ ), .A2(_04944_ ), .A3(\ID_EX_typ [7] ), .ZN(_05897_ ) );
BUF_X4 _13950_ ( .A(_02838_ ), .Z(_05898_ ) );
AOI211_X1 _13951_ ( .A(_05864_ ), .B(_05897_ ), .C1(_03083_ ), .C2(_05898_ ), .ZN(_05899_ ) );
OR2_X1 _13952_ ( .A1(_05896_ ), .A2(_05899_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
CLKBUF_X2 _13953_ ( .A(_01646_ ), .Z(_05900_ ) );
NAND3_X1 _13954_ ( .A1(_05900_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_typ [7] ), .ZN(_05901_ ) );
OAI21_X1 _13955_ ( .A(_05901_ ), .B1(_02976_ ), .B2(_04125_ ), .ZN(_05902_ ) );
AOI21_X1 _13956_ ( .A(_05884_ ), .B1(_04209_ ), .B2(_04222_ ), .ZN(_05903_ ) );
AOI21_X1 _13957_ ( .A(fanout_net_8 ), .B1(_01916_ ), .B2(_01917_ ), .ZN(_05904_ ) );
AND2_X1 _13958_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [19] ), .ZN(_05905_ ) );
NOR3_X1 _13959_ ( .A1(_05903_ ), .A2(_05904_ ), .A3(_05905_ ), .ZN(_05906_ ) );
AOI21_X1 _13960_ ( .A(_05906_ ), .B1(\ID_EX_typ [2] ), .B2(_04211_ ), .ZN(_05907_ ) );
MUX2_X1 _13961_ ( .A(_05902_ ), .B(_05907_ ), .S(_05864_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
AOI22_X1 _13962_ ( .A1(_04240_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_8 ), .B2(_01896_ ), .ZN(_05908_ ) );
BUF_X4 _13963_ ( .A(_02576_ ), .Z(_05909_ ) );
OAI211_X1 _13964_ ( .A(_05908_ ), .B(_05909_ ), .C1(fanout_net_8 ), .C2(_01895_ ), .ZN(_05910_ ) );
AOI21_X1 _13965_ ( .A(_05860_ ), .B1(_04238_ ), .B2(_04248_ ), .ZN(_05911_ ) );
BUF_X4 _13966_ ( .A(_05894_ ), .Z(_05912_ ) );
NAND2_X1 _13967_ ( .A1(_05911_ ), .A2(_05912_ ), .ZN(_05913_ ) );
MUX2_X1 _13968_ ( .A(_04241_ ), .B(_03004_ ), .S(_04812_ ), .Z(_05914_ ) );
OAI211_X1 _13969_ ( .A(_05910_ ), .B(_05913_ ), .C1(_05871_ ), .C2(_05914_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
AOI22_X1 _13970_ ( .A1(_04267_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_8 ), .B2(_01943_ ), .ZN(_05915_ ) );
BUF_X4 _13971_ ( .A(_05864_ ), .Z(_05916_ ) );
OAI211_X1 _13972_ ( .A(_05915_ ), .B(_05916_ ), .C1(fanout_net_9 ), .C2(_01942_ ), .ZN(_05917_ ) );
AND3_X1 _13973_ ( .A1(_04260_ ), .A2(_05864_ ), .A3(_04265_ ), .ZN(_05918_ ) );
NAND2_X1 _13974_ ( .A1(_05918_ ), .A2(_05912_ ), .ZN(_05919_ ) );
AOI21_X1 _13975_ ( .A(_04125_ ), .B1(_02913_ ), .B2(_02920_ ), .ZN(_05920_ ) );
AND3_X1 _13976_ ( .A1(_05900_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_typ [7] ), .ZN(_05921_ ) );
OAI21_X1 _13977_ ( .A(_05888_ ), .B1(_05920_ ), .B2(_05921_ ), .ZN(_05922_ ) );
NAND3_X1 _13978_ ( .A1(_05917_ ), .A2(_05919_ ), .A3(_05922_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
AOI22_X1 _13979_ ( .A1(_04295_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_01966_ ), .ZN(_05923_ ) );
OAI211_X1 _13980_ ( .A(_05923_ ), .B(_05909_ ), .C1(fanout_net_9 ), .C2(_01965_ ), .ZN(_05924_ ) );
AND3_X1 _13981_ ( .A1(_04292_ ), .A2(_02576_ ), .A3(_04293_ ), .ZN(_05925_ ) );
NAND2_X1 _13982_ ( .A1(_05925_ ), .A2(_05912_ ), .ZN(_05926_ ) );
MUX2_X1 _13983_ ( .A(_04272_ ), .B(_02952_ ), .S(_04812_ ), .Z(_05927_ ) );
OAI211_X1 _13984_ ( .A(_05924_ ), .B(_05926_ ), .C1(_05871_ ), .C2(_05927_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
AOI22_X1 _13985_ ( .A1(_04315_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02310_ ), .ZN(_05928_ ) );
OAI211_X1 _13986_ ( .A(_05928_ ), .B(_05870_ ), .C1(fanout_net_9 ), .C2(_02309_ ), .ZN(_05929_ ) );
AOI21_X1 _13987_ ( .A(_05860_ ), .B1(_04313_ ), .B2(_04325_ ), .ZN(_05930_ ) );
NAND2_X1 _13988_ ( .A1(_05930_ ), .A2(_05912_ ), .ZN(_05931_ ) );
MUX2_X1 _13989_ ( .A(_04991_ ), .B(_03162_ ), .S(_04812_ ), .Z(_05932_ ) );
OAI211_X1 _13990_ ( .A(_05929_ ), .B(_05931_ ), .C1(_05871_ ), .C2(_05932_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
AOI22_X1 _13991_ ( .A1(_04346_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02333_ ), .ZN(_05933_ ) );
OAI211_X1 _13992_ ( .A(_05933_ ), .B(_05870_ ), .C1(fanout_net_9 ), .C2(_02332_ ), .ZN(_05934_ ) );
AND3_X1 _13993_ ( .A1(_04343_ ), .A2(_02576_ ), .A3(_04344_ ), .ZN(_05935_ ) );
NAND2_X1 _13994_ ( .A1(_05935_ ), .A2(_05912_ ), .ZN(_05936_ ) );
MUX2_X1 _13995_ ( .A(_04347_ ), .B(_03134_ ), .S(_04812_ ), .Z(_05937_ ) );
OAI211_X1 _13996_ ( .A(_05934_ ), .B(_05936_ ), .C1(_05865_ ), .C2(_05937_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OAI21_X1 _13997_ ( .A(\ID_EX_typ [2] ), .B1(_04367_ ), .B2(_04369_ ), .ZN(_05938_ ) );
NAND2_X1 _13998_ ( .A1(_02355_ ), .A2(fanout_net_9 ), .ZN(_05939_ ) );
NAND3_X1 _13999_ ( .A1(_02354_ ), .A2(_04227_ ), .A3(_02356_ ), .ZN(_05940_ ) );
NAND3_X1 _14000_ ( .A1(_05938_ ), .A2(_05939_ ), .A3(_05940_ ), .ZN(_05941_ ) );
OR3_X1 _14001_ ( .A1(_04367_ ), .A2(_05884_ ), .A3(_04369_ ), .ZN(_05942_ ) );
NAND3_X1 _14002_ ( .A1(_05941_ ), .A2(_05864_ ), .A3(_05942_ ), .ZN(_05943_ ) );
INV_X1 _14003_ ( .A(_05943_ ), .ZN(_05944_ ) );
MUX2_X1 _14004_ ( .A(_04374_ ), .B(_03212_ ), .S(_04812_ ), .Z(_05945_ ) );
AOI21_X1 _14005_ ( .A(_05944_ ), .B1(_05862_ ), .B2(_05945_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AOI22_X1 _14006_ ( .A1(_04418_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02381_ ), .ZN(_05946_ ) );
OAI211_X1 _14007_ ( .A(_05946_ ), .B(_05916_ ), .C1(fanout_net_9 ), .C2(_02380_ ), .ZN(_05947_ ) );
AND3_X1 _14008_ ( .A1(_04414_ ), .A2(_05864_ ), .A3(_04416_ ), .ZN(_05948_ ) );
NAND2_X1 _14009_ ( .A1(_05948_ ), .A2(_05912_ ), .ZN(_05949_ ) );
AOI21_X1 _14010_ ( .A(_04125_ ), .B1(_03166_ ), .B2(_03186_ ), .ZN(_05950_ ) );
AND3_X1 _14011_ ( .A1(_05900_ ), .A2(\ID_EX_pc [12] ), .A3(\ID_EX_typ [7] ), .ZN(_05951_ ) );
OAI21_X1 _14012_ ( .A(_05888_ ), .B1(_05950_ ), .B2(_05951_ ), .ZN(_05952_ ) );
NAND3_X1 _14013_ ( .A1(_05947_ ), .A2(_05949_ ), .A3(_05952_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _14014_ ( .A(_05885_ ), .B1(_02713_ ), .B2(_02718_ ), .ZN(_05953_ ) );
AOI22_X1 _14015_ ( .A1(_02719_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_01733_ ), .ZN(_05954_ ) );
NAND3_X1 _14016_ ( .A1(_01724_ ), .A2(_04976_ ), .A3(_01731_ ), .ZN(_05955_ ) );
AOI211_X1 _14017_ ( .A(_05891_ ), .B(_05953_ ), .C1(_05954_ ), .C2(_05955_ ), .ZN(_05956_ ) );
NAND3_X1 _14018_ ( .A1(_05900_ ), .A2(_04984_ ), .A3(\ID_EX_typ [7] ), .ZN(_05957_ ) );
OAI21_X1 _14019_ ( .A(_05957_ ), .B1(_03549_ ), .B2(_04163_ ), .ZN(_05958_ ) );
AOI21_X1 _14020_ ( .A(_05956_ ), .B1(_05862_ ), .B2(_05958_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _14021_ ( .A1(_02715_ ), .A2(_04437_ ), .A3(_02717_ ), .ZN(_05959_ ) );
NAND4_X1 _14022_ ( .A1(_04436_ ), .A2(_05870_ ), .A3(_05894_ ), .A4(_05959_ ), .ZN(_05960_ ) );
MUX2_X1 _14023_ ( .A(_04442_ ), .B(_03240_ ), .S(_02838_ ), .Z(_05961_ ) );
OAI221_X1 _14024_ ( .A(_05870_ ), .B1(_05009_ ), .B2(\ID_EX_imm [11] ), .C1(_04439_ ), .C2(_05008_ ), .ZN(_05962_ ) );
AND3_X1 _14025_ ( .A1(_02270_ ), .A2(_05009_ ), .A3(_02271_ ), .ZN(_05963_ ) );
OAI221_X1 _14026_ ( .A(_05960_ ), .B1(_05865_ ), .B2(_05961_ ), .C1(_05962_ ), .C2(_05963_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI22_X1 _14027_ ( .A1(_04498_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02250_ ), .ZN(_05964_ ) );
NAND3_X1 _14028_ ( .A1(_02247_ ), .A2(_04227_ ), .A3(_02248_ ), .ZN(_05965_ ) );
AND2_X1 _14029_ ( .A1(_05964_ ), .A2(_05965_ ), .ZN(_05966_ ) );
AOI21_X1 _14030_ ( .A(_05885_ ), .B1(_04496_ ), .B2(_04509_ ), .ZN(_05967_ ) );
OAI21_X1 _14031_ ( .A(_05879_ ), .B1(_05966_ ), .B2(_05967_ ), .ZN(_05968_ ) );
MUX2_X1 _14032_ ( .A(_04500_ ), .B(_03265_ ), .S(_04812_ ), .Z(_05969_ ) );
OAI21_X1 _14033_ ( .A(_05968_ ), .B1(_05871_ ), .B2(_05969_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
AOI22_X1 _14034_ ( .A1(_04526_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02226_ ), .ZN(_05970_ ) );
OAI211_X1 _14035_ ( .A(_05970_ ), .B(_05916_ ), .C1(fanout_net_9 ), .C2(_02225_ ), .ZN(_05971_ ) );
AOI21_X1 _14036_ ( .A(_05891_ ), .B1(_04524_ ), .B2(_04525_ ), .ZN(_05972_ ) );
NAND2_X1 _14037_ ( .A1(_05972_ ), .A2(_05912_ ), .ZN(_05973_ ) );
AOI21_X1 _14038_ ( .A(_04125_ ), .B1(_03270_ ), .B2(_03290_ ), .ZN(_05974_ ) );
AND3_X1 _14039_ ( .A1(_05900_ ), .A2(\ID_EX_pc [9] ), .A3(\ID_EX_typ [7] ), .ZN(_05975_ ) );
OAI21_X1 _14040_ ( .A(_05888_ ), .B1(_05974_ ), .B2(_05975_ ), .ZN(_05976_ ) );
NAND3_X1 _14041_ ( .A1(_05971_ ), .A2(_05973_ ), .A3(_05976_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _14042_ ( .A1(_02715_ ), .A2(_04549_ ), .A3(_02717_ ), .ZN(_05977_ ) );
NAND4_X1 _14043_ ( .A1(_04548_ ), .A2(_05870_ ), .A3(_05894_ ), .A4(_05977_ ), .ZN(_05978_ ) );
MUX2_X1 _14044_ ( .A(_04553_ ), .B(_03316_ ), .S(_02838_ ), .Z(_05979_ ) );
OAI221_X1 _14045_ ( .A(_05864_ ), .B1(_05009_ ), .B2(\ID_EX_imm [8] ), .C1(_04551_ ), .C2(_05008_ ), .ZN(_05980_ ) );
AND3_X1 _14046_ ( .A1(_02200_ ), .A2(_05009_ ), .A3(_02201_ ), .ZN(_05981_ ) );
OAI221_X1 _14047_ ( .A(_05978_ ), .B1(_05979_ ), .B2(_05879_ ), .C1(_05980_ ), .C2(_05981_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
AOI22_X1 _14048_ ( .A1(_04574_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_05982_ ) );
OAI211_X1 _14049_ ( .A(_05982_ ), .B(_05916_ ), .C1(fanout_net_9 ), .C2(_02149_ ), .ZN(_05983_ ) );
AOI21_X1 _14050_ ( .A(_04125_ ), .B1(_03320_ ), .B2(_03340_ ), .ZN(_05984_ ) );
AND3_X1 _14051_ ( .A1(_05900_ ), .A2(\ID_EX_pc [7] ), .A3(\ID_EX_typ [7] ), .ZN(_05985_ ) );
OAI21_X1 _14052_ ( .A(_05888_ ), .B1(_05984_ ), .B2(_05985_ ), .ZN(_05986_ ) );
NAND2_X1 _14053_ ( .A1(_04341_ ), .A2(\mtvec [7] ), .ZN(_05987_ ) );
NAND4_X1 _14054_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][7] ), .A4(_04571_ ), .ZN(_05988_ ) );
NAND3_X1 _14055_ ( .A1(_04331_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_04332_ ), .ZN(_05989_ ) );
AND4_X1 _14056_ ( .A1(_04584_ ), .A2(_05987_ ), .A3(_05988_ ), .A4(_05989_ ), .ZN(_05990_ ) );
OAI21_X1 _14057_ ( .A(_05990_ ), .B1(_04262_ ), .B2(_04264_ ), .ZN(_05991_ ) );
NAND3_X1 _14058_ ( .A1(_04181_ ), .A2(_04582_ ), .A3(_04183_ ), .ZN(_05992_ ) );
NAND4_X1 _14059_ ( .A1(_05991_ ), .A2(_05909_ ), .A3(_05912_ ), .A4(_05992_ ), .ZN(_05993_ ) );
NAND3_X1 _14060_ ( .A1(_05983_ ), .A2(_05986_ ), .A3(_05993_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
OAI21_X1 _14061_ ( .A(\ID_EX_typ [2] ), .B1(_04603_ ), .B2(_04605_ ), .ZN(_05994_ ) );
AOI21_X1 _14062_ ( .A(fanout_net_9 ), .B1(_02169_ ), .B2(_02170_ ), .ZN(_05995_ ) );
AND2_X1 _14063_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [6] ), .ZN(_05996_ ) );
OAI21_X1 _14064_ ( .A(_05994_ ), .B1(_05995_ ), .B2(_05996_ ), .ZN(_05997_ ) );
OAI211_X1 _14065_ ( .A(_04608_ ), .B(_05894_ ), .C1(_04610_ ), .C2(_04615_ ), .ZN(_05998_ ) );
AOI21_X1 _14066_ ( .A(_05891_ ), .B1(_05997_ ), .B2(_05998_ ), .ZN(_05999_ ) );
AND3_X1 _14067_ ( .A1(_01646_ ), .A2(_04618_ ), .A3(\ID_EX_typ [7] ), .ZN(_06000_ ) );
AOI211_X1 _14068_ ( .A(_05864_ ), .B(_06000_ ), .C1(_03373_ ), .C2(_05898_ ), .ZN(_06001_ ) );
OR2_X1 _14069_ ( .A1(_05999_ ), .A2(_06001_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
NAND3_X1 _14070_ ( .A1(_02093_ ), .A2(_02835_ ), .A3(_02094_ ), .ZN(_06002_ ) );
NAND2_X1 _14071_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [5] ), .ZN(_06003_ ) );
AND2_X1 _14072_ ( .A1(_06002_ ), .A2(_06003_ ), .ZN(_06004_ ) );
AOI21_X1 _14073_ ( .A(_06004_ ), .B1(\ID_EX_typ [2] ), .B2(_04637_ ), .ZN(_06005_ ) );
NOR3_X1 _14074_ ( .A1(_04633_ ), .A2(_05885_ ), .A3(_04635_ ), .ZN(_06006_ ) );
OAI21_X1 _14075_ ( .A(_05916_ ), .B1(_06005_ ), .B2(_06006_ ), .ZN(_06007_ ) );
AND4_X1 _14076_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06008_ ) );
AOI21_X1 _14077_ ( .A(_06008_ ), .B1(_03397_ ), .B2(_05898_ ), .ZN(_06009_ ) );
OAI21_X1 _14078_ ( .A(_06007_ ), .B1(_05871_ ), .B2(_06009_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
AOI221_X4 _14079_ ( .A(_05860_ ), .B1(fanout_net_9 ), .B2(_02119_ ), .C1(_04671_ ), .C2(\ID_EX_typ [2] ), .ZN(_06010_ ) );
OAI21_X1 _14080_ ( .A(_06010_ ), .B1(fanout_net_9 ), .B2(_02118_ ), .ZN(_06011_ ) );
NAND3_X1 _14081_ ( .A1(_04670_ ), .A2(_05909_ ), .A3(_05912_ ), .ZN(_06012_ ) );
MUX2_X1 _14082_ ( .A(_04672_ ), .B(_03420_ ), .S(_02838_ ), .Z(_06013_ ) );
OAI211_X1 _14083_ ( .A(_06011_ ), .B(_06012_ ), .C1(_05865_ ), .C2(_06013_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
OAI22_X1 _14084_ ( .A1(_04699_ ), .A2(_03982_ ), .B1(_04227_ ), .B2(\ID_EX_imm [3] ), .ZN(_06014_ ) );
AOI21_X1 _14085_ ( .A(_06014_ ), .B1(_05009_ ), .B2(_03904_ ), .ZN(_06015_ ) );
NOR3_X1 _14086_ ( .A1(_04696_ ), .A2(_05885_ ), .A3(_04698_ ), .ZN(_06016_ ) );
OAI21_X1 _14087_ ( .A(_05916_ ), .B1(_06015_ ), .B2(_06016_ ), .ZN(_06017_ ) );
AND4_X1 _14088_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06018_ ) );
AOI21_X1 _14089_ ( .A(_06018_ ), .B1(_03691_ ), .B2(_05898_ ), .ZN(_06019_ ) );
OAI21_X1 _14090_ ( .A(_06017_ ), .B1(_05871_ ), .B2(_06019_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
AOI22_X1 _14091_ ( .A1(_04728_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_01969_ ), .ZN(_06020_ ) );
NAND3_X1 _14092_ ( .A1(_01989_ ), .A2(_04227_ ), .A3(_01990_ ), .ZN(_06021_ ) );
AND2_X1 _14093_ ( .A1(_06020_ ), .A2(_06021_ ), .ZN(_06022_ ) );
AOI21_X1 _14094_ ( .A(_05885_ ), .B1(_04726_ ), .B2(_04735_ ), .ZN(_06023_ ) );
OAI21_X1 _14095_ ( .A(_05916_ ), .B1(_06022_ ), .B2(_06023_ ), .ZN(_06024_ ) );
MUX2_X1 _14096_ ( .A(_04992_ ), .B(_03716_ ), .S(_04812_ ), .Z(_06025_ ) );
OAI21_X1 _14097_ ( .A(_06024_ ), .B1(_05871_ ), .B2(_06025_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
OAI22_X1 _14098_ ( .A1(_04144_ ), .A2(_05008_ ), .B1(_04976_ ), .B2(\ID_EX_imm [29] ), .ZN(_06026_ ) );
AOI21_X1 _14099_ ( .A(_06026_ ), .B1(_05009_ ), .B2(_03738_ ), .ZN(_06027_ ) );
NOR3_X1 _14100_ ( .A1(_04132_ ), .A2(_05885_ ), .A3(_04143_ ), .ZN(_06028_ ) );
OAI21_X1 _14101_ ( .A(_05865_ ), .B1(_06027_ ), .B2(_06028_ ), .ZN(_06029_ ) );
BUF_X4 _14102_ ( .A(_05861_ ), .Z(_06030_ ) );
NAND3_X1 _14103_ ( .A1(_05900_ ), .A2(_02825_ ), .A3(\ID_EX_typ [7] ), .ZN(_06031_ ) );
OAI211_X1 _14104_ ( .A(_06030_ ), .B(_06031_ ), .C1(_03594_ ), .C2(_04163_ ), .ZN(_06032_ ) );
NAND2_X1 _14105_ ( .A1(_06029_ ), .A2(_06032_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
AOI21_X1 _14106_ ( .A(fanout_net_9 ), .B1(_02011_ ), .B2(_02013_ ), .ZN(_06033_ ) );
AND2_X1 _14107_ ( .A1(fanout_net_9 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_06034_ ) );
NOR2_X1 _14108_ ( .A1(_06033_ ), .A2(_06034_ ), .ZN(_06035_ ) );
AOI21_X1 _14109_ ( .A(_05885_ ), .B1(_04747_ ), .B2(_04748_ ), .ZN(_06036_ ) );
INV_X1 _14110_ ( .A(_04749_ ), .ZN(_06037_ ) );
OAI221_X1 _14111_ ( .A(_05879_ ), .B1(_06035_ ), .B2(_06036_ ), .C1(_06037_ ), .C2(_05008_ ), .ZN(_06038_ ) );
NAND3_X1 _14112_ ( .A1(_03622_ ), .A2(_03642_ ), .A3(_05898_ ), .ZN(_06039_ ) );
OAI211_X1 _14113_ ( .A(_06039_ ), .B(_06030_ ), .C1(\ID_EX_pc [1] ), .C2(_05898_ ), .ZN(_06040_ ) );
NAND2_X1 _14114_ ( .A1(_06038_ ), .A2(_06040_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
INV_X1 _14115_ ( .A(_04816_ ), .ZN(_06041_ ) );
AOI22_X1 _14116_ ( .A1(_04816_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_03919_ ), .ZN(_06042_ ) );
OR2_X1 _14117_ ( .A1(_03645_ ), .A2(fanout_net_9 ), .ZN(_06043_ ) );
AOI221_X4 _14118_ ( .A(_05860_ ), .B1(_06041_ ), .B2(_05894_ ), .C1(_06042_ ), .C2(_06043_ ), .ZN(_06044_ ) );
MUX2_X1 _14119_ ( .A(_04800_ ), .B(_03669_ ), .S(_04812_ ), .Z(_06045_ ) );
AOI21_X1 _14120_ ( .A(_06044_ ), .B1(_05862_ ), .B2(_06045_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
OAI21_X1 _14121_ ( .A(\ID_EX_typ [2] ), .B1(_04468_ ), .B2(_04470_ ), .ZN(_06046_ ) );
AOI21_X1 _14122_ ( .A(fanout_net_9 ), .B1(_01763_ ), .B2(_01764_ ), .ZN(_06047_ ) );
AND2_X1 _14123_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [28] ), .ZN(_06048_ ) );
OAI21_X1 _14124_ ( .A(_06046_ ), .B1(_06047_ ), .B2(_06048_ ), .ZN(_06049_ ) );
OR3_X1 _14125_ ( .A1(_04468_ ), .A2(_05884_ ), .A3(_04470_ ), .ZN(_06050_ ) );
NAND2_X1 _14126_ ( .A1(_06049_ ), .A2(_06050_ ), .ZN(_06051_ ) );
MUX2_X1 _14127_ ( .A(\ID_EX_pc [28] ), .B(_03616_ ), .S(_02838_ ), .Z(_06052_ ) );
MUX2_X1 _14128_ ( .A(_06051_ ), .B(_06052_ ), .S(_05867_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
AOI22_X1 _14129_ ( .A1(_04777_ ), .A2(\ID_EX_typ [2] ), .B1(_03763_ ), .B2(_04976_ ), .ZN(_06053_ ) );
OAI211_X1 _14130_ ( .A(_06053_ ), .B(_05870_ ), .C1(_05009_ ), .C2(\ID_EX_imm [27] ), .ZN(_06054_ ) );
NAND4_X1 _14131_ ( .A1(_04774_ ), .A2(_05909_ ), .A3(_05894_ ), .A4(_04776_ ), .ZN(_06055_ ) );
AND3_X1 _14132_ ( .A1(_05900_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_06056_ ) );
AOI21_X1 _14133_ ( .A(_06056_ ), .B1(_03501_ ), .B2(_05898_ ), .ZN(_06057_ ) );
OAI211_X1 _14134_ ( .A(_06054_ ), .B(_06055_ ), .C1(_05865_ ), .C2(_06057_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
INV_X1 _14135_ ( .A(_04824_ ), .ZN(_06058_ ) );
OAI22_X1 _14136_ ( .A1(_04824_ ), .A2(_05885_ ), .B1(_04976_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06059_ ) );
AOI21_X1 _14137_ ( .A(fanout_net_9 ), .B1(_02508_ ), .B2(_02509_ ), .ZN(_06060_ ) );
OAI221_X1 _14138_ ( .A(_05909_ ), .B1(_05008_ ), .B2(_06058_ ), .C1(_06059_ ), .C2(_06060_ ), .ZN(_06061_ ) );
AND3_X1 _14139_ ( .A1(_05900_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_06062_ ) );
AOI21_X1 _14140_ ( .A(_06062_ ), .B1(_03525_ ), .B2(_05898_ ), .ZN(_06063_ ) );
OAI21_X1 _14141_ ( .A(_06061_ ), .B1(_05871_ ), .B2(_06063_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
AOI22_X1 _14142_ ( .A1(_04976_ ), .A2(_03476_ ), .B1(_04848_ ), .B2(\ID_EX_typ [2] ), .ZN(_06064_ ) );
OAI211_X1 _14143_ ( .A(_06064_ ), .B(_05870_ ), .C1(_05009_ ), .C2(\ID_EX_imm [25] ), .ZN(_06065_ ) );
OR3_X1 _14144_ ( .A1(_04262_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_04264_ ), .ZN(_06066_ ) );
NAND2_X1 _14145_ ( .A1(_04341_ ), .A2(\mtvec [25] ), .ZN(_06067_ ) );
NAND4_X1 _14146_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][25] ), .A4(_04571_ ), .ZN(_06068_ ) );
NAND3_X1 _14147_ ( .A1(_04331_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_04332_ ), .ZN(_06069_ ) );
AND4_X1 _14148_ ( .A1(_04862_ ), .A2(_06067_ ), .A3(_06068_ ), .A4(_06069_ ), .ZN(_06070_ ) );
OAI21_X1 _14149_ ( .A(_06070_ ), .B1(_04262_ ), .B2(_04264_ ), .ZN(_06071_ ) );
NAND4_X1 _14150_ ( .A1(_06066_ ), .A2(_05909_ ), .A3(_05894_ ), .A4(_06071_ ), .ZN(_06072_ ) );
AND3_X1 _14151_ ( .A1(_05900_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06073_ ) );
AOI21_X1 _14152_ ( .A(_06073_ ), .B1(_03475_ ), .B2(_05898_ ), .ZN(_06074_ ) );
OAI211_X1 _14153_ ( .A(_06065_ ), .B(_06072_ ), .C1(_05865_ ), .C2(_06074_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
AOI22_X1 _14154_ ( .A1(_04881_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02433_ ), .ZN(_06075_ ) );
OAI211_X1 _14155_ ( .A(_06075_ ), .B(_05870_ ), .C1(\ID_EX_typ [0] ), .C2(_02432_ ), .ZN(_06076_ ) );
AND3_X1 _14156_ ( .A1(_04878_ ), .A2(_02576_ ), .A3(_04879_ ), .ZN(_06077_ ) );
NAND2_X1 _14157_ ( .A1(_06077_ ), .A2(_05912_ ), .ZN(_06078_ ) );
AND3_X1 _14158_ ( .A1(_01646_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_typ [7] ), .ZN(_06079_ ) );
AOI21_X1 _14159_ ( .A(_06079_ ), .B1(_03450_ ), .B2(_05898_ ), .ZN(_06080_ ) );
OAI211_X1 _14160_ ( .A(_06076_ ), .B(_06078_ ), .C1(_05865_ ), .C2(_06080_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
AOI22_X1 _14161_ ( .A1(_04976_ ), .A2(_03058_ ), .B1(_04905_ ), .B2(\ID_EX_typ [2] ), .ZN(_06081_ ) );
OAI211_X1 _14162_ ( .A(_06081_ ), .B(_05870_ ), .C1(_05009_ ), .C2(\ID_EX_imm [23] ), .ZN(_06082_ ) );
OR3_X1 _14163_ ( .A1(_04262_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_04264_ ), .ZN(_06083_ ) );
NAND3_X1 _14164_ ( .A1(_04388_ ), .A2(\mepc [23] ), .A3(_04571_ ), .ZN(_06084_ ) );
NAND2_X1 _14165_ ( .A1(_04341_ ), .A2(\mtvec [23] ), .ZN(_06085_ ) );
NAND4_X1 _14166_ ( .A1(_02698_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][23] ), .A4(_04571_ ), .ZN(_06086_ ) );
NAND3_X1 _14167_ ( .A1(_04331_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_04332_ ), .ZN(_06087_ ) );
AND4_X1 _14168_ ( .A1(_06084_ ), .A2(_06085_ ), .A3(_06086_ ), .A4(_06087_ ), .ZN(_06088_ ) );
OAI21_X1 _14169_ ( .A(_06088_ ), .B1(_04262_ ), .B2(_04264_ ), .ZN(_06089_ ) );
NAND4_X1 _14170_ ( .A1(_06083_ ), .A2(_05909_ ), .A3(_05894_ ), .A4(_06089_ ), .ZN(_06090_ ) );
AOI21_X1 _14171_ ( .A(_04125_ ), .B1(_03036_ ), .B2(_03056_ ), .ZN(_06091_ ) );
AOI21_X1 _14172_ ( .A(_06091_ ), .B1(\ID_EX_pc [23] ), .B2(_04163_ ), .ZN(_06092_ ) );
OAI211_X1 _14173_ ( .A(_06082_ ), .B(_06090_ ), .C1(_05865_ ), .C2(_06092_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _14174_ ( .A1(_01794_ ), .A2(\ID_EX_typ [0] ), .ZN(_06093_ ) );
OAI221_X1 _14175_ ( .A(_06093_ ), .B1(\ID_EX_typ [0] ), .B2(_01793_ ), .C1(_04919_ ), .C2(_05008_ ), .ZN(_06094_ ) );
NAND3_X1 _14176_ ( .A1(_04917_ ), .A2(_05894_ ), .A3(_04918_ ), .ZN(_06095_ ) );
NAND3_X1 _14177_ ( .A1(_06094_ ), .A2(_05909_ ), .A3(_06095_ ), .ZN(_06096_ ) );
NAND4_X1 _14178_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06097_ ) );
OAI211_X1 _14179_ ( .A(_05867_ ), .B(_06097_ ), .C1(_03032_ ), .C2(_04125_ ), .ZN(_06098_ ) );
AND2_X1 _14180_ ( .A1(_06096_ ), .A2(_06098_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
NAND4_X1 _14181_ ( .A1(_02678_ ), .A2(_04204_ ), .A3(\mtvec [31] ), .A4(_02688_ ), .ZN(_06099_ ) );
NAND4_X1 _14182_ ( .A1(_02691_ ), .A2(_04231_ ), .A3(\mepc [31] ), .A4(_04205_ ), .ZN(_06100_ ) );
NAND4_X1 _14183_ ( .A1(_04204_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04205_ ), .A4(_04117_ ), .ZN(_06101_ ) );
NAND4_X1 _14184_ ( .A1(_04231_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[3][31] ), .A4(_04205_ ), .ZN(_06102_ ) );
AND4_X1 _14185_ ( .A1(_06099_ ), .A2(_06100_ ), .A3(_06101_ ), .A4(_06102_ ), .ZN(_06103_ ) );
OR2_X1 _14186_ ( .A1(_02664_ ), .A2(_06103_ ), .ZN(_06104_ ) );
NAND3_X1 _14187_ ( .A1(_02715_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_02717_ ), .ZN(_06105_ ) );
AND2_X1 _14188_ ( .A1(_06104_ ), .A2(_06105_ ), .ZN(_06106_ ) );
INV_X1 _14189_ ( .A(_06106_ ), .ZN(_06107_ ) );
OAI22_X1 _14190_ ( .A1(_06106_ ), .A2(_05885_ ), .B1(_04976_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_06108_ ) );
AND3_X1 _14191_ ( .A1(_02569_ ), .A2(_04976_ ), .A3(_02570_ ), .ZN(_06109_ ) );
OAI221_X1 _14192_ ( .A(_05879_ ), .B1(_05008_ ), .B2(_06107_ ), .C1(_06108_ ), .C2(_06109_ ), .ZN(_06110_ ) );
NAND4_X1 _14193_ ( .A1(_04990_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06111_ ) );
OAI211_X1 _14194_ ( .A(_06030_ ), .B(_06111_ ), .C1(_03571_ ), .C2(_04163_ ), .ZN(_06112_ ) );
NAND2_X1 _14195_ ( .A1(_06110_ ), .A2(_06112_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
OR3_X1 _14196_ ( .A1(_04939_ ), .A2(_05861_ ), .A3(_04941_ ), .ZN(_06113_ ) );
NOR3_X1 _14197_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_06114_ ) );
AND2_X1 _14198_ ( .A1(\ID_EX_typ [3] ), .A2(\ID_EX_typ [2] ), .ZN(_06115_ ) );
AND2_X2 _14199_ ( .A1(_06114_ ), .A2(_06115_ ), .ZN(_06116_ ) );
INV_X1 _14200_ ( .A(_06116_ ), .ZN(_06117_ ) );
BUF_X4 _14201_ ( .A(_06117_ ), .Z(_06118_ ) );
NOR2_X1 _14202_ ( .A1(_04951_ ), .A2(_06118_ ), .ZN(_06119_ ) );
AND2_X1 _14203_ ( .A1(_03083_ ), .A2(_01869_ ), .ZN(_06120_ ) );
OAI21_X1 _14204_ ( .A(_04056_ ), .B1(_04025_ ), .B2(_03008_ ), .ZN(_06121_ ) );
AOI21_X1 _14205_ ( .A(_06120_ ), .B1(_06121_ ), .B2(_03085_ ), .ZN(_06122_ ) );
XNOR2_X1 _14206_ ( .A(_06122_ ), .B(_03109_ ), .ZN(_06123_ ) );
AND3_X1 _14207_ ( .A1(_02859_ ), .A2(\ID_EX_typ [3] ), .A3(_03982_ ), .ZN(_06124_ ) );
AND2_X2 _14208_ ( .A1(_06124_ ), .A2(_03728_ ), .ZN(_06125_ ) );
AND2_X1 _14209_ ( .A1(_06123_ ), .A2(_06125_ ), .ZN(_06126_ ) );
NOR3_X2 _14210_ ( .A1(_04073_ ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_06127_ ) );
BUF_X2 _14211_ ( .A(_06115_ ), .Z(_06128_ ) );
AND3_X1 _14212_ ( .A1(_06127_ ), .A2(\ID_EX_imm [21] ), .A3(_06128_ ), .ZN(_06129_ ) );
NOR3_X1 _14213_ ( .A1(_06119_ ), .A2(_06126_ ), .A3(_06129_ ), .ZN(_06130_ ) );
AND2_X1 _14214_ ( .A1(_01648_ ), .A2(_01656_ ), .ZN(_06131_ ) );
INV_X1 _14215_ ( .A(_06131_ ), .ZN(_06132_ ) );
BUF_X4 _14216_ ( .A(_06132_ ), .Z(_06133_ ) );
OAI21_X1 _14217_ ( .A(_04161_ ), .B1(_06130_ ), .B2(_06133_ ), .ZN(_06134_ ) );
BUF_X4 _14218_ ( .A(_04076_ ), .Z(_06135_ ) );
AOI21_X1 _14219_ ( .A(_06135_ ), .B1(_03797_ ), .B2(_02403_ ), .ZN(_06136_ ) );
INV_X1 _14220_ ( .A(_01732_ ), .ZN(_06137_ ) );
BUF_X2 _14221_ ( .A(_03918_ ), .Z(_06138_ ) );
BUF_X2 _14222_ ( .A(_06138_ ), .Z(_06139_ ) );
BUF_X2 _14223_ ( .A(_06139_ ), .Z(_06140_ ) );
BUF_X2 _14224_ ( .A(_03920_ ), .Z(_06141_ ) );
BUF_X2 _14225_ ( .A(_06141_ ), .Z(_06142_ ) );
BUF_X2 _14226_ ( .A(_06142_ ), .Z(_06143_ ) );
NAND3_X1 _14227_ ( .A1(_06137_ ), .A2(_06140_ ), .A3(_06143_ ), .ZN(_06144_ ) );
BUF_X4 _14228_ ( .A(_03927_ ), .Z(_06145_ ) );
BUF_X4 _14229_ ( .A(_06145_ ), .Z(_06146_ ) );
BUF_X4 _14230_ ( .A(_03921_ ), .Z(_06147_ ) );
NAND2_X1 _14231_ ( .A1(_06147_ ), .A2(_02539_ ), .ZN(_06148_ ) );
NAND3_X1 _14232_ ( .A1(_06144_ ), .A2(_06146_ ), .A3(_06148_ ), .ZN(_06149_ ) );
BUF_X4 _14233_ ( .A(_06145_ ), .Z(_06150_ ) );
BUF_X4 _14234_ ( .A(_06150_ ), .Z(_06151_ ) );
AND2_X1 _14235_ ( .A1(_06147_ ), .A2(_02571_ ), .ZN(_06152_ ) );
OAI21_X1 _14236_ ( .A(_06149_ ), .B1(_06151_ ), .B2(_06152_ ), .ZN(_06153_ ) );
BUF_X4 _14237_ ( .A(_03909_ ), .Z(_06154_ ) );
NOR2_X1 _14238_ ( .A1(_06153_ ), .A2(_06154_ ), .ZN(_06155_ ) );
AND3_X1 _14239_ ( .A1(_06140_ ), .A2(_02514_ ), .A3(_06143_ ), .ZN(_06156_ ) );
INV_X2 _14240_ ( .A(_06145_ ), .ZN(_06157_ ) );
BUF_X4 _14241_ ( .A(_06157_ ), .Z(_06158_ ) );
AOI21_X1 _14242_ ( .A(_02456_ ), .B1(_06140_ ), .B2(_06143_ ), .ZN(_06159_ ) );
NOR3_X1 _14243_ ( .A1(_06156_ ), .A2(_06158_ ), .A3(_06159_ ), .ZN(_06160_ ) );
AND3_X1 _14244_ ( .A1(_06139_ ), .A2(_03732_ ), .A3(_06142_ ), .ZN(_06161_ ) );
AOI21_X1 _14245_ ( .A(_03502_ ), .B1(_06139_ ), .B2(_06142_ ), .ZN(_06162_ ) );
NOR3_X1 _14246_ ( .A1(_06161_ ), .A2(_06162_ ), .A3(_06146_ ), .ZN(_06163_ ) );
OAI21_X1 _14247_ ( .A(_03909_ ), .B1(_06160_ ), .B2(_06163_ ), .ZN(_06164_ ) );
AND3_X1 _14248_ ( .A1(_06140_ ), .A2(_03033_ ), .A3(_06143_ ), .ZN(_06165_ ) );
AOI21_X1 _14249_ ( .A(_01843_ ), .B1(_06140_ ), .B2(_06143_ ), .ZN(_06166_ ) );
OAI21_X1 _14250_ ( .A(_06146_ ), .B1(_06165_ ), .B2(_06166_ ), .ZN(_06167_ ) );
INV_X1 _14251_ ( .A(_02432_ ), .ZN(_06168_ ) );
AND3_X1 _14252_ ( .A1(_06140_ ), .A2(_06168_ ), .A3(_06143_ ), .ZN(_06169_ ) );
AOI21_X1 _14253_ ( .A(_01816_ ), .B1(_06140_ ), .B2(_06143_ ), .ZN(_06170_ ) );
OAI21_X1 _14254_ ( .A(_06158_ ), .B1(_06169_ ), .B2(_06170_ ), .ZN(_06171_ ) );
BUF_X4 _14255_ ( .A(_03908_ ), .Z(_06172_ ) );
NAND3_X1 _14256_ ( .A1(_06167_ ), .A2(_06171_ ), .A3(_06172_ ), .ZN(_06173_ ) );
NAND2_X1 _14257_ ( .A1(_06164_ ), .A2(_06173_ ), .ZN(_06174_ ) );
BUF_X4 _14258_ ( .A(_03912_ ), .Z(_06175_ ) );
MUX2_X1 _14259_ ( .A(_06155_ ), .B(_06174_ ), .S(_06175_ ), .Z(_06176_ ) );
BUF_X2 _14260_ ( .A(_03886_ ), .Z(_06177_ ) );
BUF_X2 _14261_ ( .A(_06177_ ), .Z(_06178_ ) );
AND2_X1 _14262_ ( .A1(_06176_ ), .A2(_06178_ ), .ZN(_06179_ ) );
AND2_X2 _14263_ ( .A1(_04074_ ), .A2(\ID_EX_typ [2] ), .ZN(_06180_ ) );
BUF_X2 _14264_ ( .A(_06180_ ), .Z(_06181_ ) );
OR2_X1 _14265_ ( .A1(_03793_ ), .A2(_03084_ ), .ZN(_06182_ ) );
AND2_X1 _14266_ ( .A1(_03807_ ), .A2(_03958_ ), .ZN(_06183_ ) );
AND3_X1 _14267_ ( .A1(_06183_ ), .A2(_03814_ ), .A3(_03819_ ), .ZN(_06184_ ) );
INV_X1 _14268_ ( .A(_06184_ ), .ZN(_06185_ ) );
OR2_X1 _14269_ ( .A1(_03881_ ), .A2(_03344_ ), .ZN(_06186_ ) );
NOR3_X1 _14270_ ( .A1(_03875_ ), .A2(_03876_ ), .A3(_06186_ ), .ZN(_06187_ ) );
NOR3_X1 _14271_ ( .A1(_03875_ ), .A2(_03876_ ), .A3(_03883_ ), .ZN(_06188_ ) );
NOR2_X1 _14272_ ( .A1(_03886_ ), .A2(_02123_ ), .ZN(_06189_ ) );
NAND2_X1 _14273_ ( .A1(_03896_ ), .A2(_06189_ ), .ZN(_06190_ ) );
INV_X1 _14274_ ( .A(_03889_ ), .ZN(_06191_ ) );
OAI21_X1 _14275_ ( .A(_06190_ ), .B1(_03891_ ), .B2(_06191_ ), .ZN(_06192_ ) );
AOI211_X1 _14276_ ( .A(_03875_ ), .B(_06187_ ), .C1(_06188_ ), .C2(_06192_ ), .ZN(_06193_ ) );
AND4_X1 _14277_ ( .A1(_03877_ ), .A2(_03882_ ), .A3(_03896_ ), .A4(_03898_ ), .ZN(_06194_ ) );
INV_X1 _14278_ ( .A(_03917_ ), .ZN(_06195_ ) );
NOR2_X1 _14279_ ( .A1(_03908_ ), .A2(_03717_ ), .ZN(_06196_ ) );
INV_X1 _14280_ ( .A(_06196_ ), .ZN(_06197_ ) );
NOR2_X1 _14281_ ( .A1(_03921_ ), .A2(_03646_ ), .ZN(_06198_ ) );
AND3_X2 _14282_ ( .A1(_03926_ ), .A2(_03928_ ), .A3(_06198_ ), .ZN(_06199_ ) );
NOR2_X4 _14283_ ( .A1(_06199_ ), .A2(_03925_ ), .ZN(_06200_ ) );
OAI221_X1 _14284_ ( .A(_06197_ ), .B1(_03904_ ), .B2(_06175_ ), .C1(_06200_ ), .C2(_03915_ ), .ZN(_06201_ ) );
NAND3_X1 _14285_ ( .A1(_06194_ ), .A2(_06195_ ), .A3(_06201_ ), .ZN(_06202_ ) );
AND2_X4 _14286_ ( .A1(_06193_ ), .A2(_06202_ ), .ZN(_06203_ ) );
NOR3_X4 _14287_ ( .A1(_06203_ ), .A2(_03865_ ), .A3(_03870_ ), .ZN(_06204_ ) );
AND2_X1 _14288_ ( .A1(_03850_ ), .A2(_03844_ ), .ZN(_06205_ ) );
AND3_X1 _14289_ ( .A1(_06205_ ), .A2(_03834_ ), .A3(_03839_ ), .ZN(_06206_ ) );
AND2_X2 _14290_ ( .A1(_03859_ ), .A2(_03855_ ), .ZN(_06207_ ) );
NAND3_X1 _14291_ ( .A1(_06204_ ), .A2(_06206_ ), .A3(_06207_ ), .ZN(_06208_ ) );
NOR2_X1 _14292_ ( .A1(_03868_ ), .A2(_03317_ ), .ZN(_06209_ ) );
INV_X1 _14293_ ( .A(_03938_ ), .ZN(_06210_ ) );
AOI21_X1 _14294_ ( .A(_03939_ ), .B1(_06209_ ), .B2(_06210_ ), .ZN(_06211_ ) );
INV_X1 _14295_ ( .A(_06211_ ), .ZN(_06212_ ) );
AND2_X1 _14296_ ( .A1(_06212_ ), .A2(_06207_ ), .ZN(_06213_ ) );
NOR2_X1 _14297_ ( .A1(_03858_ ), .A2(_03241_ ), .ZN(_06214_ ) );
NOR2_X1 _14298_ ( .A1(_03854_ ), .A2(_03266_ ), .ZN(_06215_ ) );
AND2_X1 _14299_ ( .A1(_03859_ ), .A2(_06215_ ), .ZN(_06216_ ) );
NOR3_X4 _14300_ ( .A1(_06213_ ), .A2(_06214_ ), .A3(_06216_ ), .ZN(_06217_ ) );
INV_X1 _14301_ ( .A(_06206_ ), .ZN(_06218_ ) );
NOR2_X1 _14302_ ( .A1(_06217_ ), .A2(_06218_ ), .ZN(_06219_ ) );
NOR2_X1 _14303_ ( .A1(_03833_ ), .A2(_03954_ ), .ZN(_06220_ ) );
NOR2_X1 _14304_ ( .A1(_03849_ ), .A2(_03214_ ), .ZN(_06221_ ) );
NOR2_X1 _14305_ ( .A1(_03843_ ), .A2(_03188_ ), .ZN(_06222_ ) );
AOI21_X1 _14306_ ( .A(_06221_ ), .B1(_03850_ ), .B2(_06222_ ), .ZN(_06223_ ) );
NOR3_X1 _14307_ ( .A1(_06223_ ), .A2(_03835_ ), .A3(_03840_ ), .ZN(_06224_ ) );
NOR2_X1 _14308_ ( .A1(_03838_ ), .A2(_03135_ ), .ZN(_06225_ ) );
AND2_X1 _14309_ ( .A1(_03834_ ), .A2(_06225_ ), .ZN(_06226_ ) );
NOR4_X4 _14310_ ( .A1(_06219_ ), .A2(_06220_ ), .A3(_06224_ ), .A4(_06226_ ), .ZN(_06227_ ) );
AOI21_X1 _14311_ ( .A(_06185_ ), .B1(_06208_ ), .B2(_06227_ ), .ZN(_06228_ ) );
INV_X1 _14312_ ( .A(_06228_ ), .ZN(_06229_ ) );
NOR2_X1 _14313_ ( .A1(_03810_ ), .A2(_02953_ ), .ZN(_06230_ ) );
AND2_X1 _14314_ ( .A1(_03807_ ), .A2(_06230_ ), .ZN(_06231_ ) );
NOR2_X1 _14315_ ( .A1(_03806_ ), .A2(_02922_ ), .ZN(_06232_ ) );
OAI211_X1 _14316_ ( .A(_03814_ ), .B(_03819_ ), .C1(_06231_ ), .C2(_06232_ ), .ZN(_06233_ ) );
OR2_X1 _14317_ ( .A1(_03802_ ), .A2(_02977_ ), .ZN(_06234_ ) );
NOR2_X1 _14318_ ( .A1(_03818_ ), .A2(_03005_ ), .ZN(_06235_ ) );
NAND2_X1 _14319_ ( .A1(_03814_ ), .A2(_06235_ ), .ZN(_06236_ ) );
AND3_X1 _14320_ ( .A1(_06233_ ), .A2(_06234_ ), .A3(_06236_ ), .ZN(_06237_ ) );
AND2_X1 _14321_ ( .A1(_06229_ ), .A2(_06237_ ), .ZN(_06238_ ) );
INV_X1 _14322_ ( .A(_03794_ ), .ZN(_06239_ ) );
OAI21_X1 _14323_ ( .A(_06182_ ), .B1(_06238_ ), .B2(_06239_ ), .ZN(_06240_ ) );
INV_X1 _14324_ ( .A(_03798_ ), .ZN(_06241_ ) );
XNOR2_X1 _14325_ ( .A(_06240_ ), .B(_06241_ ), .ZN(_06242_ ) );
NOR2_X1 _14326_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06243_ ) );
INV_X1 _14327_ ( .A(_06243_ ), .ZN(_06244_ ) );
NOR2_X1 _14328_ ( .A1(_03723_ ), .A2(_06244_ ), .ZN(_06245_ ) );
AOI221_X4 _14329_ ( .A(_06136_ ), .B1(_06179_ ), .B2(_06181_ ), .C1(_06242_ ), .C2(_06245_ ), .ZN(_06246_ ) );
AND2_X2 _14330_ ( .A1(_03985_ ), .A2(\ID_EX_typ [2] ), .ZN(_06247_ ) );
BUF_X4 _14331_ ( .A(_06247_ ), .Z(_06248_ ) );
BUF_X4 _14332_ ( .A(_06248_ ), .Z(_06249_ ) );
AND2_X1 _14333_ ( .A1(_06145_ ), .A2(_03921_ ), .ZN(_06250_ ) );
AND2_X4 _14334_ ( .A1(_06250_ ), .A2(_03908_ ), .ZN(_06251_ ) );
AND2_X1 _14335_ ( .A1(_06251_ ), .A2(_03912_ ), .ZN(_06252_ ) );
AND2_X4 _14336_ ( .A1(_06252_ ), .A2(_03886_ ), .ZN(_06253_ ) );
NOR2_X1 _14337_ ( .A1(_06253_ ), .A2(_06191_ ), .ZN(_06254_ ) );
INV_X1 _14338_ ( .A(_06254_ ), .ZN(_06255_ ) );
AND3_X1 _14339_ ( .A1(_03872_ ), .A2(_03873_ ), .A3(_03881_ ), .ZN(_06256_ ) );
AND2_X1 _14340_ ( .A1(_06255_ ), .A2(_06256_ ), .ZN(_06257_ ) );
NOR4_X1 _14341_ ( .A1(_06253_ ), .A2(_03874_ ), .A3(_03881_ ), .A4(_06191_ ), .ZN(_06258_ ) );
OAI21_X1 _14342_ ( .A(_02571_ ), .B1(_06257_ ), .B2(_06258_ ), .ZN(_06259_ ) );
OR3_X1 _14343_ ( .A1(_06257_ ), .A2(_03863_ ), .A3(_03868_ ), .ZN(_06260_ ) );
NAND3_X1 _14344_ ( .A1(_06255_ ), .A2(_03868_ ), .A3(_06256_ ), .ZN(_06261_ ) );
NOR2_X2 _14345_ ( .A1(_06261_ ), .A2(_03941_ ), .ZN(_06262_ ) );
INV_X1 _14346_ ( .A(_06262_ ), .ZN(_06263_ ) );
AOI21_X1 _14347_ ( .A(_06259_ ), .B1(_06260_ ), .B2(_06263_ ), .ZN(_06264_ ) );
AND2_X1 _14348_ ( .A1(_03858_ ), .A2(_03854_ ), .ZN(_06265_ ) );
AND2_X1 _14349_ ( .A1(_06262_ ), .A2(_06265_ ), .ZN(_06266_ ) );
NOR3_X1 _14350_ ( .A1(_06262_ ), .A2(_03858_ ), .A3(_03854_ ), .ZN(_06267_ ) );
OAI21_X1 _14351_ ( .A(_06264_ ), .B1(_06266_ ), .B2(_06267_ ), .ZN(_06268_ ) );
AND3_X1 _14352_ ( .A1(_03838_ ), .A2(_03849_ ), .A3(_03843_ ), .ZN(_06269_ ) );
AND4_X1 _14353_ ( .A1(_03787_ ), .A2(_03793_ ), .A3(_03782_ ), .A4(_03810_ ), .ZN(_06270_ ) );
NAND2_X1 _14354_ ( .A1(_03746_ ), .A2(_03748_ ), .ZN(_06271_ ) );
NOR4_X1 _14355_ ( .A1(_03731_ ), .A2(_03737_ ), .A3(_06271_ ), .A4(_03978_ ), .ZN(_06272_ ) );
AND4_X1 _14356_ ( .A1(_03797_ ), .A2(_03806_ ), .A3(_03802_ ), .A4(_03818_ ), .ZN(_06273_ ) );
AND2_X1 _14357_ ( .A1(_03771_ ), .A2(_03775_ ), .ZN(_06274_ ) );
AND3_X1 _14358_ ( .A1(_06274_ ), .A2(_03762_ ), .A3(_03755_ ), .ZN(_06275_ ) );
NAND4_X1 _14359_ ( .A1(_06270_ ), .A2(_06272_ ), .A3(_06273_ ), .A4(_06275_ ), .ZN(_06276_ ) );
AND4_X1 _14360_ ( .A1(_03833_ ), .A2(_06266_ ), .A3(_06269_ ), .A4(_06276_ ), .ZN(_06277_ ) );
NOR2_X2 _14361_ ( .A1(_06268_ ), .A2(_06277_ ), .ZN(_06278_ ) );
NAND4_X1 _14362_ ( .A1(_06262_ ), .A2(_03833_ ), .A3(_06265_ ), .A4(_06269_ ), .ZN(_06279_ ) );
NOR4_X1 _14363_ ( .A1(_03787_ ), .A2(_03793_ ), .A3(_03782_ ), .A4(_03810_ ), .ZN(_06280_ ) );
NOR4_X1 _14364_ ( .A1(_03833_ ), .A2(_03838_ ), .A3(_03849_ ), .A4(_03843_ ), .ZN(_06281_ ) );
NOR4_X1 _14365_ ( .A1(_03806_ ), .A2(_03802_ ), .A3(_03818_ ), .A4(_03797_ ), .ZN(_06282_ ) );
NAND3_X1 _14366_ ( .A1(_06280_ ), .A2(_06281_ ), .A3(_06282_ ), .ZN(_06283_ ) );
OR4_X1 _14367_ ( .A1(_03762_ ), .A2(_03755_ ), .A3(_03771_ ), .A4(_03775_ ), .ZN(_06284_ ) );
NAND4_X1 _14368_ ( .A1(_03731_ ), .A2(_03737_ ), .A3(_06271_ ), .A4(_03978_ ), .ZN(_06285_ ) );
OR3_X1 _14369_ ( .A1(_06283_ ), .A2(_06284_ ), .A3(_06285_ ), .ZN(_06286_ ) );
OAI21_X1 _14370_ ( .A(_06279_ ), .B1(_06266_ ), .B2(_06286_ ), .ZN(_06287_ ) );
AND2_X2 _14371_ ( .A1(_06278_ ), .A2(_06287_ ), .ZN(_06288_ ) );
XNOR2_X1 _14372_ ( .A(_06253_ ), .B(_03889_ ), .ZN(_06289_ ) );
AND2_X4 _14373_ ( .A1(_06288_ ), .A2(_06289_ ), .ZN(_06290_ ) );
INV_X1 _14374_ ( .A(_06290_ ), .ZN(_06291_ ) );
XNOR2_X1 _14375_ ( .A(_06252_ ), .B(_03886_ ), .ZN(_06292_ ) );
NOR2_X1 _14376_ ( .A1(_06292_ ), .A2(_03889_ ), .ZN(_06293_ ) );
INV_X1 _14377_ ( .A(_06293_ ), .ZN(_06294_ ) );
INV_X1 _14378_ ( .A(_06292_ ), .ZN(_06295_ ) );
XNOR2_X1 _14379_ ( .A(_06151_ ), .B(_06147_ ), .ZN(_06296_ ) );
BUF_X4 _14380_ ( .A(_06154_ ), .Z(_06297_ ) );
OR2_X1 _14381_ ( .A1(_06296_ ), .A2(_06297_ ), .ZN(_06298_ ) );
XNOR2_X1 _14382_ ( .A(_06251_ ), .B(_03911_ ), .ZN(_06299_ ) );
INV_X1 _14383_ ( .A(_06299_ ), .ZN(_06300_ ) );
BUF_X2 _14384_ ( .A(_06300_ ), .Z(_06301_ ) );
NAND4_X1 _14385_ ( .A1(_06278_ ), .A2(_06298_ ), .A3(_06301_ ), .A4(_06287_ ), .ZN(_06302_ ) );
AOI22_X1 _14386_ ( .A1(_06291_ ), .A2(_06294_ ), .B1(_06295_ ), .B2(_06302_ ), .ZN(_06303_ ) );
OAI21_X1 _14387_ ( .A(_06249_ ), .B1(_06303_ ), .B2(_06179_ ), .ZN(_06304_ ) );
INV_X1 _14388_ ( .A(_04070_ ), .ZN(_06305_ ) );
BUF_X2 _14389_ ( .A(_06139_ ), .Z(_06306_ ) );
BUF_X2 _14390_ ( .A(_06142_ ), .Z(_06307_ ) );
AND3_X1 _14391_ ( .A1(_06306_ ), .A2(_02123_ ), .A3(_06307_ ), .ZN(_06308_ ) );
BUF_X4 _14392_ ( .A(_06158_ ), .Z(_06309_ ) );
AOI21_X1 _14393_ ( .A(_02096_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_06310_ ) );
NOR3_X1 _14394_ ( .A1(_06308_ ), .A2(_06309_ ), .A3(_06310_ ), .ZN(_06311_ ) );
AND3_X1 _14395_ ( .A1(_06140_ ), .A2(_03717_ ), .A3(_06143_ ), .ZN(_06312_ ) );
AOI21_X1 _14396_ ( .A(_02069_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_06313_ ) );
NOR3_X1 _14397_ ( .A1(_06312_ ), .A2(_06313_ ), .A3(_06146_ ), .ZN(_06314_ ) );
OR3_X1 _14398_ ( .A1(_06311_ ), .A2(_06314_ ), .A3(_06154_ ), .ZN(_06315_ ) );
BUF_X4 _14399_ ( .A(_06172_ ), .Z(_06316_ ) );
BUF_X4 _14400_ ( .A(_06316_ ), .Z(_06317_ ) );
BUF_X2 _14401_ ( .A(_06158_ ), .Z(_06318_ ) );
AOI21_X1 _14402_ ( .A(_02014_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_06319_ ) );
NOR3_X1 _14403_ ( .A1(_03922_ ), .A2(_06318_ ), .A3(_06319_ ), .ZN(_06320_ ) );
OAI21_X1 _14404_ ( .A(_06315_ ), .B1(_06317_ ), .B2(_06320_ ), .ZN(_06321_ ) );
BUF_X2 _14405_ ( .A(_06177_ ), .Z(_06322_ ) );
BUF_X4 _14406_ ( .A(_03911_ ), .Z(_06323_ ) );
OR3_X1 _14407_ ( .A1(_06321_ ), .A2(_06322_ ), .A3(_06323_ ), .ZN(_06324_ ) );
BUF_X4 _14408_ ( .A(_06154_ ), .Z(_06325_ ) );
BUF_X2 _14409_ ( .A(_06139_ ), .Z(_06326_ ) );
BUF_X2 _14410_ ( .A(_06142_ ), .Z(_06327_ ) );
AND3_X1 _14411_ ( .A1(_06326_ ), .A2(_03317_ ), .A3(_06327_ ), .ZN(_06328_ ) );
BUF_X4 _14412_ ( .A(_06309_ ), .Z(_06329_ ) );
AOI21_X1 _14413_ ( .A(_02225_ ), .B1(_06326_ ), .B2(_06327_ ), .ZN(_06330_ ) );
NOR3_X1 _14414_ ( .A1(_06328_ ), .A2(_06329_ ), .A3(_06330_ ), .ZN(_06331_ ) );
AND3_X1 _14415_ ( .A1(_06306_ ), .A2(_03344_ ), .A3(_06307_ ), .ZN(_06332_ ) );
AOI21_X1 _14416_ ( .A(_02149_ ), .B1(_06326_ ), .B2(_06327_ ), .ZN(_06333_ ) );
BUF_X4 _14417_ ( .A(_06151_ ), .Z(_06334_ ) );
NOR3_X1 _14418_ ( .A1(_06332_ ), .A2(_06333_ ), .A3(_06334_ ), .ZN(_06335_ ) );
OAI21_X1 _14419_ ( .A(_06325_ ), .B1(_06331_ ), .B2(_06335_ ), .ZN(_06336_ ) );
AND3_X1 _14420_ ( .A1(_06306_ ), .A2(_03188_ ), .A3(_06307_ ), .ZN(_06337_ ) );
AOI21_X1 _14421_ ( .A(_03213_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_06338_ ) );
NOR3_X1 _14422_ ( .A1(_06337_ ), .A2(_06329_ ), .A3(_06338_ ), .ZN(_06339_ ) );
AND3_X1 _14423_ ( .A1(_06326_ ), .A2(_03266_ ), .A3(_06327_ ), .ZN(_06340_ ) );
AOI21_X1 _14424_ ( .A(_02272_ ), .B1(_06326_ ), .B2(_06327_ ), .ZN(_06341_ ) );
BUF_X4 _14425_ ( .A(_06146_ ), .Z(_06342_ ) );
NOR3_X1 _14426_ ( .A1(_06340_ ), .A2(_06341_ ), .A3(_06342_ ), .ZN(_06343_ ) );
OAI21_X1 _14427_ ( .A(_06317_ ), .B1(_06339_ ), .B2(_06343_ ), .ZN(_06344_ ) );
BUF_X4 _14428_ ( .A(_03911_ ), .Z(_06345_ ) );
NAND3_X1 _14429_ ( .A1(_06336_ ), .A2(_06344_ ), .A3(_06345_ ), .ZN(_06346_ ) );
AND3_X1 _14430_ ( .A1(_06140_ ), .A2(_03084_ ), .A3(_06143_ ), .ZN(_06347_ ) );
OR3_X1 _14431_ ( .A1(_06347_ ), .A2(_06318_ ), .A3(_06166_ ), .ZN(_06348_ ) );
BUF_X4 _14432_ ( .A(_06172_ ), .Z(_06349_ ) );
AND3_X1 _14433_ ( .A1(_06306_ ), .A2(_03005_ ), .A3(_06307_ ), .ZN(_06350_ ) );
AOI21_X1 _14434_ ( .A(_01918_ ), .B1(_06140_ ), .B2(_06143_ ), .ZN(_06351_ ) );
BUF_X2 _14435_ ( .A(_06150_ ), .Z(_06352_ ) );
OR3_X1 _14436_ ( .A1(_06350_ ), .A2(_06351_ ), .A3(_06352_ ), .ZN(_06353_ ) );
NAND3_X1 _14437_ ( .A1(_06348_ ), .A2(_06349_ ), .A3(_06353_ ), .ZN(_06354_ ) );
AND3_X1 _14438_ ( .A1(_06326_ ), .A2(_02953_ ), .A3(_06327_ ), .ZN(_06355_ ) );
AOI21_X1 _14439_ ( .A(_01942_ ), .B1(_06326_ ), .B2(_06327_ ), .ZN(_06356_ ) );
OAI21_X1 _14440_ ( .A(_06334_ ), .B1(_06355_ ), .B2(_06356_ ), .ZN(_06357_ ) );
AND3_X1 _14441_ ( .A1(_06306_ ), .A2(_03135_ ), .A3(_06307_ ), .ZN(_06358_ ) );
AOI21_X1 _14442_ ( .A(_02309_ ), .B1(_06326_ ), .B2(_06327_ ), .ZN(_06359_ ) );
OAI21_X1 _14443_ ( .A(_06329_ ), .B1(_06358_ ), .B2(_06359_ ), .ZN(_06360_ ) );
NAND2_X1 _14444_ ( .A1(_06357_ ), .A2(_06360_ ), .ZN(_06361_ ) );
NAND2_X1 _14445_ ( .A1(_06361_ ), .A2(_06325_ ), .ZN(_06362_ ) );
AND2_X1 _14446_ ( .A1(_06354_ ), .A2(_06362_ ), .ZN(_06363_ ) );
BUF_X4 _14447_ ( .A(_06323_ ), .Z(_06364_ ) );
OAI211_X1 _14448_ ( .A(_06178_ ), .B(_06346_ ), .C1(_06363_ ), .C2(_06364_ ), .ZN(_06365_ ) );
AOI21_X1 _14449_ ( .A(_06305_ ), .B1(_06324_ ), .B2(_06365_ ), .ZN(_06366_ ) );
BUF_X4 _14450_ ( .A(_03723_ ), .Z(_06367_ ) );
BUF_X4 _14451_ ( .A(_03986_ ), .Z(_06368_ ) );
AOI221_X4 _14452_ ( .A(_06366_ ), .B1(_03827_ ), .B2(_06367_ ), .C1(_03798_ ), .C2(_06368_ ), .ZN(_06369_ ) );
NAND3_X1 _14453_ ( .A1(_06246_ ), .A2(_06304_ ), .A3(_06369_ ), .ZN(_06370_ ) );
OAI21_X1 _14454_ ( .A(_06128_ ), .B1(_06127_ ), .B2(_06114_ ), .ZN(_06371_ ) );
NOR2_X1 _14455_ ( .A1(_04086_ ), .A2(\ID_EX_typ [2] ), .ZN(_06372_ ) );
OAI211_X1 _14456_ ( .A(_06372_ ), .B(_04073_ ), .C1(_03728_ ), .C2(_02832_ ), .ZN(_06373_ ) );
AND2_X1 _14457_ ( .A1(_06371_ ), .A2(_06373_ ), .ZN(_06374_ ) );
NOR2_X2 _14458_ ( .A1(_06374_ ), .A2(_06132_ ), .ZN(_06375_ ) );
INV_X1 _14459_ ( .A(_06375_ ), .ZN(_06376_ ) );
BUF_X4 _14460_ ( .A(_06376_ ), .Z(_06377_ ) );
AOI21_X1 _14461_ ( .A(_06134_ ), .B1(_06370_ ), .B2(_06377_ ), .ZN(_06378_ ) );
OAI21_X1 _14462_ ( .A(_06030_ ), .B1(_04947_ ), .B2(_01655_ ), .ZN(_06379_ ) );
OAI21_X1 _14463_ ( .A(_06113_ ), .B1(_06378_ ), .B2(_06379_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
NAND3_X1 _14464_ ( .A1(_04179_ ), .A2(_05879_ ), .A3(_04184_ ), .ZN(_06380_ ) );
BUF_X4 _14465_ ( .A(_06131_ ), .Z(_06381_ ) );
AND2_X2 _14466_ ( .A1(_06127_ ), .A2(_06115_ ), .ZN(_06382_ ) );
INV_X2 _14467_ ( .A(_06382_ ), .ZN(_06383_ ) );
OAI22_X1 _14468_ ( .A1(_04193_ ), .A2(_06118_ ), .B1(_01870_ ), .B2(_06383_ ), .ZN(_06384_ ) );
OR2_X1 _14469_ ( .A1(_06121_ ), .A2(_03085_ ), .ZN(_06385_ ) );
INV_X1 _14470_ ( .A(_06125_ ), .ZN(_06386_ ) );
BUF_X4 _14471_ ( .A(_06386_ ), .Z(_06387_ ) );
AOI21_X1 _14472_ ( .A(_06387_ ), .B1(_06121_ ), .B2(_03085_ ), .ZN(_06388_ ) );
AND2_X1 _14473_ ( .A1(_06385_ ), .A2(_06388_ ), .ZN(_06389_ ) );
OAI21_X1 _14474_ ( .A(_06381_ ), .B1(_06384_ ), .B2(_06389_ ), .ZN(_06390_ ) );
BUF_X2 _14475_ ( .A(_02840_ ), .Z(_06391_ ) );
NAND2_X1 _14476_ ( .A1(_06390_ ), .A2(_06391_ ), .ZN(_06392_ ) );
INV_X1 _14477_ ( .A(_06247_ ), .ZN(_06393_ ) );
BUF_X2 _14478_ ( .A(_06393_ ), .Z(_06394_ ) );
BUF_X2 _14479_ ( .A(_06318_ ), .Z(_06395_ ) );
INV_X1 _14480_ ( .A(_06147_ ), .ZN(_06396_ ) );
OAI21_X1 _14481_ ( .A(_06349_ ), .B1(_06395_ ), .B2(_06396_ ), .ZN(_06397_ ) );
AND3_X1 _14482_ ( .A1(_06288_ ), .A2(_06300_ ), .A3(_06397_ ), .ZN(_06398_ ) );
OAI22_X1 _14483_ ( .A1(_06398_ ), .A2(_06292_ ), .B1(_06290_ ), .B2(_06293_ ), .ZN(_06399_ ) );
BUF_X2 _14484_ ( .A(_03918_ ), .Z(_06400_ ) );
BUF_X2 _14485_ ( .A(_03920_ ), .Z(_06401_ ) );
AND3_X1 _14486_ ( .A1(_06400_ ), .A2(_02403_ ), .A3(_06401_ ), .ZN(_06402_ ) );
AOI21_X1 _14487_ ( .A(_01869_ ), .B1(_06400_ ), .B2(_06401_ ), .ZN(_06403_ ) );
OAI21_X1 _14488_ ( .A(_06145_ ), .B1(_06402_ ), .B2(_06403_ ), .ZN(_06404_ ) );
AND3_X1 _14489_ ( .A1(_06138_ ), .A2(_03058_ ), .A3(_06141_ ), .ZN(_06405_ ) );
AOI21_X1 _14490_ ( .A(_01793_ ), .B1(_06400_ ), .B2(_06401_ ), .ZN(_06406_ ) );
OAI21_X1 _14491_ ( .A(_06157_ ), .B1(_06405_ ), .B2(_06406_ ), .ZN(_06407_ ) );
AOI21_X1 _14492_ ( .A(_06154_ ), .B1(_06404_ ), .B2(_06407_ ), .ZN(_06408_ ) );
AND3_X1 _14493_ ( .A1(_06138_ ), .A2(_03476_ ), .A3(_06141_ ), .ZN(_06409_ ) );
AOI21_X1 _14494_ ( .A(_02432_ ), .B1(_06138_ ), .B2(_06141_ ), .ZN(_06410_ ) );
OAI21_X1 _14495_ ( .A(_06145_ ), .B1(_06409_ ), .B2(_06410_ ), .ZN(_06411_ ) );
AND3_X1 _14496_ ( .A1(_06138_ ), .A2(_03763_ ), .A3(_06141_ ), .ZN(_06412_ ) );
AOI21_X1 _14497_ ( .A(_02510_ ), .B1(_06138_ ), .B2(_06141_ ), .ZN(_06413_ ) );
OAI21_X1 _14498_ ( .A(_06157_ ), .B1(_06412_ ), .B2(_06413_ ), .ZN(_06414_ ) );
AOI21_X1 _14499_ ( .A(_06316_ ), .B1(_06411_ ), .B2(_06414_ ), .ZN(_06415_ ) );
NOR2_X1 _14500_ ( .A1(_06408_ ), .A2(_06415_ ), .ZN(_06416_ ) );
AND3_X1 _14501_ ( .A1(_03918_ ), .A2(_03738_ ), .A3(_03920_ ), .ZN(_06417_ ) );
AOI21_X1 _14502_ ( .A(_01765_ ), .B1(_03918_ ), .B2(_03920_ ), .ZN(_06418_ ) );
NOR2_X1 _14503_ ( .A1(_06417_ ), .A2(_06418_ ), .ZN(_06419_ ) );
MUX2_X1 _14504_ ( .A(_02571_ ), .B(_06137_ ), .S(_03921_ ), .Z(_06420_ ) );
MUX2_X1 _14505_ ( .A(_06419_ ), .B(_06420_ ), .S(_06157_ ), .Z(_06421_ ) );
BUF_X4 _14506_ ( .A(_06172_ ), .Z(_06422_ ) );
AND2_X1 _14507_ ( .A1(_06421_ ), .A2(_06422_ ), .ZN(_06423_ ) );
MUX2_X1 _14508_ ( .A(_06416_ ), .B(_06423_ ), .S(_06323_ ), .Z(_06424_ ) );
BUF_X2 _14509_ ( .A(_06322_ ), .Z(_06425_ ) );
NAND2_X1 _14510_ ( .A1(_06424_ ), .A2(_06425_ ), .ZN(_06426_ ) );
AOI21_X1 _14511_ ( .A(_06394_ ), .B1(_06399_ ), .B2(_06426_ ), .ZN(_06427_ ) );
AND3_X1 _14512_ ( .A1(_06424_ ), .A2(_06425_ ), .A3(_06180_ ), .ZN(_06428_ ) );
AOI21_X1 _14513_ ( .A(_03646_ ), .B1(_06326_ ), .B2(_06327_ ), .ZN(_06429_ ) );
AND2_X1 _14514_ ( .A1(_06429_ ), .A2(_06342_ ), .ZN(_06430_ ) );
INV_X1 _14515_ ( .A(_06430_ ), .ZN(_06431_ ) );
NOR2_X1 _14516_ ( .A1(_06147_ ), .A2(_02014_ ), .ZN(_06432_ ) );
AOI21_X1 _14517_ ( .A(_02045_ ), .B1(_06139_ ), .B2(_06142_ ), .ZN(_06433_ ) );
NOR3_X1 _14518_ ( .A1(_06432_ ), .A2(_06352_ ), .A3(_06433_ ), .ZN(_06434_ ) );
AND3_X1 _14519_ ( .A1(_06400_ ), .A2(_03904_ ), .A3(_06401_ ), .ZN(_06435_ ) );
AOI21_X1 _14520_ ( .A(_02118_ ), .B1(_06400_ ), .B2(_06401_ ), .ZN(_06436_ ) );
NOR3_X1 _14521_ ( .A1(_06435_ ), .A2(_06309_ ), .A3(_06436_ ), .ZN(_06437_ ) );
NOR2_X1 _14522_ ( .A1(_06434_ ), .A2(_06437_ ), .ZN(_06438_ ) );
MUX2_X1 _14523_ ( .A(_06431_ ), .B(_06438_ ), .S(_06422_ ), .Z(_06439_ ) );
NOR2_X1 _14524_ ( .A1(_06439_ ), .A2(_06345_ ), .ZN(_06440_ ) );
OAI21_X1 _14525_ ( .A(_04070_ ), .B1(_06440_ ), .B2(_06178_ ), .ZN(_06441_ ) );
INV_X1 _14526_ ( .A(_06177_ ), .ZN(_06442_ ) );
BUF_X2 _14527_ ( .A(_06442_ ), .Z(_06443_ ) );
AND3_X1 _14528_ ( .A1(_06139_ ), .A2(_03214_ ), .A3(_06142_ ), .ZN(_06444_ ) );
INV_X1 _14529_ ( .A(_06444_ ), .ZN(_06445_ ) );
AOI21_X1 _14530_ ( .A(_02332_ ), .B1(_06139_ ), .B2(_06142_ ), .ZN(_06446_ ) );
INV_X1 _14531_ ( .A(_06446_ ), .ZN(_06447_ ) );
NAND3_X1 _14532_ ( .A1(_06445_ ), .A2(_06329_ ), .A3(_06447_ ), .ZN(_06448_ ) );
AND3_X1 _14533_ ( .A1(_06139_ ), .A2(_03954_ ), .A3(_06142_ ), .ZN(_06449_ ) );
INV_X1 _14534_ ( .A(_06449_ ), .ZN(_06450_ ) );
AOI21_X1 _14535_ ( .A(_01965_ ), .B1(_06138_ ), .B2(_06141_ ), .ZN(_06451_ ) );
INV_X1 _14536_ ( .A(_06451_ ), .ZN(_06452_ ) );
NAND3_X1 _14537_ ( .A1(_06450_ ), .A2(_06334_ ), .A3(_06452_ ), .ZN(_06453_ ) );
AOI21_X1 _14538_ ( .A(_06422_ ), .B1(_06448_ ), .B2(_06453_ ), .ZN(_06454_ ) );
AND3_X1 _14539_ ( .A1(_06138_ ), .A2(_02977_ ), .A3(_06141_ ), .ZN(_06455_ ) );
OAI21_X1 _14540_ ( .A(_06352_ ), .B1(_06455_ ), .B2(_06403_ ), .ZN(_06456_ ) );
AND3_X1 _14541_ ( .A1(_06326_ ), .A2(_02922_ ), .A3(_06327_ ), .ZN(_06457_ ) );
AOI21_X1 _14542_ ( .A(_01895_ ), .B1(_06138_ ), .B2(_06141_ ), .ZN(_06458_ ) );
OAI21_X1 _14543_ ( .A(_06318_ ), .B1(_06457_ ), .B2(_06458_ ), .ZN(_06459_ ) );
AND3_X1 _14544_ ( .A1(_06456_ ), .A2(_06459_ ), .A3(_06316_ ), .ZN(_06460_ ) );
OR3_X1 _14545_ ( .A1(_06454_ ), .A2(_06460_ ), .A3(_06323_ ), .ZN(_06461_ ) );
AOI21_X1 _14546_ ( .A(_02249_ ), .B1(_06400_ ), .B2(_06401_ ), .ZN(_06462_ ) );
INV_X1 _14547_ ( .A(_06462_ ), .ZN(_06463_ ) );
OAI211_X1 _14548_ ( .A(_06463_ ), .B(_06329_ ), .C1(_02225_ ), .C2(_06147_ ), .ZN(_06464_ ) );
AND3_X1 _14549_ ( .A1(_06400_ ), .A2(_03241_ ), .A3(_06401_ ), .ZN(_06465_ ) );
INV_X1 _14550_ ( .A(_06465_ ), .ZN(_06466_ ) );
AOI21_X1 _14551_ ( .A(_02380_ ), .B1(_06139_ ), .B2(_06142_ ), .ZN(_06467_ ) );
INV_X1 _14552_ ( .A(_06467_ ), .ZN(_06468_ ) );
NAND3_X1 _14553_ ( .A1(_06466_ ), .A2(_06334_ ), .A3(_06468_ ), .ZN(_06469_ ) );
AND3_X1 _14554_ ( .A1(_06464_ ), .A2(_06469_ ), .A3(_06422_ ), .ZN(_06470_ ) );
NOR2_X1 _14555_ ( .A1(_06147_ ), .A2(_02096_ ), .ZN(_06471_ ) );
AOI21_X1 _14556_ ( .A(_02171_ ), .B1(_06400_ ), .B2(_06401_ ), .ZN(_06472_ ) );
OAI21_X1 _14557_ ( .A(_06329_ ), .B1(_06471_ ), .B2(_06472_ ), .ZN(_06473_ ) );
AND3_X1 _14558_ ( .A1(_06400_ ), .A2(_03342_ ), .A3(_06401_ ), .ZN(_06474_ ) );
AOI21_X1 _14559_ ( .A(_02202_ ), .B1(_06138_ ), .B2(_06141_ ), .ZN(_06475_ ) );
OAI21_X1 _14560_ ( .A(_06334_ ), .B1(_06474_ ), .B2(_06475_ ), .ZN(_06476_ ) );
AOI21_X1 _14561_ ( .A(_06349_ ), .B1(_06473_ ), .B2(_06476_ ), .ZN(_06477_ ) );
OAI21_X1 _14562_ ( .A(_06345_ ), .B1(_06470_ ), .B2(_06477_ ), .ZN(_06478_ ) );
AOI21_X1 _14563_ ( .A(_06443_ ), .B1(_06461_ ), .B2(_06478_ ), .ZN(_06479_ ) );
NOR2_X1 _14564_ ( .A1(_06441_ ), .A2(_06479_ ), .ZN(_06480_ ) );
OR3_X1 _14565_ ( .A1(_06427_ ), .A2(_06428_ ), .A3(_06480_ ), .ZN(_06481_ ) );
OAI21_X1 _14566_ ( .A(_06245_ ), .B1(_06238_ ), .B2(_06239_ ), .ZN(_06482_ ) );
AOI21_X1 _14567_ ( .A(_06482_ ), .B1(_06239_ ), .B2(_06238_ ), .ZN(_06483_ ) );
NAND3_X1 _14568_ ( .A1(_03791_ ), .A2(_03084_ ), .A3(_03792_ ), .ZN(_06484_ ) );
NAND3_X1 _14569_ ( .A1(_06182_ ), .A2(_06484_ ), .A3(_06368_ ), .ZN(_06485_ ) );
BUF_X4 _14570_ ( .A(_04075_ ), .Z(_06486_ ) );
NAND2_X1 _14571_ ( .A1(_06484_ ), .A2(_06486_ ), .ZN(_06487_ ) );
CLKBUF_X2 _14572_ ( .A(_03724_ ), .Z(_06488_ ) );
OR3_X1 _14573_ ( .A1(_03793_ ), .A2(_03084_ ), .A3(_06488_ ), .ZN(_06489_ ) );
NAND3_X1 _14574_ ( .A1(_06485_ ), .A2(_06487_ ), .A3(_06489_ ), .ZN(_06490_ ) );
OR3_X1 _14575_ ( .A1(_06481_ ), .A2(_06483_ ), .A3(_06490_ ), .ZN(_06491_ ) );
AOI21_X1 _14576_ ( .A(_06392_ ), .B1(_06491_ ), .B2(_06377_ ), .ZN(_06492_ ) );
OAI21_X1 _14577_ ( .A(_06030_ ), .B1(_04188_ ), .B2(_01655_ ), .ZN(_06493_ ) );
OAI21_X1 _14578_ ( .A(_06380_ ), .B1(_06492_ ), .B2(_06493_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OR2_X1 _14579_ ( .A1(_04211_ ), .A2(_05891_ ), .ZN(_06494_ ) );
AND2_X1 _14580_ ( .A1(_03004_ ), .A2(_01895_ ), .ZN(_06495_ ) );
INV_X1 _14581_ ( .A(_04025_ ), .ZN(_06496_ ) );
AND2_X1 _14582_ ( .A1(_06496_ ), .A2(_02955_ ), .ZN(_06497_ ) );
OR3_X1 _14583_ ( .A1(_06497_ ), .A2(_04050_ ), .A3(_04052_ ), .ZN(_06498_ ) );
AOI21_X1 _14584_ ( .A(_06495_ ), .B1(_06498_ ), .B2(_03006_ ), .ZN(_06499_ ) );
XNOR2_X1 _14585_ ( .A(_06499_ ), .B(_02978_ ), .ZN(_06500_ ) );
BUF_X2 _14586_ ( .A(_06125_ ), .Z(_06501_ ) );
NAND2_X1 _14587_ ( .A1(_06500_ ), .A2(_06501_ ), .ZN(_06502_ ) );
OR2_X1 _14588_ ( .A1(_04220_ ), .A2(_06117_ ), .ZN(_06503_ ) );
NAND3_X1 _14589_ ( .A1(_06127_ ), .A2(\ID_EX_imm [19] ), .A3(_06128_ ), .ZN(_06504_ ) );
AND3_X1 _14590_ ( .A1(_06502_ ), .A2(_06503_ ), .A3(_06504_ ), .ZN(_06505_ ) );
OAI21_X1 _14591_ ( .A(_04161_ ), .B1(_06505_ ), .B2(_06133_ ), .ZN(_06506_ ) );
OR3_X1 _14592_ ( .A1(_03922_ ), .A2(_06146_ ), .A3(_06319_ ), .ZN(_06507_ ) );
OR3_X1 _14593_ ( .A1(_06312_ ), .A2(_06158_ ), .A3(_06313_ ), .ZN(_06508_ ) );
AOI21_X1 _14594_ ( .A(_06297_ ), .B1(_06507_ ), .B2(_06508_ ), .ZN(_06509_ ) );
BUF_X2 _14595_ ( .A(_06175_ ), .Z(_06510_ ) );
AND2_X1 _14596_ ( .A1(_06509_ ), .A2(_06510_ ), .ZN(_06511_ ) );
OAI21_X1 _14597_ ( .A(_04070_ ), .B1(_06511_ ), .B2(_06178_ ), .ZN(_06512_ ) );
NOR3_X1 _14598_ ( .A1(_06332_ ), .A2(_06309_ ), .A3(_06333_ ), .ZN(_06513_ ) );
NOR3_X1 _14599_ ( .A1(_06308_ ), .A2(_06310_ ), .A3(_06151_ ), .ZN(_06514_ ) );
NOR2_X1 _14600_ ( .A1(_06513_ ), .A2(_06514_ ), .ZN(_06515_ ) );
NAND2_X1 _14601_ ( .A1(_06515_ ), .A2(_06325_ ), .ZN(_06516_ ) );
NOR3_X1 _14602_ ( .A1(_06340_ ), .A2(_06318_ ), .A3(_06341_ ), .ZN(_06517_ ) );
NOR3_X1 _14603_ ( .A1(_06328_ ), .A2(_06330_ ), .A3(_06352_ ), .ZN(_06518_ ) );
NOR2_X1 _14604_ ( .A1(_06517_ ), .A2(_06518_ ), .ZN(_06519_ ) );
NAND2_X1 _14605_ ( .A1(_06519_ ), .A2(_06349_ ), .ZN(_06520_ ) );
NAND2_X1 _14606_ ( .A1(_06516_ ), .A2(_06520_ ), .ZN(_06521_ ) );
OAI21_X1 _14607_ ( .A(_06342_ ), .B1(_06350_ ), .B2(_06351_ ), .ZN(_06522_ ) );
OAI21_X1 _14608_ ( .A(_06318_ ), .B1(_06355_ ), .B2(_06356_ ), .ZN(_06523_ ) );
NAND2_X1 _14609_ ( .A1(_06522_ ), .A2(_06523_ ), .ZN(_06524_ ) );
NOR3_X1 _14610_ ( .A1(_06358_ ), .A2(_06309_ ), .A3(_06359_ ), .ZN(_06525_ ) );
NOR3_X1 _14611_ ( .A1(_06337_ ), .A2(_06338_ ), .A3(_06151_ ), .ZN(_06526_ ) );
NOR2_X1 _14612_ ( .A1(_06525_ ), .A2(_06526_ ), .ZN(_06527_ ) );
MUX2_X1 _14613_ ( .A(_06524_ ), .B(_06527_ ), .S(_06154_ ), .Z(_06528_ ) );
MUX2_X1 _14614_ ( .A(_06521_ ), .B(_06528_ ), .S(_06510_ ), .Z(_06529_ ) );
BUF_X2 _14615_ ( .A(_06322_ ), .Z(_06530_ ) );
AOI21_X1 _14616_ ( .A(_06512_ ), .B1(_06529_ ), .B2(_06530_ ), .ZN(_06531_ ) );
NOR3_X1 _14617_ ( .A1(_06169_ ), .A2(_06158_ ), .A3(_06170_ ), .ZN(_06532_ ) );
NOR3_X1 _14618_ ( .A1(_06156_ ), .A2(_06159_ ), .A3(_06150_ ), .ZN(_06533_ ) );
OAI21_X1 _14619_ ( .A(_03909_ ), .B1(_06532_ ), .B2(_06533_ ), .ZN(_06534_ ) );
NOR3_X1 _14620_ ( .A1(_06347_ ), .A2(_06158_ ), .A3(_06351_ ), .ZN(_06535_ ) );
NOR3_X1 _14621_ ( .A1(_06165_ ), .A2(_06166_ ), .A3(_06150_ ), .ZN(_06536_ ) );
OAI21_X1 _14622_ ( .A(_06172_ ), .B1(_06535_ ), .B2(_06536_ ), .ZN(_06537_ ) );
NAND2_X1 _14623_ ( .A1(_06534_ ), .A2(_06537_ ), .ZN(_06538_ ) );
NAND2_X1 _14624_ ( .A1(_06538_ ), .A2(_06175_ ), .ZN(_06539_ ) );
AND2_X1 _14625_ ( .A1(_06152_ ), .A2(_06150_ ), .ZN(_06540_ ) );
INV_X1 _14626_ ( .A(_06540_ ), .ZN(_06541_ ) );
AOI21_X1 _14627_ ( .A(_06150_ ), .B1(_06144_ ), .B2(_06148_ ), .ZN(_06542_ ) );
NOR3_X1 _14628_ ( .A1(_06161_ ), .A2(_06158_ ), .A3(_06162_ ), .ZN(_06543_ ) );
NOR2_X1 _14629_ ( .A1(_06542_ ), .A2(_06543_ ), .ZN(_06544_ ) );
MUX2_X1 _14630_ ( .A(_06541_ ), .B(_06544_ ), .S(_06172_ ), .Z(_06545_ ) );
BUF_X4 _14631_ ( .A(_06175_ ), .Z(_06546_ ) );
OAI21_X1 _14632_ ( .A(_06539_ ), .B1(_06545_ ), .B2(_06546_ ), .ZN(_06547_ ) );
AND2_X1 _14633_ ( .A1(_06547_ ), .A2(_06177_ ), .ZN(_06548_ ) );
AND2_X2 _14634_ ( .A1(_06290_ ), .A2(_06292_ ), .ZN(_06549_ ) );
XNOR2_X1 _14635_ ( .A(_06250_ ), .B(_06316_ ), .ZN(_06550_ ) );
AND4_X1 _14636_ ( .A1(_06300_ ), .A2(_06288_ ), .A3(_06550_ ), .A4(_06289_ ), .ZN(_06551_ ) );
OR3_X1 _14637_ ( .A1(_06549_ ), .A2(_06551_ ), .A3(_06548_ ), .ZN(_06552_ ) );
AOI221_X4 _14638_ ( .A(_06531_ ), .B1(_06181_ ), .B2(_06548_ ), .C1(_06552_ ), .C2(_06248_ ), .ZN(_06553_ ) );
AND2_X1 _14639_ ( .A1(_06208_ ), .A2(_06227_ ), .ZN(_06554_ ) );
INV_X1 _14640_ ( .A(_03807_ ), .ZN(_06555_ ) );
INV_X1 _14641_ ( .A(_03958_ ), .ZN(_06556_ ) );
OR3_X1 _14642_ ( .A1(_06554_ ), .A2(_06555_ ), .A3(_06556_ ), .ZN(_06557_ ) );
AOI21_X1 _14643_ ( .A(_06232_ ), .B1(_03807_ ), .B2(_06230_ ), .ZN(_06558_ ) );
AOI21_X1 _14644_ ( .A(_03820_ ), .B1(_06557_ ), .B2(_06558_ ), .ZN(_06559_ ) );
OR3_X1 _14645_ ( .A1(_06559_ ), .A2(_03814_ ), .A3(_06235_ ), .ZN(_06560_ ) );
BUF_X2 _14646_ ( .A(_06245_ ), .Z(_06561_ ) );
OAI21_X1 _14647_ ( .A(_03814_ ), .B1(_06559_ ), .B2(_06235_ ), .ZN(_06562_ ) );
NAND3_X1 _14648_ ( .A1(_06560_ ), .A2(_06561_ ), .A3(_06562_ ), .ZN(_06563_ ) );
AOI21_X1 _14649_ ( .A(_01918_ ), .B1(_03800_ ), .B2(_03801_ ), .ZN(_06564_ ) );
BUF_X4 _14650_ ( .A(_06135_ ), .Z(_06565_ ) );
OAI22_X1 _14651_ ( .A1(_06234_ ), .A2(_06488_ ), .B1(_06564_ ), .B2(_06565_ ), .ZN(_06566_ ) );
BUF_X2 _14652_ ( .A(_06368_ ), .Z(_06567_ ) );
AOI21_X1 _14653_ ( .A(_06566_ ), .B1(_03814_ ), .B2(_06567_ ), .ZN(_06568_ ) );
NAND3_X1 _14654_ ( .A1(_06553_ ), .A2(_06563_ ), .A3(_06568_ ), .ZN(_06569_ ) );
AOI21_X1 _14655_ ( .A(_06506_ ), .B1(_06569_ ), .B2(_06377_ ), .ZN(_06570_ ) );
OAI21_X1 _14656_ ( .A(_06030_ ), .B1(_04214_ ), .B2(_01655_ ), .ZN(_06571_ ) );
OAI21_X1 _14657_ ( .A(_06494_ ), .B1(_06570_ ), .B2(_06571_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
INV_X1 _14658_ ( .A(_05911_ ), .ZN(_06572_ ) );
BUF_X4 _14659_ ( .A(_06132_ ), .Z(_06573_ ) );
AOI21_X1 _14660_ ( .A(_06386_ ), .B1(_06498_ ), .B2(_03006_ ), .ZN(_06574_ ) );
OAI21_X1 _14661_ ( .A(_06574_ ), .B1(_03006_ ), .B2(_06498_ ), .ZN(_06575_ ) );
BUF_X4 _14662_ ( .A(_06116_ ), .Z(_06576_ ) );
BUF_X4 _14663_ ( .A(_06382_ ), .Z(_06577_ ) );
AOI22_X1 _14664_ ( .A1(_04245_ ), .A2(_06576_ ), .B1(\ID_EX_imm [18] ), .B2(_06577_ ), .ZN(_06578_ ) );
AOI21_X1 _14665_ ( .A(_06573_ ), .B1(_06575_ ), .B2(_06578_ ), .ZN(_06579_ ) );
OR2_X1 _14666_ ( .A1(_06579_ ), .A2(_01650_ ), .ZN(_06580_ ) );
NOR2_X1 _14667_ ( .A1(_06290_ ), .A2(_06293_ ), .ZN(_06581_ ) );
AND2_X1 _14668_ ( .A1(_06288_ ), .A2(_06550_ ), .ZN(_06582_ ) );
INV_X1 _14669_ ( .A(_06582_ ), .ZN(_06583_ ) );
NOR2_X1 _14670_ ( .A1(_06395_ ), .A2(_06147_ ), .ZN(_06584_ ) );
OR3_X1 _14671_ ( .A1(_06583_ ), .A2(_06584_ ), .A3(_06299_ ), .ZN(_06585_ ) );
AOI21_X1 _14672_ ( .A(_06581_ ), .B1(_06585_ ), .B2(_06295_ ), .ZN(_06586_ ) );
NOR3_X1 _14673_ ( .A1(_06405_ ), .A2(_06318_ ), .A3(_06406_ ), .ZN(_06587_ ) );
NOR3_X1 _14674_ ( .A1(_06409_ ), .A2(_06410_ ), .A3(_06352_ ), .ZN(_06588_ ) );
OAI21_X1 _14675_ ( .A(_06297_ ), .B1(_06587_ ), .B2(_06588_ ), .ZN(_06589_ ) );
OAI21_X1 _14676_ ( .A(_06342_ ), .B1(_06455_ ), .B2(_06458_ ), .ZN(_06590_ ) );
OAI21_X1 _14677_ ( .A(_06318_ ), .B1(_06402_ ), .B2(_06403_ ), .ZN(_06591_ ) );
NAND3_X1 _14678_ ( .A1(_06590_ ), .A2(_06591_ ), .A3(_06316_ ), .ZN(_06592_ ) );
AND2_X1 _14679_ ( .A1(_06589_ ), .A2(_06592_ ), .ZN(_06593_ ) );
NAND3_X1 _14680_ ( .A1(_06420_ ), .A2(_06154_ ), .A3(_06334_ ), .ZN(_06594_ ) );
NOR3_X1 _14681_ ( .A1(_06412_ ), .A2(_06309_ ), .A3(_06413_ ), .ZN(_06595_ ) );
NOR3_X1 _14682_ ( .A1(_06417_ ), .A2(_06418_ ), .A3(_06151_ ), .ZN(_06596_ ) );
OAI21_X1 _14683_ ( .A(_06316_ ), .B1(_06595_ ), .B2(_06596_ ), .ZN(_06597_ ) );
AND2_X1 _14684_ ( .A1(_06594_ ), .A2(_06597_ ), .ZN(_06598_ ) );
MUX2_X1 _14685_ ( .A(_06593_ ), .B(_06598_ ), .S(_06345_ ), .Z(_06599_ ) );
BUF_X2 _14686_ ( .A(_06443_ ), .Z(_06600_ ) );
NOR2_X1 _14687_ ( .A1(_06599_ ), .A2(_06600_ ), .ZN(_06601_ ) );
OAI21_X1 _14688_ ( .A(_06249_ ), .B1(_06586_ ), .B2(_06601_ ), .ZN(_06602_ ) );
AOI21_X1 _14689_ ( .A(_06565_ ), .B1(_03818_ ), .B2(_03005_ ), .ZN(_06603_ ) );
OAI21_X1 _14690_ ( .A(_06157_ ), .B1(_06396_ ), .B2(_03646_ ), .ZN(_06604_ ) );
AOI21_X1 _14691_ ( .A(_06433_ ), .B1(_06396_ ), .B2(_02041_ ), .ZN(_06605_ ) );
OAI21_X1 _14692_ ( .A(_06604_ ), .B1(_06605_ ), .B2(_06158_ ), .ZN(_06606_ ) );
BUF_X4 _14693_ ( .A(_06325_ ), .Z(_06607_ ) );
NOR2_X1 _14694_ ( .A1(_06606_ ), .A2(_06607_ ), .ZN(_06608_ ) );
BUF_X2 _14695_ ( .A(_06510_ ), .Z(_06609_ ) );
AND2_X1 _14696_ ( .A1(_06608_ ), .A2(_06609_ ), .ZN(_06610_ ) );
OAI21_X1 _14697_ ( .A(_04070_ ), .B1(_06610_ ), .B2(_06530_ ), .ZN(_06611_ ) );
OAI21_X1 _14698_ ( .A(_06334_ ), .B1(_06457_ ), .B2(_06458_ ), .ZN(_06612_ ) );
OAI21_X1 _14699_ ( .A(_06395_ ), .B1(_06449_ ), .B2(_06451_ ), .ZN(_06613_ ) );
NAND2_X1 _14700_ ( .A1(_06612_ ), .A2(_06613_ ), .ZN(_06614_ ) );
OAI21_X1 _14701_ ( .A(_06352_ ), .B1(_06444_ ), .B2(_06446_ ), .ZN(_06615_ ) );
OAI21_X1 _14702_ ( .A(_06309_ ), .B1(_06465_ ), .B2(_06467_ ), .ZN(_06616_ ) );
NAND2_X1 _14703_ ( .A1(_06615_ ), .A2(_06616_ ), .ZN(_06617_ ) );
BUF_X4 _14704_ ( .A(_06297_ ), .Z(_06618_ ) );
MUX2_X1 _14705_ ( .A(_06614_ ), .B(_06617_ ), .S(_06618_ ), .Z(_06619_ ) );
BUF_X4 _14706_ ( .A(_06422_ ), .Z(_06620_ ) );
AND3_X1 _14707_ ( .A1(_06400_ ), .A2(_03292_ ), .A3(_06401_ ), .ZN(_06621_ ) );
NOR3_X1 _14708_ ( .A1(_06621_ ), .A2(_06309_ ), .A3(_06462_ ), .ZN(_06622_ ) );
NOR3_X1 _14709_ ( .A1(_06474_ ), .A2(_06475_ ), .A3(_06146_ ), .ZN(_06623_ ) );
OAI21_X1 _14710_ ( .A(_06620_ ), .B1(_06622_ ), .B2(_06623_ ), .ZN(_06624_ ) );
NOR3_X1 _14711_ ( .A1(_06471_ ), .A2(_06157_ ), .A3(_06472_ ), .ZN(_06625_ ) );
NOR3_X1 _14712_ ( .A1(_06435_ ), .A2(_06436_ ), .A3(_06150_ ), .ZN(_06626_ ) );
OAI21_X1 _14713_ ( .A(_06618_ ), .B1(_06625_ ), .B2(_06626_ ), .ZN(_06627_ ) );
AND2_X1 _14714_ ( .A1(_06624_ ), .A2(_06627_ ), .ZN(_06628_ ) );
MUX2_X1 _14715_ ( .A(_06619_ ), .B(_06628_ ), .S(_06364_ ), .Z(_06629_ ) );
BUF_X2 _14716_ ( .A(_06425_ ), .Z(_06630_ ) );
AOI21_X1 _14717_ ( .A(_06611_ ), .B1(_06629_ ), .B2(_06630_ ), .ZN(_06631_ ) );
AOI211_X1 _14718_ ( .A(_06603_ ), .B(_06631_ ), .C1(_03819_ ), .C2(_06567_ ), .ZN(_06632_ ) );
AND3_X1 _14719_ ( .A1(_06557_ ), .A2(_03820_ ), .A3(_06558_ ), .ZN(_06633_ ) );
INV_X1 _14720_ ( .A(_06245_ ), .ZN(_06634_ ) );
NOR3_X1 _14721_ ( .A1(_06633_ ), .A2(_06559_ ), .A3(_06634_ ), .ZN(_06635_ ) );
AOI221_X4 _14722_ ( .A(_06635_ ), .B1(_06235_ ), .B2(_06367_ ), .C1(_06181_ ), .C2(_06601_ ), .ZN(_06636_ ) );
NAND3_X1 _14723_ ( .A1(_06602_ ), .A2(_06632_ ), .A3(_06636_ ), .ZN(_06637_ ) );
AOI21_X1 _14724_ ( .A(_06580_ ), .B1(_06637_ ), .B2(_06377_ ), .ZN(_06638_ ) );
OAI21_X1 _14725_ ( .A(_06030_ ), .B1(_04242_ ), .B2(_01655_ ), .ZN(_06639_ ) );
OAI21_X1 _14726_ ( .A(_06572_ ), .B1(_06638_ ), .B2(_06639_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
INV_X1 _14727_ ( .A(_05918_ ), .ZN(_06640_ ) );
OAI22_X1 _14728_ ( .A1(_04278_ ), .A2(_06118_ ), .B1(_01943_ ), .B2(_06383_ ), .ZN(_06641_ ) );
AOI21_X1 _14729_ ( .A(_04048_ ), .B1(_06496_ ), .B2(_02954_ ), .ZN(_06642_ ) );
XNOR2_X1 _14730_ ( .A(_06642_ ), .B(_02923_ ), .ZN(_06643_ ) );
AOI21_X1 _14731_ ( .A(_06641_ ), .B1(_06643_ ), .B2(_06501_ ), .ZN(_06644_ ) );
OAI21_X1 _14732_ ( .A(_04161_ ), .B1(_06644_ ), .B2(_06133_ ), .ZN(_06645_ ) );
BUF_X2 _14733_ ( .A(_06288_ ), .Z(_06646_ ) );
NAND4_X1 _14734_ ( .A1(_06646_ ), .A2(_06296_ ), .A3(_06301_ ), .A4(_06550_ ), .ZN(_06647_ ) );
AOI22_X1 _14735_ ( .A1(_06291_ ), .A2(_06294_ ), .B1(_06295_ ), .B2(_06647_ ), .ZN(_06648_ ) );
OR3_X1 _14736_ ( .A1(_06160_ ), .A2(_06163_ ), .A3(_03909_ ), .ZN(_06649_ ) );
NAND2_X1 _14737_ ( .A1(_06153_ ), .A2(_06297_ ), .ZN(_06650_ ) );
AOI21_X1 _14738_ ( .A(_06546_ ), .B1(_06649_ ), .B2(_06650_ ), .ZN(_06651_ ) );
NAND3_X1 _14739_ ( .A1(_06167_ ), .A2(_06171_ ), .A3(_06154_ ), .ZN(_06652_ ) );
OAI21_X1 _14740_ ( .A(_06352_ ), .B1(_06350_ ), .B2(_06356_ ), .ZN(_06653_ ) );
OAI21_X1 _14741_ ( .A(_06309_ ), .B1(_06347_ ), .B2(_06351_ ), .ZN(_06654_ ) );
NAND3_X1 _14742_ ( .A1(_06653_ ), .A2(_06654_ ), .A3(_06316_ ), .ZN(_06655_ ) );
AND3_X1 _14743_ ( .A1(_06652_ ), .A2(_06655_ ), .A3(_06175_ ), .ZN(_06656_ ) );
NOR3_X1 _14744_ ( .A1(_06651_ ), .A2(_06600_ ), .A3(_06656_ ), .ZN(_06657_ ) );
OAI21_X1 _14745_ ( .A(_06249_ ), .B1(_06648_ ), .B2(_06657_ ), .ZN(_06658_ ) );
CLKBUF_X2 _14746_ ( .A(_06634_ ), .Z(_06659_ ) );
AOI21_X1 _14747_ ( .A(_06556_ ), .B1(_06208_ ), .B2(_06227_ ), .ZN(_06660_ ) );
NOR2_X1 _14748_ ( .A1(_06660_ ), .A2(_06230_ ), .ZN(_06661_ ) );
AOI21_X1 _14749_ ( .A(_06659_ ), .B1(_06661_ ), .B2(_06555_ ), .ZN(_06662_ ) );
OAI21_X1 _14750_ ( .A(_06662_ ), .B1(_06555_ ), .B2(_06661_ ), .ZN(_06663_ ) );
NOR2_X1 _14751_ ( .A1(_06339_ ), .A2(_06343_ ), .ZN(_06664_ ) );
MUX2_X1 _14752_ ( .A(_06361_ ), .B(_06664_ ), .S(_06618_ ), .Z(_06665_ ) );
NAND2_X1 _14753_ ( .A1(_06665_ ), .A2(_06609_ ), .ZN(_06666_ ) );
BUF_X2 _14754_ ( .A(_06178_ ), .Z(_06667_ ) );
BUF_X4 _14755_ ( .A(_06546_ ), .Z(_06668_ ) );
BUF_X4 _14756_ ( .A(_06668_ ), .Z(_06669_ ) );
OAI21_X1 _14757_ ( .A(_06607_ ), .B1(_06311_ ), .B2(_06314_ ), .ZN(_06670_ ) );
OAI21_X1 _14758_ ( .A(_06620_ ), .B1(_06331_ ), .B2(_06335_ ), .ZN(_06671_ ) );
NAND2_X1 _14759_ ( .A1(_06670_ ), .A2(_06671_ ), .ZN(_06672_ ) );
OAI211_X1 _14760_ ( .A(_06666_ ), .B(_06667_ ), .C1(_06669_ ), .C2(_06672_ ), .ZN(_06673_ ) );
BUF_X4 _14761_ ( .A(_06620_ ), .Z(_06674_ ) );
NAND4_X1 _14762_ ( .A1(_06320_ ), .A2(_06600_ ), .A3(_06669_ ), .A4(_06674_ ), .ZN(_06675_ ) );
AOI21_X1 _14763_ ( .A(_06305_ ), .B1(_06673_ ), .B2(_06675_ ), .ZN(_06676_ ) );
AOI21_X1 _14764_ ( .A(_06565_ ), .B1(_03806_ ), .B2(_02922_ ), .ZN(_06677_ ) );
NOR2_X1 _14765_ ( .A1(_06651_ ), .A2(_06656_ ), .ZN(_06678_ ) );
AND3_X1 _14766_ ( .A1(_06678_ ), .A2(_06667_ ), .A3(_06181_ ), .ZN(_06679_ ) );
OR3_X1 _14767_ ( .A1(_03806_ ), .A2(_02922_ ), .A3(_06488_ ), .ZN(_06680_ ) );
OAI21_X1 _14768_ ( .A(_06680_ ), .B1(_06555_ ), .B2(_03987_ ), .ZN(_06681_ ) );
NOR4_X1 _14769_ ( .A1(_06676_ ), .A2(_06677_ ), .A3(_06679_ ), .A4(_06681_ ), .ZN(_06682_ ) );
NAND3_X1 _14770_ ( .A1(_06658_ ), .A2(_06663_ ), .A3(_06682_ ), .ZN(_06683_ ) );
AOI21_X1 _14771_ ( .A(_06645_ ), .B1(_06683_ ), .B2(_06377_ ), .ZN(_06684_ ) );
BUF_X2 _14772_ ( .A(_01649_ ), .Z(_06685_ ) );
NAND2_X1 _14773_ ( .A1(_04274_ ), .A2(_06685_ ), .ZN(_06686_ ) );
NAND2_X1 _14774_ ( .A1(_06686_ ), .A2(_05862_ ), .ZN(_06687_ ) );
OAI21_X1 _14775_ ( .A(_06640_ ), .B1(_06684_ ), .B2(_06687_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
INV_X1 _14776_ ( .A(_05925_ ), .ZN(_06688_ ) );
INV_X1 _14777_ ( .A(_06289_ ), .ZN(_06689_ ) );
INV_X1 _14778_ ( .A(_06646_ ), .ZN(_06690_ ) );
INV_X1 _14779_ ( .A(_06252_ ), .ZN(_06691_ ) );
AOI211_X1 _14780_ ( .A(_06689_ ), .B(_06690_ ), .C1(_06630_ ), .C2(_06691_ ), .ZN(_06692_ ) );
OR3_X1 _14781_ ( .A1(_06455_ ), .A2(_06458_ ), .A3(_06145_ ), .ZN(_06693_ ) );
OAI211_X1 _14782_ ( .A(_06452_ ), .B(_06145_ ), .C1(_01942_ ), .C2(_03921_ ), .ZN(_06694_ ) );
AND3_X1 _14783_ ( .A1(_06693_ ), .A2(_06694_ ), .A3(_03908_ ), .ZN(_06695_ ) );
AOI21_X1 _14784_ ( .A(_03908_ ), .B1(_06404_ ), .B2(_06407_ ), .ZN(_06696_ ) );
NOR2_X1 _14785_ ( .A1(_06695_ ), .A2(_06696_ ), .ZN(_06697_ ) );
AND2_X1 _14786_ ( .A1(_06411_ ), .A2(_06414_ ), .ZN(_06698_ ) );
MUX2_X1 _14787_ ( .A(_06698_ ), .B(_06421_ ), .S(_03909_ ), .Z(_06699_ ) );
MUX2_X1 _14788_ ( .A(_06697_ ), .B(_06699_ ), .S(_03911_ ), .Z(_06700_ ) );
AND2_X1 _14789_ ( .A1(_06700_ ), .A2(_06630_ ), .ZN(_06701_ ) );
OAI21_X1 _14790_ ( .A(_06249_ ), .B1(_06692_ ), .B2(_06701_ ), .ZN(_06702_ ) );
OAI21_X1 _14791_ ( .A(_06245_ ), .B1(_06554_ ), .B2(_06556_ ), .ZN(_06703_ ) );
AOI21_X1 _14792_ ( .A(_06703_ ), .B1(_06556_ ), .B2(_06554_ ), .ZN(_06704_ ) );
AND3_X1 _14793_ ( .A1(_06700_ ), .A2(_06667_ ), .A3(_06181_ ), .ZN(_06705_ ) );
AOI21_X1 _14794_ ( .A(_06565_ ), .B1(_03810_ ), .B2(_02953_ ), .ZN(_06706_ ) );
AND3_X1 _14795_ ( .A1(_06429_ ), .A2(_06172_ ), .A3(_06352_ ), .ZN(_06707_ ) );
BUF_X4 _14796_ ( .A(_06546_ ), .Z(_06708_ ) );
NAND2_X1 _14797_ ( .A1(_06707_ ), .A2(_06708_ ), .ZN(_06709_ ) );
AOI21_X1 _14798_ ( .A(_06305_ ), .B1(_06709_ ), .B2(_06443_ ), .ZN(_06710_ ) );
NAND3_X1 _14799_ ( .A1(_06448_ ), .A2(_06453_ ), .A3(_06317_ ), .ZN(_06711_ ) );
NAND3_X1 _14800_ ( .A1(_06464_ ), .A2(_06469_ ), .A3(_06325_ ), .ZN(_06712_ ) );
AOI21_X1 _14801_ ( .A(_06323_ ), .B1(_06711_ ), .B2(_06712_ ), .ZN(_06713_ ) );
NAND2_X1 _14802_ ( .A1(_06438_ ), .A2(_06618_ ), .ZN(_06714_ ) );
NAND2_X1 _14803_ ( .A1(_06473_ ), .A2(_06476_ ), .ZN(_06715_ ) );
NAND2_X1 _14804_ ( .A1(_06715_ ), .A2(_06620_ ), .ZN(_06716_ ) );
NAND2_X1 _14805_ ( .A1(_06714_ ), .A2(_06716_ ), .ZN(_06717_ ) );
AOI21_X1 _14806_ ( .A(_06713_ ), .B1(_06717_ ), .B2(_06364_ ), .ZN(_06718_ ) );
OAI21_X1 _14807_ ( .A(_06710_ ), .B1(_06718_ ), .B2(_06600_ ), .ZN(_06719_ ) );
NAND3_X1 _14808_ ( .A1(_03811_ ), .A2(_01965_ ), .A3(_06367_ ), .ZN(_06720_ ) );
OAI211_X1 _14809_ ( .A(_06719_ ), .B(_06720_ ), .C1(_06556_ ), .C2(_03987_ ), .ZN(_06721_ ) );
NOR4_X1 _14810_ ( .A1(_06704_ ), .A2(_06705_ ), .A3(_06706_ ), .A4(_06721_ ), .ZN(_06722_ ) );
AOI21_X1 _14811_ ( .A(_06375_ ), .B1(_06702_ ), .B2(_06722_ ), .ZN(_06723_ ) );
AOI21_X1 _14812_ ( .A(_06387_ ), .B1(_06496_ ), .B2(_02954_ ), .ZN(_06724_ ) );
OAI21_X1 _14813_ ( .A(_06724_ ), .B1(_02954_ ), .B2(_06496_ ), .ZN(_06725_ ) );
AOI22_X1 _14814_ ( .A1(_04298_ ), .A2(_06576_ ), .B1(\ID_EX_imm [16] ), .B2(_06577_ ), .ZN(_06726_ ) );
AOI21_X1 _14815_ ( .A(_06133_ ), .B1(_06725_ ), .B2(_06726_ ), .ZN(_06727_ ) );
NOR3_X1 _14816_ ( .A1(_06723_ ), .A2(_06685_ ), .A3(_06727_ ), .ZN(_06728_ ) );
BUF_X4 _14817_ ( .A(_01654_ ), .Z(_06729_ ) );
OAI21_X1 _14818_ ( .A(_06030_ ), .B1(_04296_ ), .B2(_06729_ ), .ZN(_06730_ ) );
OAI21_X1 _14819_ ( .A(_06688_ ), .B1(_06728_ ), .B2(_06730_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
NAND2_X1 _14820_ ( .A1(_04003_ ), .A2(_03319_ ), .ZN(_06731_ ) );
AND2_X1 _14821_ ( .A1(_06731_ ), .A2(_04022_ ), .ZN(_06732_ ) );
INV_X1 _14822_ ( .A(_03189_ ), .ZN(_06733_ ) );
NOR2_X1 _14823_ ( .A1(_06732_ ), .A2(_06733_ ), .ZN(_06734_ ) );
NOR2_X1 _14824_ ( .A1(_06734_ ), .A2(_04010_ ), .ZN(_06735_ ) );
INV_X1 _14825_ ( .A(_06735_ ), .ZN(_06736_ ) );
AOI21_X1 _14826_ ( .A(_04011_ ), .B1(_06736_ ), .B2(_04009_ ), .ZN(_06737_ ) );
NOR2_X1 _14827_ ( .A1(_06737_ ), .A2(_03137_ ), .ZN(_06738_ ) );
INV_X1 _14828_ ( .A(_06738_ ), .ZN(_06739_ ) );
AND3_X1 _14829_ ( .A1(_06739_ ), .A2(_03163_ ), .A3(_04006_ ), .ZN(_06740_ ) );
AOI21_X1 _14830_ ( .A(_03163_ ), .B1(_06739_ ), .B2(_04006_ ), .ZN(_06741_ ) );
NOR3_X1 _14831_ ( .A1(_06740_ ), .A2(_06741_ ), .A3(_06387_ ), .ZN(_06742_ ) );
OAI22_X1 _14832_ ( .A1(_04323_ ), .A2(_06118_ ), .B1(_02310_ ), .B2(_06383_ ), .ZN(_06743_ ) );
OAI21_X1 _14833_ ( .A(_06381_ ), .B1(_06742_ ), .B2(_06743_ ), .ZN(_06744_ ) );
NAND2_X1 _14834_ ( .A1(_06744_ ), .A2(_06391_ ), .ZN(_06745_ ) );
INV_X1 _14835_ ( .A(_03850_ ), .ZN(_06746_ ) );
AND2_X1 _14836_ ( .A1(_06204_ ), .A2(_06207_ ), .ZN(_06747_ ) );
INV_X1 _14837_ ( .A(_06747_ ), .ZN(_06748_ ) );
AOI211_X1 _14838_ ( .A(_06746_ ), .B(_03845_ ), .C1(_06748_ ), .C2(_06217_ ), .ZN(_06749_ ) );
INV_X1 _14839_ ( .A(_06749_ ), .ZN(_06750_ ) );
AOI21_X1 _14840_ ( .A(_03840_ ), .B1(_06750_ ), .B2(_06223_ ), .ZN(_06751_ ) );
OR3_X1 _14841_ ( .A1(_06751_ ), .A2(_03834_ ), .A3(_06225_ ), .ZN(_06752_ ) );
OAI21_X1 _14842_ ( .A(_03834_ ), .B1(_06751_ ), .B2(_06225_ ), .ZN(_06753_ ) );
NAND3_X1 _14843_ ( .A1(_06752_ ), .A2(_06561_ ), .A3(_06753_ ), .ZN(_06754_ ) );
NAND4_X1 _14844_ ( .A1(_06646_ ), .A2(_06248_ ), .A3(_06292_ ), .A4(_06289_ ), .ZN(_06755_ ) );
OAI21_X1 _14845_ ( .A(_06297_ ), .B1(_06542_ ), .B2(_06543_ ), .ZN(_06756_ ) );
OAI21_X1 _14846_ ( .A(_06422_ ), .B1(_06532_ ), .B2(_06533_ ), .ZN(_06757_ ) );
NAND2_X1 _14847_ ( .A1(_06756_ ), .A2(_06757_ ), .ZN(_06758_ ) );
NAND2_X1 _14848_ ( .A1(_06758_ ), .A2(_06364_ ), .ZN(_06759_ ) );
OAI21_X1 _14849_ ( .A(_06618_ ), .B1(_06535_ ), .B2(_06536_ ), .ZN(_06760_ ) );
NOR3_X1 _14850_ ( .A1(_06355_ ), .A2(_06329_ ), .A3(_06359_ ), .ZN(_06761_ ) );
NOR3_X1 _14851_ ( .A1(_06350_ ), .A2(_06356_ ), .A3(_06342_ ), .ZN(_06762_ ) );
OAI21_X1 _14852_ ( .A(_06317_ ), .B1(_06761_ ), .B2(_06762_ ), .ZN(_06763_ ) );
AND2_X1 _14853_ ( .A1(_06760_ ), .A2(_06763_ ), .ZN(_06764_ ) );
BUF_X2 _14854_ ( .A(_06323_ ), .Z(_06765_ ) );
OAI211_X1 _14855_ ( .A(_06759_ ), .B(_06425_ ), .C1(_06764_ ), .C2(_06765_ ), .ZN(_06766_ ) );
OR2_X1 _14856_ ( .A1(_06180_ ), .A2(_06247_ ), .ZN(_06767_ ) );
AND3_X1 _14857_ ( .A1(_06152_ ), .A2(_06172_ ), .A3(_06352_ ), .ZN(_06768_ ) );
AND2_X1 _14858_ ( .A1(_06768_ ), .A2(_06175_ ), .ZN(_06769_ ) );
OAI211_X1 _14859_ ( .A(_06766_ ), .B(_06767_ ), .C1(_06667_ ), .C2(_06769_ ), .ZN(_06770_ ) );
NOR2_X1 _14860_ ( .A1(_06515_ ), .A2(_06297_ ), .ZN(_06771_ ) );
AOI21_X1 _14861_ ( .A(_06316_ ), .B1(_06507_ ), .B2(_06508_ ), .ZN(_06772_ ) );
OR3_X1 _14862_ ( .A1(_06771_ ), .A2(_06772_ ), .A3(_06546_ ), .ZN(_06773_ ) );
OAI21_X1 _14863_ ( .A(_06618_ ), .B1(_06517_ ), .B2(_06518_ ), .ZN(_06774_ ) );
OAI21_X1 _14864_ ( .A(_06317_ ), .B1(_06525_ ), .B2(_06526_ ), .ZN(_06775_ ) );
NAND3_X1 _14865_ ( .A1(_06774_ ), .A2(_06775_ ), .A3(_06708_ ), .ZN(_06776_ ) );
AND2_X2 _14866_ ( .A1(_06177_ ), .A2(_04070_ ), .ZN(_06777_ ) );
BUF_X2 _14867_ ( .A(_06777_ ), .Z(_06778_ ) );
NAND3_X1 _14868_ ( .A1(_06773_ ), .A2(_06776_ ), .A3(_06778_ ), .ZN(_06779_ ) );
NAND2_X1 _14869_ ( .A1(_03834_ ), .A2(_06368_ ), .ZN(_06780_ ) );
AOI21_X1 _14870_ ( .A(_06135_ ), .B1(_03833_ ), .B2(_03954_ ), .ZN(_06781_ ) );
AOI21_X1 _14871_ ( .A(_06781_ ), .B1(_06220_ ), .B2(_06367_ ), .ZN(_06782_ ) );
AND2_X1 _14872_ ( .A1(_06780_ ), .A2(_06782_ ), .ZN(_06783_ ) );
AND4_X1 _14873_ ( .A1(_06755_ ), .A2(_06770_ ), .A3(_06779_ ), .A4(_06783_ ), .ZN(_06784_ ) );
AOI21_X1 _14874_ ( .A(_06375_ ), .B1(_06754_ ), .B2(_06784_ ), .ZN(_06785_ ) );
OAI221_X1 _14875_ ( .A(_05888_ ), .B1(_06391_ ), .B2(_04317_ ), .C1(_06745_ ), .C2(_06785_ ), .ZN(_06786_ ) );
INV_X1 _14876_ ( .A(_05930_ ), .ZN(_06787_ ) );
NAND2_X1 _14877_ ( .A1(_06786_ ), .A2(_06787_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
AND2_X1 _14878_ ( .A1(_06646_ ), .A2(_06301_ ), .ZN(_06788_ ) );
AND2_X2 _14879_ ( .A1(_06289_ ), .A2(_06292_ ), .ZN(_06789_ ) );
AND2_X1 _14880_ ( .A1(_06788_ ), .A2(_06789_ ), .ZN(_06790_ ) );
INV_X1 _14881_ ( .A(_06790_ ), .ZN(_06791_ ) );
NAND3_X1 _14882_ ( .A1(_06396_ ), .A2(_06422_ ), .A3(_06334_ ), .ZN(_06792_ ) );
AND3_X1 _14883_ ( .A1(_06278_ ), .A2(_06287_ ), .A3(_06792_ ), .ZN(_06793_ ) );
BUF_X4 _14884_ ( .A(_06789_ ), .Z(_06794_ ) );
OAI21_X1 _14885_ ( .A(_06297_ ), .B1(_06595_ ), .B2(_06596_ ), .ZN(_06795_ ) );
OAI21_X1 _14886_ ( .A(_06422_ ), .B1(_06587_ ), .B2(_06588_ ), .ZN(_06796_ ) );
NAND2_X1 _14887_ ( .A1(_06795_ ), .A2(_06796_ ), .ZN(_06797_ ) );
NAND2_X1 _14888_ ( .A1(_06797_ ), .A2(_06364_ ), .ZN(_06798_ ) );
NOR3_X1 _14889_ ( .A1(_06449_ ), .A2(_06395_ ), .A3(_06446_ ), .ZN(_06799_ ) );
NOR3_X1 _14890_ ( .A1(_06457_ ), .A2(_06451_ ), .A3(_06334_ ), .ZN(_06800_ ) );
OAI21_X1 _14891_ ( .A(_06620_ ), .B1(_06799_ ), .B2(_06800_ ), .ZN(_06801_ ) );
NAND3_X1 _14892_ ( .A1(_06590_ ), .A2(_06591_ ), .A3(_06325_ ), .ZN(_06802_ ) );
AND2_X1 _14893_ ( .A1(_06801_ ), .A2(_06802_ ), .ZN(_06803_ ) );
OAI211_X1 _14894_ ( .A(_06798_ ), .B(_06425_ ), .C1(_06765_ ), .C2(_06803_ ), .ZN(_06804_ ) );
AND3_X1 _14895_ ( .A1(_06420_ ), .A2(_06172_ ), .A3(_06151_ ), .ZN(_06805_ ) );
AND2_X1 _14896_ ( .A1(_06805_ ), .A2(_06175_ ), .ZN(_06806_ ) );
OR2_X1 _14897_ ( .A1(_06806_ ), .A2(_06178_ ), .ZN(_06807_ ) );
AOI22_X1 _14898_ ( .A1(_06793_ ), .A2(_06794_ ), .B1(_06804_ ), .B2(_06807_ ), .ZN(_06808_ ) );
AOI21_X1 _14899_ ( .A(_06394_ ), .B1(_06791_ ), .B2(_06808_ ), .ZN(_06809_ ) );
NOR2_X1 _14900_ ( .A1(_06625_ ), .A2(_06626_ ), .ZN(_06810_ ) );
MUX2_X1 _14901_ ( .A(_06606_ ), .B(_06810_ ), .S(_06172_ ), .Z(_06811_ ) );
NAND2_X1 _14902_ ( .A1(_06811_ ), .A2(_03911_ ), .ZN(_06812_ ) );
OAI21_X1 _14903_ ( .A(_06154_ ), .B1(_06622_ ), .B2(_06623_ ), .ZN(_06813_ ) );
NAND3_X1 _14904_ ( .A1(_06615_ ), .A2(_06616_ ), .A3(_06316_ ), .ZN(_06814_ ) );
NAND3_X1 _14905_ ( .A1(_06813_ ), .A2(_06175_ ), .A3(_06814_ ), .ZN(_06815_ ) );
AND3_X1 _14906_ ( .A1(_06812_ ), .A2(_06777_ ), .A3(_06815_ ), .ZN(_06816_ ) );
AOI221_X4 _14907_ ( .A(_06816_ ), .B1(_06225_ ), .B2(_06367_ ), .C1(_03839_ ), .C2(_03986_ ), .ZN(_06817_ ) );
BUF_X2 _14908_ ( .A(_06181_ ), .Z(_06818_ ) );
NAND3_X1 _14909_ ( .A1(_06807_ ), .A2(_06818_ ), .A3(_06804_ ), .ZN(_06819_ ) );
OAI21_X1 _14910_ ( .A(_06486_ ), .B1(_03936_ ), .B2(_02332_ ), .ZN(_06820_ ) );
NAND3_X1 _14911_ ( .A1(_06817_ ), .A2(_06819_ ), .A3(_06820_ ), .ZN(_06821_ ) );
NOR2_X1 _14912_ ( .A1(_06809_ ), .A2(_06821_ ), .ZN(_06822_ ) );
AND3_X1 _14913_ ( .A1(_06750_ ), .A2(_03840_ ), .A3(_06223_ ), .ZN(_06823_ ) );
OR3_X1 _14914_ ( .A1(_06823_ ), .A2(_06751_ ), .A3(_06659_ ), .ZN(_06824_ ) );
AOI21_X1 _14915_ ( .A(_06375_ ), .B1(_06822_ ), .B2(_06824_ ), .ZN(_06825_ ) );
NAND2_X1 _14916_ ( .A1(_06737_ ), .A2(_03137_ ), .ZN(_06826_ ) );
NAND3_X1 _14917_ ( .A1(_06739_ ), .A2(_06501_ ), .A3(_06826_ ), .ZN(_06827_ ) );
AOI22_X1 _14918_ ( .A1(_04351_ ), .A2(_06576_ ), .B1(\ID_EX_imm [14] ), .B2(_06577_ ), .ZN(_06828_ ) );
AOI21_X1 _14919_ ( .A(_06573_ ), .B1(_06827_ ), .B2(_06828_ ), .ZN(_06829_ ) );
OR2_X1 _14920_ ( .A1(_06829_ ), .A2(_06685_ ), .ZN(_06830_ ) );
OAI221_X1 _14921_ ( .A(_05888_ ), .B1(_06391_ ), .B2(_04348_ ), .C1(_06825_ ), .C2(_06830_ ), .ZN(_06831_ ) );
INV_X1 _14922_ ( .A(_05935_ ), .ZN(_06832_ ) );
NAND2_X1 _14923_ ( .A1(_06831_ ), .A2(_06832_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
OR3_X1 _14924_ ( .A1(_04367_ ), .A2(_05861_ ), .A3(_04369_ ), .ZN(_06833_ ) );
AOI21_X1 _14925_ ( .A(_06386_ ), .B1(_06736_ ), .B2(_03215_ ), .ZN(_06834_ ) );
OAI21_X1 _14926_ ( .A(_06834_ ), .B1(_03215_ ), .B2(_06736_ ), .ZN(_06835_ ) );
OR2_X1 _14927_ ( .A1(_04380_ ), .A2(_06117_ ), .ZN(_06836_ ) );
NAND3_X1 _14928_ ( .A1(_06127_ ), .A2(\ID_EX_imm [13] ), .A3(_06128_ ), .ZN(_06837_ ) );
AND3_X1 _14929_ ( .A1(_06835_ ), .A2(_06836_ ), .A3(_06837_ ), .ZN(_06838_ ) );
OAI21_X1 _14930_ ( .A(_01654_ ), .B1(_06838_ ), .B2(_06133_ ), .ZN(_06839_ ) );
OAI211_X1 _14931_ ( .A(_06646_ ), .B(_06794_ ), .C1(_06298_ ), .C2(_06301_ ), .ZN(_06840_ ) );
NAND2_X1 _14932_ ( .A1(_06174_ ), .A2(_06765_ ), .ZN(_06841_ ) );
BUF_X2 _14933_ ( .A(_06364_ ), .Z(_06842_ ) );
NAND3_X1 _14934_ ( .A1(_06653_ ), .A2(_06654_ ), .A3(_06297_ ), .ZN(_06843_ ) );
OAI21_X1 _14935_ ( .A(_06342_ ), .B1(_06358_ ), .B2(_06338_ ), .ZN(_06844_ ) );
OAI21_X1 _14936_ ( .A(_06329_ ), .B1(_06355_ ), .B2(_06359_ ), .ZN(_06845_ ) );
NAND3_X1 _14937_ ( .A1(_06844_ ), .A2(_06845_ ), .A3(_06422_ ), .ZN(_06846_ ) );
AND2_X1 _14938_ ( .A1(_06843_ ), .A2(_06846_ ), .ZN(_06847_ ) );
OAI211_X1 _14939_ ( .A(_06841_ ), .B(_06530_ ), .C1(_06842_ ), .C2(_06847_ ), .ZN(_06848_ ) );
NOR3_X1 _14940_ ( .A1(_06153_ ), .A2(_06323_ ), .A3(_06618_ ), .ZN(_06849_ ) );
OR2_X1 _14941_ ( .A1(_06849_ ), .A2(_06425_ ), .ZN(_06850_ ) );
NAND2_X1 _14942_ ( .A1(_06848_ ), .A2(_06850_ ), .ZN(_06851_ ) );
AOI21_X1 _14943_ ( .A(_06394_ ), .B1(_06840_ ), .B2(_06851_ ), .ZN(_06852_ ) );
AND3_X1 _14944_ ( .A1(_06848_ ), .A2(_06818_ ), .A3(_06850_ ), .ZN(_06853_ ) );
NAND2_X1 _14945_ ( .A1(_06321_ ), .A2(_06364_ ), .ZN(_06854_ ) );
NAND3_X1 _14946_ ( .A1(_06336_ ), .A2(_06344_ ), .A3(_06708_ ), .ZN(_06855_ ) );
AND3_X1 _14947_ ( .A1(_06854_ ), .A2(_06855_ ), .A3(_06778_ ), .ZN(_06856_ ) );
NOR3_X1 _14948_ ( .A1(_06852_ ), .A2(_06853_ ), .A3(_06856_ ), .ZN(_06857_ ) );
AOI21_X1 _14949_ ( .A(_03845_ ), .B1(_06748_ ), .B2(_06217_ ), .ZN(_06858_ ) );
OR3_X1 _14950_ ( .A1(_06858_ ), .A2(_03850_ ), .A3(_06222_ ), .ZN(_06859_ ) );
OAI21_X1 _14951_ ( .A(_03850_ ), .B1(_06858_ ), .B2(_06222_ ), .ZN(_06860_ ) );
NAND3_X1 _14952_ ( .A1(_06859_ ), .A2(_06561_ ), .A3(_06860_ ), .ZN(_06861_ ) );
AND2_X1 _14953_ ( .A1(_03850_ ), .A2(_06567_ ), .ZN(_06862_ ) );
NOR3_X1 _14954_ ( .A1(_03849_ ), .A2(_03214_ ), .A3(_06488_ ), .ZN(_06863_ ) );
AOI21_X1 _14955_ ( .A(_06565_ ), .B1(_03849_ ), .B2(_03214_ ), .ZN(_06864_ ) );
NOR3_X1 _14956_ ( .A1(_06862_ ), .A2(_06863_ ), .A3(_06864_ ), .ZN(_06865_ ) );
NAND3_X1 _14957_ ( .A1(_06857_ ), .A2(_06861_ ), .A3(_06865_ ), .ZN(_06866_ ) );
AOI21_X1 _14958_ ( .A(_06839_ ), .B1(_06866_ ), .B2(_06377_ ), .ZN(_06867_ ) );
OAI21_X1 _14959_ ( .A(_06030_ ), .B1(_04375_ ), .B2(_06729_ ), .ZN(_06868_ ) );
OAI21_X1 _14960_ ( .A(_06833_ ), .B1(_06867_ ), .B2(_06868_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
INV_X1 _14961_ ( .A(_05948_ ), .ZN(_06869_ ) );
AND3_X1 _14962_ ( .A1(_06731_ ), .A2(_06733_ ), .A3(_04022_ ), .ZN(_06870_ ) );
OR3_X1 _14963_ ( .A1(_06734_ ), .A2(_06386_ ), .A3(_06870_ ), .ZN(_06871_ ) );
AOI22_X1 _14964_ ( .A1(_04421_ ), .A2(_06576_ ), .B1(\ID_EX_imm [12] ), .B2(_06577_ ), .ZN(_06872_ ) );
AOI21_X1 _14965_ ( .A(_06573_ ), .B1(_06871_ ), .B2(_06872_ ), .ZN(_06873_ ) );
OR2_X1 _14966_ ( .A1(_06873_ ), .A2(_01650_ ), .ZN(_06874_ ) );
OAI211_X1 _14967_ ( .A(_06646_ ), .B(_06794_ ), .C1(_06301_ ), .C2(_06397_ ), .ZN(_06875_ ) );
OR2_X1 _14968_ ( .A1(_06875_ ), .A2(_06394_ ), .ZN(_06876_ ) );
AND3_X1 _14969_ ( .A1(_06748_ ), .A2(_03845_ ), .A3(_06217_ ), .ZN(_06877_ ) );
OR3_X1 _14970_ ( .A1(_06877_ ), .A2(_06858_ ), .A3(_06659_ ), .ZN(_06878_ ) );
OAI21_X1 _14971_ ( .A(_06150_ ), .B1(_06444_ ), .B2(_06467_ ), .ZN(_06879_ ) );
OAI21_X1 _14972_ ( .A(_06157_ ), .B1(_06449_ ), .B2(_06446_ ), .ZN(_06880_ ) );
NAND2_X1 _14973_ ( .A1(_06879_ ), .A2(_06880_ ), .ZN(_06881_ ) );
AND2_X1 _14974_ ( .A1(_06693_ ), .A2(_06694_ ), .ZN(_06882_ ) );
MUX2_X1 _14975_ ( .A(_06881_ ), .B(_06882_ ), .S(_06618_ ), .Z(_06883_ ) );
NAND2_X1 _14976_ ( .A1(_06883_ ), .A2(_06609_ ), .ZN(_06884_ ) );
OAI211_X1 _14977_ ( .A(_06884_ ), .B(_06667_ ), .C1(_06669_ ), .C2(_06416_ ), .ZN(_06885_ ) );
NAND4_X1 _14978_ ( .A1(_06421_ ), .A2(_06600_ ), .A3(_06669_ ), .A4(_06674_ ), .ZN(_06886_ ) );
INV_X1 _14979_ ( .A(_06180_ ), .ZN(_06887_ ) );
AOI22_X1 _14980_ ( .A1(_06885_ ), .A2(_06886_ ), .B1(_06394_ ), .B2(_06887_ ), .ZN(_06888_ ) );
NOR2_X1 _14981_ ( .A1(_06439_ ), .A2(_06708_ ), .ZN(_06889_ ) );
NOR3_X1 _14982_ ( .A1(_06470_ ), .A2(_06323_ ), .A3(_06477_ ), .ZN(_06890_ ) );
OAI21_X1 _14983_ ( .A(_06667_ ), .B1(_06889_ ), .B2(_06890_ ), .ZN(_06891_ ) );
NOR2_X1 _14984_ ( .A1(_06891_ ), .A2(_06305_ ), .ZN(_06892_ ) );
NOR3_X1 _14985_ ( .A1(_03843_ ), .A2(_03188_ ), .A3(_06488_ ), .ZN(_06893_ ) );
OAI21_X1 _14986_ ( .A(_04075_ ), .B1(_03950_ ), .B2(_02380_ ), .ZN(_06894_ ) );
OAI21_X1 _14987_ ( .A(_06894_ ), .B1(_03845_ ), .B2(_03987_ ), .ZN(_06895_ ) );
NOR4_X1 _14988_ ( .A1(_06888_ ), .A2(_06892_ ), .A3(_06893_ ), .A4(_06895_ ), .ZN(_06896_ ) );
NAND3_X1 _14989_ ( .A1(_06876_ ), .A2(_06878_ ), .A3(_06896_ ), .ZN(_06897_ ) );
AOI21_X1 _14990_ ( .A(_06874_ ), .B1(_06897_ ), .B2(_06377_ ), .ZN(_06898_ ) );
OAI21_X1 _14991_ ( .A(_06030_ ), .B1(_04419_ ), .B2(_06729_ ), .ZN(_06899_ ) );
OAI21_X1 _14992_ ( .A(_06869_ ), .B1(_06898_ ), .B2(_06899_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
OR2_X1 _14993_ ( .A1(_02719_ ), .A2(_05891_ ), .ZN(_06900_ ) );
OR2_X1 _14994_ ( .A1(_02858_ ), .A2(_01654_ ), .ZN(_06901_ ) );
AOI22_X1 _14995_ ( .A1(_02830_ ), .A2(_06576_ ), .B1(\ID_EX_imm [30] ), .B2(_06577_ ), .ZN(_06902_ ) );
AOI211_X1 _14996_ ( .A(_03110_ ), .B(_03008_ ), .C1(_04004_ ), .C2(_04024_ ), .ZN(_06903_ ) );
OAI21_X1 _14997_ ( .A(_03527_ ), .B1(_06903_ ), .B2(_04067_ ), .ZN(_06904_ ) );
AND2_X1 _14998_ ( .A1(_06904_ ), .A2(_04039_ ), .ZN(_06905_ ) );
AOI21_X1 _14999_ ( .A(_03738_ ), .B1(_03593_ ), .B2(_03574_ ), .ZN(_06906_ ) );
INV_X1 _15000_ ( .A(_03617_ ), .ZN(_06907_ ) );
NOR4_X1 _15001_ ( .A1(_06905_ ), .A2(_06906_ ), .A3(_04043_ ), .A4(_06907_ ), .ZN(_06908_ ) );
OR2_X1 _15002_ ( .A1(_06908_ ), .A2(_04047_ ), .ZN(_06909_ ) );
AOI21_X1 _15003_ ( .A(_06387_ ), .B1(_06909_ ), .B2(_03550_ ), .ZN(_06910_ ) );
OAI21_X1 _15004_ ( .A(_06910_ ), .B1(_03550_ ), .B2(_06909_ ), .ZN(_06911_ ) );
AOI21_X1 _15005_ ( .A(_06573_ ), .B1(_06902_ ), .B2(_06911_ ), .ZN(_06912_ ) );
OR2_X1 _15006_ ( .A1(_06912_ ), .A2(_06685_ ), .ZN(_06913_ ) );
NAND3_X1 _15007_ ( .A1(_06806_ ), .A2(_06177_ ), .A3(_06180_ ), .ZN(_06914_ ) );
NAND3_X1 _15008_ ( .A1(_06137_ ), .A2(_03978_ ), .A3(_03723_ ), .ZN(_06915_ ) );
INV_X1 _15009_ ( .A(_03745_ ), .ZN(_06916_ ) );
OAI211_X1 _15010_ ( .A(_06914_ ), .B(_06915_ ), .C1(_06916_ ), .C2(_03987_ ), .ZN(_06917_ ) );
NOR2_X1 _15011_ ( .A1(_06177_ ), .A2(_06305_ ), .ZN(_06918_ ) );
AND3_X1 _15012_ ( .A1(_06812_ ), .A2(_06815_ ), .A3(_06918_ ), .ZN(_06919_ ) );
NOR2_X1 _15013_ ( .A1(_03743_ ), .A2(_06135_ ), .ZN(_06920_ ) );
OR3_X1 _15014_ ( .A1(_06917_ ), .A2(_06919_ ), .A3(_06920_ ), .ZN(_06921_ ) );
OR3_X1 _15015_ ( .A1(_06402_ ), .A2(_06309_ ), .A3(_06406_ ), .ZN(_06922_ ) );
OR3_X1 _15016_ ( .A1(_06455_ ), .A2(_06403_ ), .A3(_06151_ ), .ZN(_06923_ ) );
NAND2_X1 _15017_ ( .A1(_06922_ ), .A2(_06923_ ), .ZN(_06924_ ) );
NAND2_X1 _15018_ ( .A1(_06924_ ), .A2(_06317_ ), .ZN(_06925_ ) );
NAND3_X1 _15019_ ( .A1(_06612_ ), .A2(_06613_ ), .A3(_06325_ ), .ZN(_06926_ ) );
NAND2_X1 _15020_ ( .A1(_06925_ ), .A2(_06926_ ), .ZN(_06927_ ) );
NOR2_X1 _15021_ ( .A1(_06409_ ), .A2(_06413_ ), .ZN(_06928_ ) );
NAND2_X1 _15022_ ( .A1(_06928_ ), .A2(_06342_ ), .ZN(_06929_ ) );
OR3_X1 _15023_ ( .A1(_06405_ ), .A2(_06410_ ), .A3(_06146_ ), .ZN(_06930_ ) );
NAND2_X1 _15024_ ( .A1(_06929_ ), .A2(_06930_ ), .ZN(_06931_ ) );
NOR2_X1 _15025_ ( .A1(_06412_ ), .A2(_06418_ ), .ZN(_06932_ ) );
AOI21_X1 _15026_ ( .A(_06417_ ), .B1(_01732_ ), .B2(_06147_ ), .ZN(_06933_ ) );
MUX2_X1 _15027_ ( .A(_06932_ ), .B(_06933_ ), .S(_06352_ ), .Z(_06934_ ) );
MUX2_X1 _15028_ ( .A(_06931_ ), .B(_06934_ ), .S(_06349_ ), .Z(_06935_ ) );
MUX2_X1 _15029_ ( .A(_06927_ ), .B(_06935_ ), .S(_06708_ ), .Z(_06936_ ) );
OAI211_X1 _15030_ ( .A(_06288_ ), .B(_06792_ ), .C1(_06289_ ), .C2(_06293_ ), .ZN(_06937_ ) );
INV_X1 _15031_ ( .A(_06937_ ), .ZN(_06938_ ) );
AND2_X1 _15032_ ( .A1(_06806_ ), .A2(_06177_ ), .ZN(_06939_ ) );
AND4_X1 _15033_ ( .A1(_06300_ ), .A2(_06278_ ), .A3(_06287_ ), .A4(_06293_ ), .ZN(_06940_ ) );
OR4_X1 _15034_ ( .A1(_06549_ ), .A2(_06938_ ), .A3(_06939_ ), .A4(_06940_ ), .ZN(_06941_ ) );
AOI221_X2 _15035_ ( .A(_06921_ ), .B1(_06777_ ), .B2(_06936_ ), .C1(_06941_ ), .C2(_06247_ ), .ZN(_06942_ ) );
NOR3_X1 _15036_ ( .A1(_03788_ ), .A2(_03784_ ), .A3(_03789_ ), .ZN(_06943_ ) );
AND3_X1 _15037_ ( .A1(_06943_ ), .A2(_03794_ ), .A3(_03798_ ), .ZN(_06944_ ) );
INV_X1 _15038_ ( .A(_06944_ ), .ZN(_06945_ ) );
AOI211_X1 _15039_ ( .A(_06185_ ), .B(_06945_ ), .C1(_06208_ ), .C2(_06227_ ), .ZN(_06946_ ) );
NOR2_X1 _15040_ ( .A1(_06237_ ), .A2(_06945_ ), .ZN(_06947_ ) );
NOR4_X1 _15041_ ( .A1(_03826_ ), .A2(_03793_ ), .A3(_03827_ ), .A4(_03084_ ), .ZN(_06948_ ) );
OR2_X1 _15042_ ( .A1(_06948_ ), .A2(_03827_ ), .ZN(_06949_ ) );
AND2_X1 _15043_ ( .A1(_06949_ ), .A2(_06943_ ), .ZN(_06950_ ) );
NOR4_X1 _15044_ ( .A1(_03788_ ), .A2(_03033_ ), .A3(_03789_ ), .A4(_03782_ ), .ZN(_06951_ ) );
NOR4_X1 _15045_ ( .A1(_06947_ ), .A2(_03788_ ), .A3(_06950_ ), .A4(_06951_ ), .ZN(_06952_ ) );
INV_X1 _15046_ ( .A(_06952_ ), .ZN(_06953_ ) );
OAI211_X1 _15047_ ( .A(_03772_ ), .B(_03778_ ), .C1(_06946_ ), .C2(_06953_ ), .ZN(_06954_ ) );
NOR2_X1 _15048_ ( .A1(_03771_ ), .A2(_06168_ ), .ZN(_06955_ ) );
AOI21_X1 _15049_ ( .A(_03776_ ), .B1(_03778_ ), .B2(_06955_ ), .ZN(_06956_ ) );
AOI211_X2 _15050_ ( .A(_03767_ ), .B(_03759_ ), .C1(_06954_ ), .C2(_06956_ ), .ZN(_06957_ ) );
INV_X1 _15051_ ( .A(_03765_ ), .ZN(_06958_ ) );
AOI21_X1 _15052_ ( .A(_03764_ ), .B1(_06958_ ), .B2(_03756_ ), .ZN(_06959_ ) );
INV_X1 _15053_ ( .A(_06959_ ), .ZN(_06960_ ) );
OAI211_X1 _15054_ ( .A(_03739_ ), .B(_03733_ ), .C1(_06957_ ), .C2(_06960_ ), .ZN(_06961_ ) );
AND3_X1 _15055_ ( .A1(_03739_ ), .A2(_01765_ ), .A3(_03731_ ), .ZN(_06962_ ) );
AOI21_X1 _15056_ ( .A(_06962_ ), .B1(_02539_ ), .B2(_03737_ ), .ZN(_06963_ ) );
AND3_X1 _15057_ ( .A1(_06961_ ), .A2(_06916_ ), .A3(_06963_ ), .ZN(_06964_ ) );
AOI21_X1 _15058_ ( .A(_06916_ ), .B1(_06961_ ), .B2(_06963_ ), .ZN(_06965_ ) );
OR3_X1 _15059_ ( .A1(_06964_ ), .A2(_06965_ ), .A3(_06659_ ), .ZN(_06966_ ) );
AOI21_X1 _15060_ ( .A(_06375_ ), .B1(_06942_ ), .B2(_06966_ ), .ZN(_06967_ ) );
OAI21_X1 _15061_ ( .A(_06901_ ), .B1(_06913_ ), .B2(_06967_ ), .ZN(_06968_ ) );
OAI21_X1 _15062_ ( .A(_06900_ ), .B1(_06968_ ), .B2(_05865_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _15063_ ( .A1(_04436_ ), .A2(_05879_ ), .A3(_04438_ ), .ZN(_06969_ ) );
NAND4_X1 _15064_ ( .A1(_06278_ ), .A2(_06287_ ), .A3(_06550_ ), .A4(_06794_ ), .ZN(_06970_ ) );
OAI21_X1 _15065_ ( .A(_06600_ ), .B1(_06545_ ), .B2(_06765_ ), .ZN(_06971_ ) );
OAI21_X1 _15066_ ( .A(_06325_ ), .B1(_06761_ ), .B2(_06762_ ), .ZN(_06972_ ) );
NOR3_X1 _15067_ ( .A1(_06337_ ), .A2(_06329_ ), .A3(_06341_ ), .ZN(_06973_ ) );
NOR3_X1 _15068_ ( .A1(_06358_ ), .A2(_06338_ ), .A3(_06342_ ), .ZN(_06974_ ) );
OAI21_X1 _15069_ ( .A(_06349_ ), .B1(_06973_ ), .B2(_06974_ ), .ZN(_06975_ ) );
NAND2_X1 _15070_ ( .A1(_06972_ ), .A2(_06975_ ), .ZN(_06976_ ) );
NAND2_X1 _15071_ ( .A1(_06976_ ), .A2(_06609_ ), .ZN(_06977_ ) );
NAND2_X1 _15072_ ( .A1(_06538_ ), .A2(_06765_ ), .ZN(_06978_ ) );
NAND3_X1 _15073_ ( .A1(_06977_ ), .A2(_06978_ ), .A3(_06530_ ), .ZN(_06979_ ) );
NAND2_X1 _15074_ ( .A1(_06971_ ), .A2(_06979_ ), .ZN(_06980_ ) );
INV_X1 _15075_ ( .A(_06788_ ), .ZN(_06981_ ) );
INV_X1 _15076_ ( .A(_06794_ ), .ZN(_06982_ ) );
OAI211_X1 _15077_ ( .A(_06970_ ), .B(_06980_ ), .C1(_06981_ ), .C2(_06982_ ), .ZN(_06983_ ) );
NAND2_X1 _15078_ ( .A1(_06983_ ), .A2(_06249_ ), .ZN(_06984_ ) );
INV_X1 _15079_ ( .A(_03855_ ), .ZN(_06985_ ) );
INV_X1 _15080_ ( .A(_06204_ ), .ZN(_06986_ ) );
AOI21_X1 _15081_ ( .A(_06985_ ), .B1(_06986_ ), .B2(_06211_ ), .ZN(_06987_ ) );
OR3_X1 _15082_ ( .A1(_06987_ ), .A2(_03859_ ), .A3(_06215_ ), .ZN(_06988_ ) );
OAI21_X1 _15083_ ( .A(_03859_ ), .B1(_06987_ ), .B2(_06215_ ), .ZN(_06989_ ) );
NAND3_X1 _15084_ ( .A1(_06988_ ), .A2(_06561_ ), .A3(_06989_ ), .ZN(_06990_ ) );
NAND3_X1 _15085_ ( .A1(_06971_ ), .A2(_06979_ ), .A3(_06181_ ), .ZN(_06991_ ) );
OR3_X1 _15086_ ( .A1(_03858_ ), .A2(_03241_ ), .A3(_06488_ ), .ZN(_06992_ ) );
AOI21_X1 _15087_ ( .A(_06135_ ), .B1(_03858_ ), .B2(_03241_ ), .ZN(_06993_ ) );
NAND2_X1 _15088_ ( .A1(_06521_ ), .A2(_06708_ ), .ZN(_06994_ ) );
OR2_X1 _15089_ ( .A1(_06509_ ), .A2(_06546_ ), .ZN(_06995_ ) );
AND3_X1 _15090_ ( .A1(_06994_ ), .A2(_06777_ ), .A3(_06995_ ), .ZN(_06996_ ) );
AOI211_X1 _15091_ ( .A(_06993_ ), .B(_06996_ ), .C1(_03859_ ), .C2(_06368_ ), .ZN(_06997_ ) );
AND4_X1 _15092_ ( .A1(_06990_ ), .A2(_06991_ ), .A3(_06992_ ), .A4(_06997_ ), .ZN(_06998_ ) );
AOI21_X1 _15093_ ( .A(_06375_ ), .B1(_06984_ ), .B2(_06998_ ), .ZN(_06999_ ) );
AND2_X1 _15094_ ( .A1(_03318_ ), .A2(_03293_ ), .ZN(_07000_ ) );
AOI21_X1 _15095_ ( .A(_04017_ ), .B1(_04003_ ), .B2(_07000_ ), .ZN(_07001_ ) );
XNOR2_X1 _15096_ ( .A(_03265_ ), .B(_02249_ ), .ZN(_07002_ ) );
NOR2_X1 _15097_ ( .A1(_07001_ ), .A2(_07002_ ), .ZN(_07003_ ) );
OR3_X1 _15098_ ( .A1(_07003_ ), .A2(_03242_ ), .A3(_04020_ ), .ZN(_07004_ ) );
OAI21_X1 _15099_ ( .A(_03242_ ), .B1(_07003_ ), .B2(_04020_ ), .ZN(_07005_ ) );
NAND3_X1 _15100_ ( .A1(_07004_ ), .A2(_06501_ ), .A3(_07005_ ), .ZN(_07006_ ) );
OR2_X1 _15101_ ( .A1(_04449_ ), .A2(_06117_ ), .ZN(_07007_ ) );
NAND3_X1 _15102_ ( .A1(_06127_ ), .A2(\ID_EX_imm [11] ), .A3(_06128_ ), .ZN(_07008_ ) );
AND2_X1 _15103_ ( .A1(_07007_ ), .A2(_07008_ ), .ZN(_07009_ ) );
AOI21_X1 _15104_ ( .A(_06133_ ), .B1(_07006_ ), .B2(_07009_ ), .ZN(_07010_ ) );
NOR3_X1 _15105_ ( .A1(_06999_ ), .A2(_06685_ ), .A3(_07010_ ), .ZN(_07011_ ) );
BUF_X4 _15106_ ( .A(_05861_ ), .Z(_07012_ ) );
OAI21_X1 _15107_ ( .A(_07012_ ), .B1(_04443_ ), .B2(_06729_ ), .ZN(_07013_ ) );
OAI21_X1 _15108_ ( .A(_06969_ ), .B1(_07011_ ), .B2(_07013_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OR2_X1 _15109_ ( .A1(_04498_ ), .A2(_05891_ ), .ZN(_07014_ ) );
AND2_X1 _15110_ ( .A1(_07001_ ), .A2(_07002_ ), .ZN(_07015_ ) );
OR3_X1 _15111_ ( .A1(_07015_ ), .A2(_07003_ ), .A3(_06386_ ), .ZN(_07016_ ) );
AOI22_X1 _15112_ ( .A1(_04506_ ), .A2(_06576_ ), .B1(\ID_EX_imm [10] ), .B2(_06577_ ), .ZN(_07017_ ) );
AOI21_X1 _15113_ ( .A(_06573_ ), .B1(_07016_ ), .B2(_07017_ ), .ZN(_07018_ ) );
OR2_X1 _15114_ ( .A1(_07018_ ), .A2(_01650_ ), .ZN(_07019_ ) );
OAI21_X1 _15115_ ( .A(_06981_ ), .B1(_06583_ ), .B2(_06584_ ), .ZN(_07020_ ) );
NAND3_X1 _15116_ ( .A1(_07020_ ), .A2(_06249_ ), .A3(_06794_ ), .ZN(_07021_ ) );
NOR3_X1 _15117_ ( .A1(_06204_ ), .A2(_03855_ ), .A3(_06212_ ), .ZN(_07022_ ) );
OR3_X1 _15118_ ( .A1(_06987_ ), .A2(_06659_ ), .A3(_07022_ ), .ZN(_07023_ ) );
OAI21_X1 _15119_ ( .A(_06607_ ), .B1(_06799_ ), .B2(_06800_ ), .ZN(_07024_ ) );
NOR3_X1 _15120_ ( .A1(_06465_ ), .A2(_06395_ ), .A3(_06462_ ), .ZN(_07025_ ) );
BUF_X4 _15121_ ( .A(_06342_ ), .Z(_07026_ ) );
NOR3_X1 _15122_ ( .A1(_06444_ ), .A2(_06467_ ), .A3(_07026_ ), .ZN(_07027_ ) );
OAI21_X1 _15123_ ( .A(_06620_ ), .B1(_07025_ ), .B2(_07027_ ), .ZN(_07028_ ) );
NAND2_X1 _15124_ ( .A1(_07024_ ), .A2(_07028_ ), .ZN(_07029_ ) );
NAND2_X1 _15125_ ( .A1(_07029_ ), .A2(_06609_ ), .ZN(_07030_ ) );
OAI211_X1 _15126_ ( .A(_07030_ ), .B(_06530_ ), .C1(_06669_ ), .C2(_06593_ ), .ZN(_07031_ ) );
AOI21_X1 _15127_ ( .A(_03911_ ), .B1(_06594_ ), .B2(_06597_ ), .ZN(_07032_ ) );
OAI211_X1 _15128_ ( .A(_07031_ ), .B(_06767_ ), .C1(_06630_ ), .C2(_07032_ ), .ZN(_07033_ ) );
BUF_X4 _15129_ ( .A(_06367_ ), .Z(_07034_ ) );
NAND3_X1 _15130_ ( .A1(_03946_ ), .A2(_02249_ ), .A3(_07034_ ), .ZN(_07035_ ) );
AOI21_X1 _15131_ ( .A(_06565_ ), .B1(_03854_ ), .B2(_03266_ ), .ZN(_07036_ ) );
AOI21_X1 _15132_ ( .A(_07036_ ), .B1(_03855_ ), .B2(_06567_ ), .ZN(_07037_ ) );
NAND3_X1 _15133_ ( .A1(_06627_ ), .A2(_06624_ ), .A3(_06609_ ), .ZN(_07038_ ) );
OAI21_X1 _15134_ ( .A(_06765_ ), .B1(_06606_ ), .B2(_06607_ ), .ZN(_07039_ ) );
NAND3_X1 _15135_ ( .A1(_07038_ ), .A2(_06778_ ), .A3(_07039_ ), .ZN(_07040_ ) );
AND4_X1 _15136_ ( .A1(_07033_ ), .A2(_07035_ ), .A3(_07037_ ), .A4(_07040_ ), .ZN(_07041_ ) );
NAND3_X1 _15137_ ( .A1(_07021_ ), .A2(_07023_ ), .A3(_07041_ ), .ZN(_07042_ ) );
AOI21_X1 _15138_ ( .A(_07019_ ), .B1(_07042_ ), .B2(_06377_ ), .ZN(_07043_ ) );
OAI21_X1 _15139_ ( .A(_07012_ ), .B1(_04501_ ), .B2(_06729_ ), .ZN(_07044_ ) );
OAI21_X1 _15140_ ( .A(_07014_ ), .B1(_07043_ ), .B2(_07044_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
INV_X1 _15141_ ( .A(_05972_ ), .ZN(_07045_ ) );
NOR3_X1 _15142_ ( .A1(_06340_ ), .A2(_06318_ ), .A3(_06330_ ), .ZN(_07046_ ) );
NOR3_X1 _15143_ ( .A1(_06337_ ), .A2(_06341_ ), .A3(_06342_ ), .ZN(_07047_ ) );
NOR3_X1 _15144_ ( .A1(_07046_ ), .A2(_07047_ ), .A3(_06325_ ), .ZN(_07048_ ) );
AOI21_X1 _15145_ ( .A(_06349_ ), .B1(_06844_ ), .B2(_06845_ ), .ZN(_07049_ ) );
OAI21_X1 _15146_ ( .A(_06708_ ), .B1(_07048_ ), .B2(_07049_ ), .ZN(_07050_ ) );
NAND3_X1 _15147_ ( .A1(_06652_ ), .A2(_06655_ ), .A3(_06345_ ), .ZN(_07051_ ) );
AND3_X1 _15148_ ( .A1(_07050_ ), .A2(_06178_ ), .A3(_07051_ ), .ZN(_07052_ ) );
AND4_X1 _15149_ ( .A1(_06443_ ), .A2(_06649_ ), .A3(_06650_ ), .A4(_06668_ ), .ZN(_07053_ ) );
AOI211_X1 _15150_ ( .A(_07052_ ), .B(_07053_ ), .C1(_06788_ ), .C2(_06794_ ), .ZN(_07054_ ) );
NAND4_X1 _15151_ ( .A1(_06582_ ), .A2(_06296_ ), .A3(_06299_ ), .A4(_06794_ ), .ZN(_07055_ ) );
AOI21_X1 _15152_ ( .A(_06394_ ), .B1(_07054_ ), .B2(_07055_ ), .ZN(_07056_ ) );
OR2_X1 _15153_ ( .A1(_06203_ ), .A2(_03870_ ), .ZN(_07057_ ) );
INV_X1 _15154_ ( .A(_06209_ ), .ZN(_07058_ ) );
AND3_X1 _15155_ ( .A1(_07057_ ), .A2(_03865_ ), .A3(_07058_ ), .ZN(_07059_ ) );
AOI21_X1 _15156_ ( .A(_03865_ ), .B1(_07057_ ), .B2(_07058_ ), .ZN(_07060_ ) );
OR3_X1 _15157_ ( .A1(_07059_ ), .A2(_07060_ ), .A3(_06634_ ), .ZN(_07061_ ) );
OAI21_X1 _15158_ ( .A(_06818_ ), .B1(_07052_ ), .B2(_07053_ ), .ZN(_07062_ ) );
AOI22_X1 _15159_ ( .A1(_03864_ ), .A2(_06567_ ), .B1(_03939_ ), .B2(_07034_ ), .ZN(_07063_ ) );
NAND2_X1 _15160_ ( .A1(_06672_ ), .A2(_06609_ ), .ZN(_07064_ ) );
NAND3_X1 _15161_ ( .A1(_06320_ ), .A2(_06765_ ), .A3(_06674_ ), .ZN(_07065_ ) );
NAND2_X1 _15162_ ( .A1(_07064_ ), .A2(_07065_ ), .ZN(_07066_ ) );
AOI22_X1 _15163_ ( .A1(_07066_ ), .A2(_06778_ ), .B1(_06210_ ), .B2(_06486_ ), .ZN(_07067_ ) );
NAND4_X1 _15164_ ( .A1(_07061_ ), .A2(_07062_ ), .A3(_07063_ ), .A4(_07067_ ), .ZN(_07068_ ) );
OAI21_X1 _15165_ ( .A(_06376_ ), .B1(_07056_ ), .B2(_07068_ ), .ZN(_07069_ ) );
NAND2_X1 _15166_ ( .A1(_03316_ ), .A2(_02202_ ), .ZN(_07070_ ) );
NOR2_X1 _15167_ ( .A1(_03316_ ), .A2(_02202_ ), .ZN(_07071_ ) );
OAI21_X1 _15168_ ( .A(_07070_ ), .B1(_04002_ ), .B2(_07071_ ), .ZN(_07072_ ) );
AOI21_X1 _15169_ ( .A(_06387_ ), .B1(_07072_ ), .B2(_03293_ ), .ZN(_07073_ ) );
OAI21_X1 _15170_ ( .A(_07073_ ), .B1(_03293_ ), .B2(_07072_ ), .ZN(_07074_ ) );
OR2_X1 _15171_ ( .A1(_04531_ ), .A2(_06117_ ), .ZN(_07075_ ) );
NAND3_X1 _15172_ ( .A1(_06127_ ), .A2(\ID_EX_imm [9] ), .A3(_06128_ ), .ZN(_07076_ ) );
NAND3_X1 _15173_ ( .A1(_07074_ ), .A2(_07075_ ), .A3(_07076_ ), .ZN(_07077_ ) );
NAND2_X1 _15174_ ( .A1(_07077_ ), .A2(_06381_ ), .ZN(_07078_ ) );
AND3_X1 _15175_ ( .A1(_07069_ ), .A2(_06391_ ), .A3(_07078_ ), .ZN(_07079_ ) );
NAND2_X1 _15176_ ( .A1(_04528_ ), .A2(_06685_ ), .ZN(_07080_ ) );
NAND2_X1 _15177_ ( .A1(_07080_ ), .A2(_05862_ ), .ZN(_07081_ ) );
OAI21_X1 _15178_ ( .A(_07045_ ), .B1(_07079_ ), .B2(_07081_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
NOR2_X1 _15179_ ( .A1(_06251_ ), .A2(_06345_ ), .ZN(_07082_ ) );
INV_X1 _15180_ ( .A(_07082_ ), .ZN(_07083_ ) );
NAND4_X1 _15181_ ( .A1(_06646_ ), .A2(_06292_ ), .A3(_07083_ ), .A4(_06289_ ), .ZN(_07084_ ) );
OR3_X1 _15182_ ( .A1(_06621_ ), .A2(_06157_ ), .A3(_06475_ ), .ZN(_07085_ ) );
NAND3_X1 _15183_ ( .A1(_06466_ ), .A2(_06157_ ), .A3(_06463_ ), .ZN(_07086_ ) );
AND2_X1 _15184_ ( .A1(_07085_ ), .A2(_07086_ ), .ZN(_07087_ ) );
MUX2_X1 _15185_ ( .A(_06881_ ), .B(_07087_ ), .S(_03908_ ), .Z(_07088_ ) );
NAND2_X1 _15186_ ( .A1(_07088_ ), .A2(_06546_ ), .ZN(_07089_ ) );
OAI211_X1 _15187_ ( .A(_07089_ ), .B(_06322_ ), .C1(_06510_ ), .C2(_06697_ ), .ZN(_07090_ ) );
NAND3_X1 _15188_ ( .A1(_06699_ ), .A2(_06442_ ), .A3(_06708_ ), .ZN(_07091_ ) );
AND2_X1 _15189_ ( .A1(_07090_ ), .A2(_07091_ ), .ZN(_07092_ ) );
AOI21_X1 _15190_ ( .A(_06394_ ), .B1(_07084_ ), .B2(_07092_ ), .ZN(_07093_ ) );
AOI21_X1 _15191_ ( .A(_06887_ ), .B1(_07090_ ), .B2(_07091_ ), .ZN(_07094_ ) );
NAND2_X1 _15192_ ( .A1(_06717_ ), .A2(_06668_ ), .ZN(_07095_ ) );
OR2_X1 _15193_ ( .A1(_06707_ ), .A2(_06510_ ), .ZN(_07096_ ) );
AND3_X1 _15194_ ( .A1(_07095_ ), .A2(_06777_ ), .A3(_07096_ ), .ZN(_07097_ ) );
OR3_X1 _15195_ ( .A1(_07093_ ), .A2(_07094_ ), .A3(_07097_ ), .ZN(_07098_ ) );
OAI21_X1 _15196_ ( .A(_06245_ ), .B1(_06203_ ), .B2(_03870_ ), .ZN(_07099_ ) );
AOI21_X1 _15197_ ( .A(_07099_ ), .B1(_03870_ ), .B2(_06203_ ), .ZN(_07100_ ) );
NAND3_X1 _15198_ ( .A1(_03866_ ), .A2(_03317_ ), .A3(_03867_ ), .ZN(_07101_ ) );
AOI22_X1 _15199_ ( .A1(_06209_ ), .A2(_07034_ ), .B1(_07101_ ), .B2(_06486_ ), .ZN(_07102_ ) );
OAI21_X1 _15200_ ( .A(_07102_ ), .B1(_03870_ ), .B2(_03987_ ), .ZN(_07103_ ) );
NOR3_X1 _15201_ ( .A1(_07098_ ), .A2(_07100_ ), .A3(_07103_ ), .ZN(_07104_ ) );
NOR2_X1 _15202_ ( .A1(_07104_ ), .A2(_06375_ ), .ZN(_07105_ ) );
AOI21_X1 _15203_ ( .A(_06387_ ), .B1(_04003_ ), .B2(_03318_ ), .ZN(_07106_ ) );
OAI21_X1 _15204_ ( .A(_07106_ ), .B1(_03318_ ), .B2(_04003_ ), .ZN(_07107_ ) );
AOI22_X1 _15205_ ( .A1(_04556_ ), .A2(_06576_ ), .B1(\ID_EX_imm [8] ), .B2(_06577_ ), .ZN(_07108_ ) );
AOI21_X1 _15206_ ( .A(_06573_ ), .B1(_07107_ ), .B2(_07108_ ), .ZN(_07109_ ) );
OR2_X1 _15207_ ( .A1(_07109_ ), .A2(_06685_ ), .ZN(_07110_ ) );
OAI221_X1 _15208_ ( .A(_05888_ ), .B1(_06391_ ), .B2(_04554_ ), .C1(_07105_ ), .C2(_07110_ ), .ZN(_07111_ ) );
NAND3_X1 _15209_ ( .A1(_04548_ ), .A2(_05879_ ), .A3(_04550_ ), .ZN(_07112_ ) );
NAND2_X1 _15210_ ( .A1(_07111_ ), .A2(_07112_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
OAI21_X1 _15211_ ( .A(_05916_ ), .B1(_04566_ ), .B2(_04573_ ), .ZN(_07113_ ) );
AND2_X1 _15212_ ( .A1(_03994_ ), .A2(_03995_ ), .ZN(_07114_ ) );
AOI21_X1 _15213_ ( .A(_04000_ ), .B1(_07114_ ), .B2(_03422_ ), .ZN(_07115_ ) );
INV_X1 _15214_ ( .A(_03374_ ), .ZN(_07116_ ) );
NOR2_X1 _15215_ ( .A1(_07115_ ), .A2(_07116_ ), .ZN(_07117_ ) );
AOI21_X1 _15216_ ( .A(_07117_ ), .B1(_02171_ ), .B2(_03373_ ), .ZN(_07118_ ) );
XNOR2_X1 _15217_ ( .A(_07118_ ), .B(_03343_ ), .ZN(_07119_ ) );
NAND2_X1 _15218_ ( .A1(_07119_ ), .A2(_06501_ ), .ZN(_07120_ ) );
OR2_X1 _15219_ ( .A1(_04580_ ), .A2(_06117_ ), .ZN(_07121_ ) );
NAND3_X1 _15220_ ( .A1(_06127_ ), .A2(\ID_EX_imm [7] ), .A3(_06128_ ), .ZN(_07122_ ) );
AND3_X1 _15221_ ( .A1(_07120_ ), .A2(_07121_ ), .A3(_07122_ ), .ZN(_07123_ ) );
OAI21_X1 _15222_ ( .A(_01654_ ), .B1(_07123_ ), .B2(_06133_ ), .ZN(_07124_ ) );
NAND4_X1 _15223_ ( .A1(_06646_ ), .A2(_06248_ ), .A3(_06301_ ), .A4(_06794_ ), .ZN(_07125_ ) );
NAND2_X1 _15224_ ( .A1(_06201_ ), .A2(_06195_ ), .ZN(_07126_ ) );
NOR2_X1 _15225_ ( .A1(_07126_ ), .A2(_03899_ ), .ZN(_07127_ ) );
NOR3_X1 _15226_ ( .A1(_07127_ ), .A2(_03890_ ), .A3(_06189_ ), .ZN(_07128_ ) );
OR3_X1 _15227_ ( .A1(_07128_ ), .A2(_03883_ ), .A3(_03892_ ), .ZN(_07129_ ) );
AND3_X1 _15228_ ( .A1(_07129_ ), .A2(_03878_ ), .A3(_06186_ ), .ZN(_07130_ ) );
AOI21_X1 _15229_ ( .A(_03878_ ), .B1(_07129_ ), .B2(_06186_ ), .ZN(_07131_ ) );
OR3_X1 _15230_ ( .A1(_07130_ ), .A2(_07131_ ), .A3(_06659_ ), .ZN(_07132_ ) );
OR3_X1 _15231_ ( .A1(_06328_ ), .A2(_06318_ ), .A3(_06333_ ), .ZN(_07133_ ) );
OR3_X1 _15232_ ( .A1(_06340_ ), .A2(_06330_ ), .A3(_06151_ ), .ZN(_07134_ ) );
AND3_X1 _15233_ ( .A1(_07133_ ), .A2(_07134_ ), .A3(_06317_ ), .ZN(_07135_ ) );
NOR3_X1 _15234_ ( .A1(_06973_ ), .A2(_06974_ ), .A3(_06317_ ), .ZN(_07136_ ) );
NOR3_X1 _15235_ ( .A1(_07135_ ), .A2(_06345_ ), .A3(_07136_ ), .ZN(_07137_ ) );
AOI21_X1 _15236_ ( .A(_06510_ ), .B1(_06760_ ), .B2(_06763_ ), .ZN(_07138_ ) );
OR3_X1 _15237_ ( .A1(_07137_ ), .A2(_06443_ ), .A3(_07138_ ), .ZN(_07139_ ) );
MUX2_X1 _15238_ ( .A(_06768_ ), .B(_06758_ ), .S(_06510_ ), .Z(_07140_ ) );
OAI211_X1 _15239_ ( .A(_07139_ ), .B(_06767_ ), .C1(_06630_ ), .C2(_07140_ ), .ZN(_07141_ ) );
NOR2_X1 _15240_ ( .A1(_06771_ ), .A2(_06772_ ), .ZN(_07142_ ) );
INV_X1 _15241_ ( .A(_06777_ ), .ZN(_07143_ ) );
OR3_X1 _15242_ ( .A1(_07142_ ), .A2(_06842_ ), .A3(_07143_ ), .ZN(_07144_ ) );
OR3_X1 _15243_ ( .A1(_03874_ ), .A2(_03342_ ), .A3(_06488_ ), .ZN(_07145_ ) );
NOR2_X1 _15244_ ( .A1(_03876_ ), .A2(_06565_ ), .ZN(_07146_ ) );
AOI21_X1 _15245_ ( .A(_07146_ ), .B1(_03877_ ), .B2(_06368_ ), .ZN(_07147_ ) );
AND4_X1 _15246_ ( .A1(_07141_ ), .A2(_07144_ ), .A3(_07145_ ), .A4(_07147_ ), .ZN(_07148_ ) );
NAND3_X1 _15247_ ( .A1(_07125_ ), .A2(_07132_ ), .A3(_07148_ ), .ZN(_07149_ ) );
AOI21_X1 _15248_ ( .A(_07124_ ), .B1(_07149_ ), .B2(_06377_ ), .ZN(_07150_ ) );
OAI21_X1 _15249_ ( .A(_07012_ ), .B1(_04576_ ), .B2(_06729_ ), .ZN(_07151_ ) );
OAI21_X1 _15250_ ( .A(_07113_ ), .B1(_07150_ ), .B2(_07151_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
OR3_X1 _15251_ ( .A1(_04603_ ), .A2(_05861_ ), .A3(_04605_ ), .ZN(_07152_ ) );
AND3_X1 _15252_ ( .A1(_06793_ ), .A2(_06301_ ), .A3(_06789_ ), .ZN(_07153_ ) );
MUX2_X1 _15253_ ( .A(_06805_ ), .B(_06797_ ), .S(_06510_ ), .Z(_07154_ ) );
NAND2_X1 _15254_ ( .A1(_07154_ ), .A2(_06443_ ), .ZN(_07155_ ) );
OAI21_X1 _15255_ ( .A(_06607_ ), .B1(_07025_ ), .B2(_07027_ ), .ZN(_07156_ ) );
OAI21_X1 _15256_ ( .A(_07026_ ), .B1(_06474_ ), .B2(_06472_ ), .ZN(_07157_ ) );
OAI21_X1 _15257_ ( .A(_06395_ ), .B1(_06621_ ), .B2(_06475_ ), .ZN(_07158_ ) );
NAND3_X1 _15258_ ( .A1(_07157_ ), .A2(_07158_ ), .A3(_06620_ ), .ZN(_07159_ ) );
NAND3_X1 _15259_ ( .A1(_07156_ ), .A2(_06668_ ), .A3(_07159_ ), .ZN(_07160_ ) );
NAND3_X1 _15260_ ( .A1(_06801_ ), .A2(_06364_ ), .A3(_06802_ ), .ZN(_07161_ ) );
NAND3_X1 _15261_ ( .A1(_07160_ ), .A2(_07161_ ), .A3(_06425_ ), .ZN(_07162_ ) );
NAND2_X1 _15262_ ( .A1(_07155_ ), .A2(_07162_ ), .ZN(_07163_ ) );
OAI21_X1 _15263_ ( .A(_06248_ ), .B1(_07153_ ), .B2(_07163_ ), .ZN(_07164_ ) );
OAI21_X1 _15264_ ( .A(_03883_ ), .B1(_07128_ ), .B2(_03892_ ), .ZN(_07165_ ) );
NAND3_X1 _15265_ ( .A1(_07129_ ), .A2(_06561_ ), .A3(_07165_ ), .ZN(_07166_ ) );
NAND2_X1 _15266_ ( .A1(_07163_ ), .A2(_06818_ ), .ZN(_07167_ ) );
NOR3_X1 _15267_ ( .A1(_06811_ ), .A2(_06323_ ), .A3(_07143_ ), .ZN(_07168_ ) );
NAND3_X1 _15268_ ( .A1(_03344_ ), .A2(_03879_ ), .A3(_03880_ ), .ZN(_07169_ ) );
AOI221_X4 _15269_ ( .A(_07168_ ), .B1(_07169_ ), .B2(_04075_ ), .C1(_03882_ ), .C2(_03986_ ), .ZN(_07170_ ) );
AND4_X1 _15270_ ( .A1(_07164_ ), .A2(_07166_ ), .A3(_07167_ ), .A4(_07170_ ), .ZN(_07171_ ) );
OR3_X1 _15271_ ( .A1(_03881_ ), .A2(_03344_ ), .A3(_06488_ ), .ZN(_07172_ ) );
AOI21_X1 _15272_ ( .A(_06375_ ), .B1(_07171_ ), .B2(_07172_ ), .ZN(_07173_ ) );
AND2_X1 _15273_ ( .A1(_07115_ ), .A2(_07116_ ), .ZN(_07174_ ) );
OR3_X1 _15274_ ( .A1(_07174_ ), .A2(_07117_ ), .A3(_06387_ ), .ZN(_07175_ ) );
AOI22_X1 _15275_ ( .A1(_04621_ ), .A2(_06576_ ), .B1(\ID_EX_imm [6] ), .B2(_06577_ ), .ZN(_07176_ ) );
AOI21_X1 _15276_ ( .A(_06133_ ), .B1(_07175_ ), .B2(_07176_ ), .ZN(_07177_ ) );
NOR3_X1 _15277_ ( .A1(_07173_ ), .A2(_06685_ ), .A3(_07177_ ), .ZN(_07178_ ) );
OAI21_X1 _15278_ ( .A(_07012_ ), .B1(_04619_ ), .B2(_06729_ ), .ZN(_07179_ ) );
OAI21_X1 _15279_ ( .A(_07152_ ), .B1(_07178_ ), .B2(_07179_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
AND2_X1 _15280_ ( .A1(_04638_ ), .A2(_01649_ ), .ZN(_07180_ ) );
AND4_X1 _15281_ ( .A1(_06298_ ), .A2(_06288_ ), .A3(_06300_ ), .A4(_06789_ ), .ZN(_07181_ ) );
NAND2_X1 _15282_ ( .A1(_06176_ ), .A2(_06442_ ), .ZN(_07182_ ) );
OAI21_X1 _15283_ ( .A(_06297_ ), .B1(_07046_ ), .B2(_07047_ ), .ZN(_07183_ ) );
OAI21_X1 _15284_ ( .A(_06334_ ), .B1(_06332_ ), .B2(_06310_ ), .ZN(_07184_ ) );
OAI21_X1 _15285_ ( .A(_06329_ ), .B1(_06328_ ), .B2(_06333_ ), .ZN(_07185_ ) );
NAND3_X1 _15286_ ( .A1(_07184_ ), .A2(_07185_ ), .A3(_06349_ ), .ZN(_07186_ ) );
NAND3_X1 _15287_ ( .A1(_07183_ ), .A2(_06546_ ), .A3(_07186_ ), .ZN(_07187_ ) );
NAND3_X1 _15288_ ( .A1(_06843_ ), .A2(_06846_ ), .A3(_06323_ ), .ZN(_07188_ ) );
NAND3_X1 _15289_ ( .A1(_07187_ ), .A2(_06322_ ), .A3(_07188_ ), .ZN(_07189_ ) );
NAND2_X1 _15290_ ( .A1(_07182_ ), .A2(_07189_ ), .ZN(_07190_ ) );
OAI21_X1 _15291_ ( .A(_06247_ ), .B1(_07181_ ), .B2(_07190_ ), .ZN(_07191_ ) );
NAND2_X1 _15292_ ( .A1(_07190_ ), .A2(_06181_ ), .ZN(_07192_ ) );
OR3_X1 _15293_ ( .A1(_06321_ ), .A2(_06345_ ), .A3(_07143_ ), .ZN(_07193_ ) );
AND3_X1 _15294_ ( .A1(_07191_ ), .A2(_07192_ ), .A3(_07193_ ), .ZN(_07194_ ) );
NAND2_X1 _15295_ ( .A1(_03896_ ), .A2(_06567_ ), .ZN(_07195_ ) );
NAND3_X1 _15296_ ( .A1(_03889_ ), .A2(_02096_ ), .A3(_07034_ ), .ZN(_07196_ ) );
OAI21_X1 _15297_ ( .A(_06486_ ), .B1(_03889_ ), .B2(_02096_ ), .ZN(_07197_ ) );
NAND4_X1 _15298_ ( .A1(_07194_ ), .A2(_07195_ ), .A3(_07196_ ), .A4(_07197_ ), .ZN(_07198_ ) );
OR3_X1 _15299_ ( .A1(_07127_ ), .A2(_03896_ ), .A3(_06189_ ), .ZN(_07199_ ) );
OAI21_X1 _15300_ ( .A(_03896_ ), .B1(_07127_ ), .B2(_06189_ ), .ZN(_07200_ ) );
AND3_X1 _15301_ ( .A1(_07199_ ), .A2(_06245_ ), .A3(_07200_ ), .ZN(_07201_ ) );
OAI21_X1 _15302_ ( .A(_06376_ ), .B1(_07198_ ), .B2(_07201_ ), .ZN(_07202_ ) );
AND3_X1 _15303_ ( .A1(_03994_ ), .A2(_03995_ ), .A3(_03421_ ), .ZN(_07203_ ) );
OR3_X1 _15304_ ( .A1(_07203_ ), .A2(_03398_ ), .A3(_03998_ ), .ZN(_07204_ ) );
OAI21_X1 _15305_ ( .A(_03398_ ), .B1(_07203_ ), .B2(_03998_ ), .ZN(_07205_ ) );
NAND3_X1 _15306_ ( .A1(_07204_ ), .A2(_06501_ ), .A3(_07205_ ), .ZN(_07206_ ) );
OR2_X1 _15307_ ( .A1(_04642_ ), .A2(_06117_ ), .ZN(_07207_ ) );
NAND3_X1 _15308_ ( .A1(_06127_ ), .A2(\ID_EX_imm [5] ), .A3(_06128_ ), .ZN(_07208_ ) );
NAND3_X1 _15309_ ( .A1(_07206_ ), .A2(_07207_ ), .A3(_07208_ ), .ZN(_07209_ ) );
AOI21_X1 _15310_ ( .A(_01650_ ), .B1(_07209_ ), .B2(_06381_ ), .ZN(_07210_ ) );
AOI21_X1 _15311_ ( .A(_07180_ ), .B1(_07202_ ), .B2(_07210_ ), .ZN(_07211_ ) );
MUX2_X1 _15312_ ( .A(_04636_ ), .B(_07211_ ), .S(_05867_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
OR3_X1 _15313_ ( .A1(_04667_ ), .A2(_05861_ ), .A3(_04669_ ), .ZN(_07212_ ) );
NAND4_X1 _15314_ ( .A1(_06646_ ), .A2(_06301_ ), .A3(_06397_ ), .A4(_06794_ ), .ZN(_07213_ ) );
OR2_X1 _15315_ ( .A1(_07087_ ), .A2(_06349_ ), .ZN(_07214_ ) );
NOR3_X1 _15316_ ( .A1(_06471_ ), .A2(_06157_ ), .A3(_06436_ ), .ZN(_07215_ ) );
NOR3_X1 _15317_ ( .A1(_06474_ ), .A2(_06472_ ), .A3(_06145_ ), .ZN(_07216_ ) );
OAI21_X1 _15318_ ( .A(_06317_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07217_ ) );
AND3_X1 _15319_ ( .A1(_07214_ ), .A2(_06510_ ), .A3(_07217_ ), .ZN(_07218_ ) );
AOI211_X1 _15320_ ( .A(_06443_ ), .B(_07218_ ), .C1(_06842_ ), .C2(_06883_ ), .ZN(_07219_ ) );
AND2_X1 _15321_ ( .A1(_06424_ ), .A2(_06443_ ), .ZN(_07220_ ) );
NOR2_X1 _15322_ ( .A1(_07219_ ), .A2(_07220_ ), .ZN(_07221_ ) );
AOI21_X1 _15323_ ( .A(_06394_ ), .B1(_07213_ ), .B2(_07221_ ), .ZN(_07222_ ) );
OAI21_X1 _15324_ ( .A(_06818_ ), .B1(_07219_ ), .B2(_07220_ ), .ZN(_07223_ ) );
AOI21_X1 _15325_ ( .A(_06634_ ), .B1(_07126_ ), .B2(_03899_ ), .ZN(_07224_ ) );
OAI21_X1 _15326_ ( .A(_07224_ ), .B1(_03899_ ), .B2(_07126_ ), .ZN(_07225_ ) );
NAND3_X1 _15327_ ( .A1(_06600_ ), .A2(_02118_ ), .A3(_07034_ ), .ZN(_07226_ ) );
AOI21_X1 _15328_ ( .A(_06135_ ), .B1(_06322_ ), .B2(_02123_ ), .ZN(_07227_ ) );
AOI221_X4 _15329_ ( .A(_07227_ ), .B1(_03898_ ), .B2(_03986_ ), .C1(_06440_ ), .C2(_06777_ ), .ZN(_07228_ ) );
NAND4_X1 _15330_ ( .A1(_07223_ ), .A2(_07225_ ), .A3(_07226_ ), .A4(_07228_ ), .ZN(_07229_ ) );
OAI21_X1 _15331_ ( .A(_06376_ ), .B1(_07222_ ), .B2(_07229_ ), .ZN(_07230_ ) );
AOI21_X1 _15332_ ( .A(_03421_ ), .B1(_03994_ ), .B2(_03995_ ), .ZN(_07231_ ) );
NOR3_X1 _15333_ ( .A1(_07203_ ), .A2(_07231_ ), .A3(_06387_ ), .ZN(_07232_ ) );
OAI22_X1 _15334_ ( .A1(_04675_ ), .A2(_06118_ ), .B1(_02119_ ), .B2(_06383_ ), .ZN(_07233_ ) );
OAI21_X1 _15335_ ( .A(_06381_ ), .B1(_07232_ ), .B2(_07233_ ), .ZN(_07234_ ) );
AND3_X1 _15336_ ( .A1(_07230_ ), .A2(_06391_ ), .A3(_07234_ ), .ZN(_07235_ ) );
OAI21_X1 _15337_ ( .A(_07012_ ), .B1(_01655_ ), .B2(_04673_ ), .ZN(_07236_ ) );
OAI21_X1 _15338_ ( .A(_07212_ ), .B1(_07235_ ), .B2(_07236_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
OR3_X1 _15339_ ( .A1(_04696_ ), .A2(_05861_ ), .A3(_04698_ ), .ZN(_07237_ ) );
OR2_X1 _15340_ ( .A1(_03993_ ), .A2(_03719_ ), .ZN(_07238_ ) );
AND3_X1 _15341_ ( .A1(_07238_ ), .A2(_03693_ ), .A3(_03989_ ), .ZN(_07239_ ) );
AOI21_X1 _15342_ ( .A(_03693_ ), .B1(_07238_ ), .B2(_03989_ ), .ZN(_07240_ ) );
OR3_X1 _15343_ ( .A1(_07239_ ), .A2(_07240_ ), .A3(_06386_ ), .ZN(_07241_ ) );
AOI22_X1 _15344_ ( .A1(_04704_ ), .A2(_06576_ ), .B1(\ID_EX_imm [3] ), .B2(_06577_ ), .ZN(_07242_ ) );
AOI21_X1 _15345_ ( .A(_06573_ ), .B1(_07241_ ), .B2(_07242_ ), .ZN(_07243_ ) );
OR2_X1 _15346_ ( .A1(_07243_ ), .A2(_01650_ ), .ZN(_07244_ ) );
NAND2_X1 _15347_ ( .A1(_06547_ ), .A2(_06443_ ), .ZN(_07245_ ) );
OAI21_X1 _15348_ ( .A(_06395_ ), .B1(_06332_ ), .B2(_06310_ ), .ZN(_07246_ ) );
NOR2_X1 _15349_ ( .A1(_06308_ ), .A2(_06313_ ), .ZN(_07247_ ) );
OAI211_X1 _15350_ ( .A(_07246_ ), .B(_06349_ ), .C1(_07247_ ), .C2(_06395_ ), .ZN(_07248_ ) );
AND2_X1 _15351_ ( .A1(_07133_ ), .A2(_07134_ ), .ZN(_07249_ ) );
OAI211_X1 _15352_ ( .A(_06510_ ), .B(_07248_ ), .C1(_07249_ ), .C2(_06620_ ), .ZN(_07250_ ) );
OAI211_X1 _15353_ ( .A(_07250_ ), .B(_06322_ ), .C1(_06668_ ), .C2(_06976_ ), .ZN(_07251_ ) );
AOI21_X1 _15354_ ( .A(_06887_ ), .B1(_07245_ ), .B2(_07251_ ), .ZN(_07252_ ) );
AND3_X1 _15355_ ( .A1(_06288_ ), .A2(_06300_ ), .A3(_06550_ ), .ZN(_07253_ ) );
NAND2_X1 _15356_ ( .A1(_07253_ ), .A2(_06789_ ), .ZN(_07254_ ) );
NAND3_X1 _15357_ ( .A1(_07254_ ), .A2(_07251_ ), .A3(_07245_ ), .ZN(_07255_ ) );
AOI221_X4 _15358_ ( .A(_07252_ ), .B1(_06511_ ), .B2(_06778_ ), .C1(_07255_ ), .C2(_06248_ ), .ZN(_07256_ ) );
NOR2_X1 _15359_ ( .A1(_06200_ ), .A2(_03915_ ), .ZN(_07257_ ) );
OAI21_X1 _15360_ ( .A(_03905_ ), .B1(_07257_ ), .B2(_06196_ ), .ZN(_07258_ ) );
OAI221_X1 _15361_ ( .A(_06197_ ), .B1(_03916_ ), .B2(_03917_ ), .C1(_06200_ ), .C2(_03915_ ), .ZN(_07259_ ) );
NAND3_X1 _15362_ ( .A1(_07258_ ), .A2(_06561_ ), .A3(_07259_ ), .ZN(_07260_ ) );
AND3_X1 _15363_ ( .A1(_06765_ ), .A2(_02069_ ), .A3(_06367_ ), .ZN(_07261_ ) );
AOI221_X4 _15364_ ( .A(_07261_ ), .B1(_06195_ ), .B2(_06486_ ), .C1(_03905_ ), .C2(_06368_ ), .ZN(_07262_ ) );
NAND3_X1 _15365_ ( .A1(_07256_ ), .A2(_07260_ ), .A3(_07262_ ), .ZN(_07263_ ) );
AOI21_X1 _15366_ ( .A(_07244_ ), .B1(_07263_ ), .B2(_06377_ ), .ZN(_07264_ ) );
OAI21_X1 _15367_ ( .A(_07012_ ), .B1(_01655_ ), .B2(_04701_ ), .ZN(_07265_ ) );
OAI21_X1 _15368_ ( .A(_07237_ ), .B1(_07264_ ), .B2(_07265_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
OR2_X1 _15369_ ( .A1(_04728_ ), .A2(_05891_ ), .ZN(_07266_ ) );
NAND2_X1 _15370_ ( .A1(_03993_ ), .A2(_03719_ ), .ZN(_07267_ ) );
NAND3_X1 _15371_ ( .A1(_07238_ ), .A2(_06501_ ), .A3(_07267_ ), .ZN(_07268_ ) );
AOI22_X1 _15372_ ( .A1(_04731_ ), .A2(_06576_ ), .B1(\ID_EX_imm [2] ), .B2(_06577_ ), .ZN(_07269_ ) );
AOI21_X1 _15373_ ( .A(_06573_ ), .B1(_07268_ ), .B2(_07269_ ), .ZN(_07270_ ) );
OR2_X1 _15374_ ( .A1(_07270_ ), .A2(_01650_ ), .ZN(_07271_ ) );
NOR4_X1 _15375_ ( .A1(_06583_ ), .A2(_06584_ ), .A3(_06299_ ), .A4(_06982_ ), .ZN(_07272_ ) );
OR2_X1 _15376_ ( .A1(_06599_ ), .A2(_06667_ ), .ZN(_07273_ ) );
NOR3_X1 _15377_ ( .A1(_06471_ ), .A2(_07026_ ), .A3(_06436_ ), .ZN(_07274_ ) );
NOR2_X1 _15378_ ( .A1(_06435_ ), .A2(_06433_ ), .ZN(_07275_ ) );
AOI211_X1 _15379_ ( .A(_06607_ ), .B(_07274_ ), .C1(_07026_ ), .C2(_07275_ ), .ZN(_07276_ ) );
AOI21_X1 _15380_ ( .A(_06674_ ), .B1(_07157_ ), .B2(_07158_ ), .ZN(_07277_ ) );
OAI21_X1 _15381_ ( .A(_06669_ ), .B1(_07276_ ), .B2(_07277_ ), .ZN(_07278_ ) );
OAI211_X1 _15382_ ( .A(_07278_ ), .B(_06630_ ), .C1(_06669_ ), .C2(_07029_ ), .ZN(_07279_ ) );
NAND2_X1 _15383_ ( .A1(_07273_ ), .A2(_07279_ ), .ZN(_07280_ ) );
OAI21_X1 _15384_ ( .A(_06249_ ), .B1(_07272_ ), .B2(_07280_ ), .ZN(_07281_ ) );
NAND2_X1 _15385_ ( .A1(_07280_ ), .A2(_06818_ ), .ZN(_07282_ ) );
NAND3_X1 _15386_ ( .A1(_06608_ ), .A2(_06669_ ), .A3(_06778_ ), .ZN(_07283_ ) );
AOI21_X1 _15387_ ( .A(_06634_ ), .B1(_06200_ ), .B2(_03915_ ), .ZN(_07284_ ) );
OAI21_X1 _15388_ ( .A(_07284_ ), .B1(_03915_ ), .B2(_06200_ ), .ZN(_07285_ ) );
NAND3_X1 _15389_ ( .A1(_06607_ ), .A2(_02045_ ), .A3(_07034_ ), .ZN(_07286_ ) );
AOI21_X1 _15390_ ( .A(_06135_ ), .B1(_06674_ ), .B2(_03717_ ), .ZN(_07287_ ) );
AOI21_X1 _15391_ ( .A(_07287_ ), .B1(_03914_ ), .B2(_06368_ ), .ZN(_07288_ ) );
AND4_X1 _15392_ ( .A1(_07283_ ), .A2(_07285_ ), .A3(_07286_ ), .A4(_07288_ ), .ZN(_07289_ ) );
NAND3_X1 _15393_ ( .A1(_07281_ ), .A2(_07282_ ), .A3(_07289_ ), .ZN(_07290_ ) );
BUF_X4 _15394_ ( .A(_06376_ ), .Z(_07291_ ) );
AOI21_X1 _15395_ ( .A(_07271_ ), .B1(_07290_ ), .B2(_07291_ ), .ZN(_07292_ ) );
OAI21_X1 _15396_ ( .A(_07012_ ), .B1(_01655_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07293_ ) );
OAI21_X1 _15397_ ( .A(_07266_ ), .B1(_07292_ ), .B2(_07293_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
OR2_X1 _15398_ ( .A1(_02665_ ), .A2(\EX_LS_result_csreg_mem [29] ), .ZN(_07294_ ) );
INV_X1 _15399_ ( .A(_04165_ ), .ZN(_07295_ ) );
OAI211_X1 _15400_ ( .A(_07294_ ), .B(_05909_ ), .C1(_07295_ ), .C2(_04142_ ), .ZN(_07296_ ) );
OAI22_X1 _15401_ ( .A1(_04128_ ), .A2(_06118_ ), .B1(_02540_ ), .B2(_06383_ ), .ZN(_07297_ ) );
NOR2_X1 _15402_ ( .A1(_06905_ ), .A2(_06907_ ), .ZN(_07298_ ) );
OR3_X1 _15403_ ( .A1(_07298_ ), .A2(_03595_ ), .A3(_04044_ ), .ZN(_07299_ ) );
OAI21_X1 _15404_ ( .A(_03595_ ), .B1(_07298_ ), .B2(_04044_ ), .ZN(_07300_ ) );
AND3_X1 _15405_ ( .A1(_07299_ ), .A2(_06501_ ), .A3(_07300_ ), .ZN(_07301_ ) );
OAI21_X1 _15406_ ( .A(_06381_ ), .B1(_07297_ ), .B2(_07301_ ), .ZN(_07302_ ) );
NAND2_X1 _15407_ ( .A1(_07302_ ), .A2(_04161_ ), .ZN(_07303_ ) );
NOR2_X1 _15408_ ( .A1(_06957_ ), .A2(_06960_ ), .ZN(_07304_ ) );
NOR2_X1 _15409_ ( .A1(_07304_ ), .A2(_03734_ ), .ZN(_07305_ ) );
AND2_X1 _15410_ ( .A1(_03731_ ), .A2(_01765_ ), .ZN(_07306_ ) );
OR3_X1 _15411_ ( .A1(_07305_ ), .A2(_03739_ ), .A3(_07306_ ), .ZN(_07307_ ) );
OAI21_X1 _15412_ ( .A(_03739_ ), .B1(_07305_ ), .B2(_07306_ ), .ZN(_07308_ ) );
AND3_X1 _15413_ ( .A1(_07307_ ), .A2(_06561_ ), .A3(_07308_ ), .ZN(_07309_ ) );
AOI22_X1 _15414_ ( .A1(_06290_ ), .A2(_06292_ ), .B1(_06667_ ), .B2(_06849_ ), .ZN(_07310_ ) );
OAI211_X1 _15415_ ( .A(_06646_ ), .B(_06293_ ), .C1(_06298_ ), .C2(_06301_ ), .ZN(_07311_ ) );
AOI21_X1 _15416_ ( .A(_06394_ ), .B1(_07310_ ), .B2(_07311_ ), .ZN(_07312_ ) );
NAND3_X1 _15417_ ( .A1(_06854_ ), .A2(_06855_ ), .A3(_06918_ ), .ZN(_07313_ ) );
NAND3_X1 _15418_ ( .A1(_06849_ ), .A2(_06425_ ), .A3(_06180_ ), .ZN(_07314_ ) );
NAND2_X1 _15419_ ( .A1(_03739_ ), .A2(_03986_ ), .ZN(_07315_ ) );
NAND3_X1 _15420_ ( .A1(_03737_ ), .A2(_02539_ ), .A3(_06367_ ), .ZN(_07316_ ) );
AND4_X1 _15421_ ( .A1(_07313_ ), .A2(_07314_ ), .A3(_07315_ ), .A4(_07316_ ), .ZN(_07317_ ) );
NOR2_X1 _15422_ ( .A1(_06156_ ), .A2(_06162_ ), .ZN(_07318_ ) );
AOI21_X1 _15423_ ( .A(_02539_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_07319_ ) );
NOR2_X1 _15424_ ( .A1(_06161_ ), .A2(_07319_ ), .ZN(_07320_ ) );
MUX2_X1 _15425_ ( .A(_07318_ ), .B(_07320_ ), .S(_07026_ ), .Z(_07321_ ) );
NAND2_X1 _15426_ ( .A1(_07321_ ), .A2(_06674_ ), .ZN(_07322_ ) );
NAND2_X1 _15427_ ( .A1(_07322_ ), .A2(_06609_ ), .ZN(_07323_ ) );
OR3_X1 _15428_ ( .A1(_06169_ ), .A2(_06395_ ), .A3(_06159_ ), .ZN(_07324_ ) );
OR3_X1 _15429_ ( .A1(_06165_ ), .A2(_06170_ ), .A3(_07026_ ), .ZN(_07325_ ) );
AOI21_X1 _15430_ ( .A(_06674_ ), .B1(_07324_ ), .B2(_07325_ ), .ZN(_07326_ ) );
OAI221_X1 _15431_ ( .A(_06778_ ), .B1(_06363_ ), .B2(_06609_ ), .C1(_07323_ ), .C2(_07326_ ), .ZN(_07327_ ) );
OAI21_X1 _15432_ ( .A(_06486_ ), .B1(_03737_ ), .B2(_02539_ ), .ZN(_07328_ ) );
NAND3_X1 _15433_ ( .A1(_07317_ ), .A2(_07327_ ), .A3(_07328_ ), .ZN(_07329_ ) );
OR3_X2 _15434_ ( .A1(_07309_ ), .A2(_07312_ ), .A3(_07329_ ), .ZN(_07330_ ) );
AOI21_X1 _15435_ ( .A(_07303_ ), .B1(_07330_ ), .B2(_07291_ ), .ZN(_07331_ ) );
OAI21_X1 _15436_ ( .A(_07012_ ), .B1(_04157_ ), .B2(_06729_ ), .ZN(_07332_ ) );
OAI21_X1 _15437_ ( .A(_07296_ ), .B1(_07331_ ), .B2(_07332_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
OR2_X1 _15438_ ( .A1(_04749_ ), .A2(_05891_ ), .ZN(_07333_ ) );
AOI21_X1 _15439_ ( .A(_06386_ ), .B1(_03644_ ), .B2(_03991_ ), .ZN(_07334_ ) );
OAI21_X1 _15440_ ( .A(_07334_ ), .B1(_03644_ ), .B2(_03991_ ), .ZN(_07335_ ) );
AOI22_X1 _15441_ ( .A1(_04751_ ), .A2(_06116_ ), .B1(\ID_EX_imm [1] ), .B2(_06382_ ), .ZN(_07336_ ) );
AOI21_X1 _15442_ ( .A(_06573_ ), .B1(_07335_ ), .B2(_07336_ ), .ZN(_07337_ ) );
OR2_X1 _15443_ ( .A1(_07337_ ), .A2(_01650_ ), .ZN(_07338_ ) );
AND3_X1 _15444_ ( .A1(_07253_ ), .A2(_06296_ ), .A3(_06789_ ), .ZN(_07339_ ) );
OR3_X1 _15445_ ( .A1(_06651_ ), .A2(_06322_ ), .A3(_06656_ ), .ZN(_07340_ ) );
NOR3_X1 _15446_ ( .A1(_07048_ ), .A2(_06708_ ), .A3(_07049_ ), .ZN(_07341_ ) );
OAI21_X1 _15447_ ( .A(_07026_ ), .B1(_06312_ ), .B2(_06319_ ), .ZN(_07342_ ) );
OAI211_X1 _15448_ ( .A(_07342_ ), .B(_06317_ ), .C1(_07247_ ), .C2(_07026_ ), .ZN(_07343_ ) );
NAND3_X1 _15449_ ( .A1(_07184_ ), .A2(_07185_ ), .A3(_06618_ ), .ZN(_07344_ ) );
AOI21_X1 _15450_ ( .A(_06345_ ), .B1(_07343_ ), .B2(_07344_ ), .ZN(_07345_ ) );
OAI21_X1 _15451_ ( .A(_06178_ ), .B1(_07341_ ), .B2(_07345_ ), .ZN(_07346_ ) );
NAND2_X1 _15452_ ( .A1(_07340_ ), .A2(_07346_ ), .ZN(_07347_ ) );
OAI21_X1 _15453_ ( .A(_06248_ ), .B1(_07339_ ), .B2(_07347_ ), .ZN(_07348_ ) );
NAND2_X1 _15454_ ( .A1(_07347_ ), .A2(_06818_ ), .ZN(_07349_ ) );
NAND4_X1 _15455_ ( .A1(_06320_ ), .A2(_06667_ ), .A3(_06669_ ), .A4(_06674_ ), .ZN(_07350_ ) );
OAI211_X1 _15456_ ( .A(_07348_ ), .B(_07349_ ), .C1(_06305_ ), .C2(_07350_ ), .ZN(_07351_ ) );
AOI21_X1 _15457_ ( .A(_06198_ ), .B1(_03926_ ), .B2(_03928_ ), .ZN(_07352_ ) );
NOR3_X1 _15458_ ( .A1(_06199_ ), .A2(_07352_ ), .A3(_06659_ ), .ZN(_07353_ ) );
AOI22_X1 _15459_ ( .A1(_03928_ ), .A2(_06486_ ), .B1(_03925_ ), .B2(_07034_ ), .ZN(_07354_ ) );
NAND3_X1 _15460_ ( .A1(_03926_ ), .A2(_03928_ ), .A3(_06567_ ), .ZN(_07355_ ) );
NAND2_X1 _15461_ ( .A1(_07354_ ), .A2(_07355_ ), .ZN(_07356_ ) );
OR3_X1 _15462_ ( .A1(_07351_ ), .A2(_07353_ ), .A3(_07356_ ), .ZN(_07357_ ) );
AOI21_X1 _15463_ ( .A(_07338_ ), .B1(_07357_ ), .B2(_07291_ ), .ZN(_07358_ ) );
OAI21_X1 _15464_ ( .A(_07012_ ), .B1(_01655_ ), .B2(\ID_EX_pc [1] ), .ZN(_07359_ ) );
OAI21_X1 _15465_ ( .A(_07333_ ), .B1(_07358_ ), .B2(_07359_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
NAND3_X1 _15466_ ( .A1(_03722_ ), .A2(_06372_ ), .A3(_03728_ ), .ZN(_07360_ ) );
NAND4_X1 _15467_ ( .A1(_02859_ ), .A2(\ID_EX_typ [4] ), .A3(\ID_EX_typ [3] ), .A4(_03982_ ), .ZN(_07361_ ) );
NAND2_X1 _15468_ ( .A1(_07360_ ), .A2(_07361_ ), .ZN(_07362_ ) );
AND2_X1 _15469_ ( .A1(_03981_ ), .A2(_07362_ ), .ZN(_07363_ ) );
NAND3_X1 _15470_ ( .A1(_04798_ ), .A2(_06128_ ), .A3(_06114_ ), .ZN(_07364_ ) );
OAI221_X1 _15471_ ( .A(_07364_ ), .B1(_03919_ ), .B2(_06383_ ), .C1(_03670_ ), .C2(_06386_ ), .ZN(_07365_ ) );
OAI21_X1 _15472_ ( .A(_06381_ ), .B1(_07363_ ), .B2(_07365_ ), .ZN(_07366_ ) );
OAI21_X1 _15473_ ( .A(_03983_ ), .B1(_06271_ ), .B2(_04029_ ), .ZN(_07367_ ) );
AOI21_X1 _15474_ ( .A(_07367_ ), .B1(_03977_ ), .B2(_03979_ ), .ZN(_07368_ ) );
AND3_X1 _15475_ ( .A1(_03973_ ), .A2(_03976_ ), .A3(_07368_ ), .ZN(_07369_ ) );
NAND4_X1 _15476_ ( .A1(_06278_ ), .A2(_03889_ ), .A3(_06253_ ), .A4(_06287_ ), .ZN(_07370_ ) );
AND2_X1 _15477_ ( .A1(_06700_ ), .A2(_06442_ ), .ZN(_07371_ ) );
AND2_X1 _15478_ ( .A1(_06147_ ), .A2(_03646_ ), .ZN(_07372_ ) );
OAI21_X1 _15479_ ( .A(_06145_ ), .B1(_07372_ ), .B2(_06432_ ), .ZN(_07373_ ) );
OAI211_X1 _15480_ ( .A(_07373_ ), .B(_03908_ ), .C1(_06150_ ), .C2(_07275_ ), .ZN(_07374_ ) );
OAI21_X1 _15481_ ( .A(_03909_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07375_ ) );
AND3_X1 _15482_ ( .A1(_07374_ ), .A2(_06175_ ), .A3(_07375_ ), .ZN(_07376_ ) );
AOI211_X1 _15483_ ( .A(_06442_ ), .B(_07376_ ), .C1(_07088_ ), .C2(_03911_ ), .ZN(_07377_ ) );
NOR2_X1 _15484_ ( .A1(_07371_ ), .A2(_07377_ ), .ZN(_07378_ ) );
AOI21_X1 _15485_ ( .A(_06393_ ), .B1(_07370_ ), .B2(_07378_ ), .ZN(_07379_ ) );
NOR2_X1 _15486_ ( .A1(_07378_ ), .A2(_06887_ ), .ZN(_07380_ ) );
AND4_X1 _15487_ ( .A1(_06177_ ), .A2(_06707_ ), .A3(_06546_ ), .A4(_04070_ ), .ZN(_07381_ ) );
OR4_X1 _15488_ ( .A1(_07369_ ), .A2(_07379_ ), .A3(_07380_ ), .A4(_07381_ ), .ZN(_07382_ ) );
NOR3_X1 _15489_ ( .A1(_07372_ ), .A2(_06198_ ), .A3(_06634_ ), .ZN(_07383_ ) );
OAI21_X1 _15490_ ( .A(_03986_ ), .B1(_06429_ ), .B2(_03922_ ), .ZN(_07384_ ) );
NAND3_X1 _15491_ ( .A1(_06396_ ), .A2(_03645_ ), .A3(_03723_ ), .ZN(_07385_ ) );
OAI211_X1 _15492_ ( .A(_07384_ ), .B(_07385_ ), .C1(_06135_ ), .C2(_07372_ ), .ZN(_07386_ ) );
NOR3_X1 _15493_ ( .A1(_07382_ ), .A2(_07383_ ), .A3(_07386_ ), .ZN(_07387_ ) );
OAI21_X1 _15494_ ( .A(_07366_ ), .B1(_07387_ ), .B2(_06375_ ), .ZN(_07388_ ) );
MUX2_X1 _15495_ ( .A(\ID_EX_pc [0] ), .B(_07388_ ), .S(_02840_ ), .Z(_07389_ ) );
MUX2_X1 _15496_ ( .A(_06041_ ), .B(_07389_ ), .S(_05867_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
OR3_X1 _15497_ ( .A1(_04468_ ), .A2(_05861_ ), .A3(_04470_ ), .ZN(_07390_ ) );
NOR2_X1 _15498_ ( .A1(_04476_ ), .A2(_06118_ ), .ZN(_07391_ ) );
OAI21_X1 _15499_ ( .A(_06125_ ), .B1(_06905_ ), .B2(_06907_ ), .ZN(_07392_ ) );
AOI21_X1 _15500_ ( .A(_07392_ ), .B1(_06907_ ), .B2(_06905_ ), .ZN(_07393_ ) );
AND3_X1 _15501_ ( .A1(_06127_ ), .A2(\ID_EX_imm [28] ), .A3(_06128_ ), .ZN(_07394_ ) );
NOR3_X1 _15502_ ( .A1(_07391_ ), .A2(_07393_ ), .A3(_07394_ ), .ZN(_07395_ ) );
OAI21_X1 _15503_ ( .A(_01654_ ), .B1(_07395_ ), .B2(_06133_ ), .ZN(_07396_ ) );
OR3_X1 _15504_ ( .A1(_06889_ ), .A2(_06178_ ), .A3(_06890_ ), .ZN(_07397_ ) );
OAI21_X1 _15505_ ( .A(_07026_ ), .B1(_06405_ ), .B2(_06410_ ), .ZN(_07398_ ) );
OAI21_X1 _15506_ ( .A(_06395_ ), .B1(_06402_ ), .B2(_06406_ ), .ZN(_07399_ ) );
AND3_X1 _15507_ ( .A1(_07398_ ), .A2(_07399_ ), .A3(_06325_ ), .ZN(_07400_ ) );
MUX2_X1 _15508_ ( .A(_06928_ ), .B(_06932_ ), .S(_07026_ ), .Z(_07401_ ) );
AOI211_X1 _15509_ ( .A(_06364_ ), .B(_07400_ ), .C1(_06674_ ), .C2(_07401_ ), .ZN(_07402_ ) );
NOR3_X1 _15510_ ( .A1(_06454_ ), .A2(_06460_ ), .A3(_06668_ ), .ZN(_07403_ ) );
OAI21_X1 _15511_ ( .A(_06530_ ), .B1(_07402_ ), .B2(_07403_ ), .ZN(_07404_ ) );
NAND3_X1 _15512_ ( .A1(_07397_ ), .A2(_07404_ ), .A3(_04070_ ), .ZN(_07405_ ) );
NAND3_X1 _15513_ ( .A1(_06421_ ), .A2(_06668_ ), .A3(_06674_ ), .ZN(_07406_ ) );
OR3_X1 _15514_ ( .A1(_07406_ ), .A2(_06600_ ), .A3(_06887_ ), .ZN(_07407_ ) );
AND3_X1 _15515_ ( .A1(_06288_ ), .A2(_06299_ ), .A3(_06397_ ), .ZN(_07408_ ) );
OAI21_X1 _15516_ ( .A(_07408_ ), .B1(_06290_ ), .B2(_06293_ ), .ZN(_07409_ ) );
INV_X1 _15517_ ( .A(_07409_ ), .ZN(_07410_ ) );
NOR2_X1 _15518_ ( .A1(_07406_ ), .A2(_06443_ ), .ZN(_07411_ ) );
NOR4_X1 _15519_ ( .A1(_07410_ ), .A2(_06549_ ), .A3(_06940_ ), .A4(_07411_ ), .ZN(_07412_ ) );
OAI211_X1 _15520_ ( .A(_07405_ ), .B(_07407_ ), .C1(_07412_ ), .C2(_06394_ ), .ZN(_07413_ ) );
OAI21_X1 _15521_ ( .A(_06245_ ), .B1(_07304_ ), .B2(_03734_ ), .ZN(_07414_ ) );
AOI21_X1 _15522_ ( .A(_07414_ ), .B1(_03734_ ), .B2(_07304_ ), .ZN(_07415_ ) );
NAND2_X1 _15523_ ( .A1(_03733_ ), .A2(_06567_ ), .ZN(_07416_ ) );
NAND3_X1 _15524_ ( .A1(_03731_ ), .A2(_01765_ ), .A3(_07034_ ), .ZN(_07417_ ) );
OAI21_X1 _15525_ ( .A(_06486_ ), .B1(_03731_ ), .B2(_01765_ ), .ZN(_07418_ ) );
NAND3_X1 _15526_ ( .A1(_07416_ ), .A2(_07417_ ), .A3(_07418_ ), .ZN(_07419_ ) );
OR3_X1 _15527_ ( .A1(_07413_ ), .A2(_07415_ ), .A3(_07419_ ), .ZN(_07420_ ) );
AOI21_X1 _15528_ ( .A(_07396_ ), .B1(_07420_ ), .B2(_07291_ ), .ZN(_07421_ ) );
OAI21_X1 _15529_ ( .A(_07012_ ), .B1(_04473_ ), .B2(_06729_ ), .ZN(_07422_ ) );
OAI21_X1 _15530_ ( .A(_07390_ ), .B1(_07421_ ), .B2(_07422_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND3_X1 _15531_ ( .A1(_04774_ ), .A2(_05879_ ), .A3(_04776_ ), .ZN(_07423_ ) );
OAI22_X1 _15532_ ( .A1(_04784_ ), .A2(_06118_ ), .B1(_02485_ ), .B2(_06383_ ), .ZN(_07424_ ) );
OAI21_X1 _15533_ ( .A(_03480_ ), .B1(_06903_ ), .B2(_04067_ ), .ZN(_07425_ ) );
NAND3_X1 _15534_ ( .A1(_07425_ ), .A2(_03478_ ), .A3(_04033_ ), .ZN(_07426_ ) );
AND2_X1 _15535_ ( .A1(_07426_ ), .A2(_03526_ ), .ZN(_07427_ ) );
OR3_X1 _15536_ ( .A1(_07427_ ), .A2(_03503_ ), .A3(_04037_ ), .ZN(_07428_ ) );
OAI21_X1 _15537_ ( .A(_03503_ ), .B1(_07427_ ), .B2(_04037_ ), .ZN(_07429_ ) );
AND3_X1 _15538_ ( .A1(_07428_ ), .A2(_06501_ ), .A3(_07429_ ), .ZN(_07430_ ) );
OAI21_X1 _15539_ ( .A(_06381_ ), .B1(_07424_ ), .B2(_07430_ ), .ZN(_07431_ ) );
NAND2_X1 _15540_ ( .A1(_07431_ ), .A2(_04161_ ), .ZN(_07432_ ) );
NOR2_X1 _15541_ ( .A1(_06545_ ), .A2(_06345_ ), .ZN(_07433_ ) );
AND3_X1 _15542_ ( .A1(_07433_ ), .A2(_06178_ ), .A3(_06180_ ), .ZN(_07434_ ) );
INV_X1 _15543_ ( .A(_06549_ ), .ZN(_07435_ ) );
INV_X1 _15544_ ( .A(_06940_ ), .ZN(_07436_ ) );
OAI211_X1 _15545_ ( .A(_06288_ ), .B(_06550_ ), .C1(_06289_ ), .C2(_06293_ ), .ZN(_07437_ ) );
NAND2_X1 _15546_ ( .A1(_07433_ ), .A2(_06425_ ), .ZN(_07438_ ) );
NAND4_X1 _15547_ ( .A1(_07435_ ), .A2(_07436_ ), .A3(_07437_ ), .A4(_07438_ ), .ZN(_07439_ ) );
AOI21_X1 _15548_ ( .A(_07434_ ), .B1(_07439_ ), .B2(_06248_ ), .ZN(_07440_ ) );
NAND3_X1 _15549_ ( .A1(_06994_ ), .A2(_06918_ ), .A3(_06995_ ), .ZN(_07441_ ) );
AND2_X1 _15550_ ( .A1(_06528_ ), .A2(_06842_ ), .ZN(_07442_ ) );
NAND2_X1 _15551_ ( .A1(_07318_ ), .A2(_06151_ ), .ZN(_07443_ ) );
OR3_X1 _15552_ ( .A1(_06169_ ), .A2(_06159_ ), .A3(_06150_ ), .ZN(_07444_ ) );
NAND2_X1 _15553_ ( .A1(_07443_ ), .A2(_07444_ ), .ZN(_07445_ ) );
OR3_X1 _15554_ ( .A1(_06165_ ), .A2(_06158_ ), .A3(_06170_ ), .ZN(_07446_ ) );
OR3_X1 _15555_ ( .A1(_06347_ ), .A2(_06166_ ), .A3(_06146_ ), .ZN(_07447_ ) );
NAND2_X1 _15556_ ( .A1(_07446_ ), .A2(_07447_ ), .ZN(_07448_ ) );
MUX2_X1 _15557_ ( .A(_07445_ ), .B(_07448_ ), .S(_06607_ ), .Z(_07449_ ) );
OAI21_X1 _15558_ ( .A(_06778_ ), .B1(_07449_ ), .B2(_06842_ ), .ZN(_07450_ ) );
OAI211_X1 _15559_ ( .A(_07440_ ), .B(_07441_ ), .C1(_07442_ ), .C2(_07450_ ), .ZN(_07451_ ) );
AOI21_X1 _15560_ ( .A(_03759_ ), .B1(_06954_ ), .B2(_06956_ ), .ZN(_07452_ ) );
OR3_X1 _15561_ ( .A1(_07452_ ), .A2(_03766_ ), .A3(_03756_ ), .ZN(_07453_ ) );
OAI21_X1 _15562_ ( .A(_03766_ ), .B1(_07452_ ), .B2(_03756_ ), .ZN(_07454_ ) );
AND3_X1 _15563_ ( .A1(_07453_ ), .A2(_06561_ ), .A3(_07454_ ), .ZN(_07455_ ) );
AOI22_X1 _15564_ ( .A1(_06958_ ), .A2(_06486_ ), .B1(_03764_ ), .B2(_06367_ ), .ZN(_07456_ ) );
OAI21_X1 _15565_ ( .A(_07456_ ), .B1(_03767_ ), .B2(_03987_ ), .ZN(_07457_ ) );
OR3_X1 _15566_ ( .A1(_07451_ ), .A2(_07455_ ), .A3(_07457_ ), .ZN(_07458_ ) );
AOI21_X1 _15567_ ( .A(_07432_ ), .B1(_07458_ ), .B2(_07291_ ), .ZN(_07459_ ) );
OAI21_X1 _15568_ ( .A(_05867_ ), .B1(_04779_ ), .B2(_06729_ ), .ZN(_07460_ ) );
OAI21_X1 _15569_ ( .A(_07423_ ), .B1(_07459_ ), .B2(_07460_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
OR2_X1 _15570_ ( .A1(_04824_ ), .A2(_05891_ ), .ZN(_07461_ ) );
OAI22_X1 _15571_ ( .A1(_04827_ ), .A2(_06118_ ), .B1(_02511_ ), .B2(_06383_ ), .ZN(_07462_ ) );
NOR2_X1 _15572_ ( .A1(_07426_ ), .A2(_03526_ ), .ZN(_07463_ ) );
NOR3_X1 _15573_ ( .A1(_07427_ ), .A2(_07463_ ), .A3(_06387_ ), .ZN(_07464_ ) );
OAI21_X1 _15574_ ( .A(_06381_ ), .B1(_07462_ ), .B2(_07464_ ), .ZN(_07465_ ) );
NAND2_X1 _15575_ ( .A1(_07465_ ), .A2(_04161_ ), .ZN(_07466_ ) );
AND2_X1 _15576_ ( .A1(_07032_ ), .A2(_06322_ ), .ZN(_07467_ ) );
OR3_X1 _15577_ ( .A1(_06549_ ), .A2(_06940_ ), .A3(_07467_ ), .ZN(_07468_ ) );
NOR3_X1 _15578_ ( .A1(_06581_ ), .A2(_06583_ ), .A3(_06584_ ), .ZN(_07469_ ) );
OAI21_X1 _15579_ ( .A(_06248_ ), .B1(_07468_ ), .B2(_07469_ ), .ZN(_07470_ ) );
NAND3_X1 _15580_ ( .A1(_07032_ ), .A2(_06630_ ), .A3(_06818_ ), .ZN(_07471_ ) );
AOI22_X1 _15581_ ( .A1(_03758_ ), .A2(_06567_ ), .B1(_03756_ ), .B2(_07034_ ), .ZN(_07472_ ) );
NAND3_X1 _15582_ ( .A1(_07470_ ), .A2(_07471_ ), .A3(_07472_ ), .ZN(_07473_ ) );
AND3_X1 _15583_ ( .A1(_06954_ ), .A2(_03759_ ), .A3(_06956_ ), .ZN(_07474_ ) );
NOR3_X1 _15584_ ( .A1(_07474_ ), .A2(_07452_ ), .A3(_06659_ ), .ZN(_07475_ ) );
NAND3_X1 _15585_ ( .A1(_07038_ ), .A2(_06918_ ), .A3(_07039_ ), .ZN(_07476_ ) );
MUX2_X1 _15586_ ( .A(_06931_ ), .B(_06924_ ), .S(_06607_ ), .Z(_07477_ ) );
OAI21_X1 _15587_ ( .A(_06778_ ), .B1(_07477_ ), .B2(_06842_ ), .ZN(_07478_ ) );
AND2_X1 _15588_ ( .A1(_06619_ ), .A2(_06842_ ), .ZN(_07479_ ) );
OAI221_X1 _15589_ ( .A(_07476_ ), .B1(_03757_ ), .B2(_06565_ ), .C1(_07478_ ), .C2(_07479_ ), .ZN(_07480_ ) );
OR3_X1 _15590_ ( .A1(_07473_ ), .A2(_07475_ ), .A3(_07480_ ), .ZN(_07481_ ) );
AOI21_X1 _15591_ ( .A(_07466_ ), .B1(_07481_ ), .B2(_07291_ ), .ZN(_07482_ ) );
NAND2_X1 _15592_ ( .A1(_04825_ ), .A2(_06685_ ), .ZN(_07483_ ) );
NAND2_X1 _15593_ ( .A1(_07483_ ), .A2(_05888_ ), .ZN(_07484_ ) );
OAI21_X1 _15594_ ( .A(_07461_ ), .B1(_07482_ ), .B2(_07484_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
OAI21_X1 _15595_ ( .A(_05916_ ), .B1(_04841_ ), .B2(_04847_ ), .ZN(_07485_ ) );
OAI22_X1 _15596_ ( .A1(_04859_ ), .A2(_06117_ ), .B1(_02457_ ), .B2(_06383_ ), .ZN(_07486_ ) );
NOR2_X1 _15597_ ( .A1(_06903_ ), .A2(_04067_ ), .ZN(_07487_ ) );
INV_X1 _15598_ ( .A(_03451_ ), .ZN(_07488_ ) );
NOR2_X1 _15599_ ( .A1(_07487_ ), .A2(_07488_ ), .ZN(_07489_ ) );
NOR2_X1 _15600_ ( .A1(_03450_ ), .A2(_06168_ ), .ZN(_07490_ ) );
OAI21_X1 _15601_ ( .A(_03479_ ), .B1(_07489_ ), .B2(_07490_ ), .ZN(_07491_ ) );
NOR3_X1 _15602_ ( .A1(_07489_ ), .A2(_03479_ ), .A3(_07490_ ), .ZN(_07492_ ) );
NOR2_X1 _15603_ ( .A1(_07492_ ), .A2(_06387_ ), .ZN(_07493_ ) );
AOI21_X1 _15604_ ( .A(_07486_ ), .B1(_07491_ ), .B2(_07493_ ), .ZN(_07494_ ) );
OAI21_X1 _15605_ ( .A(_01654_ ), .B1(_07494_ ), .B2(_06133_ ), .ZN(_07495_ ) );
AND3_X1 _15606_ ( .A1(_06649_ ), .A2(_06650_ ), .A3(_06708_ ), .ZN(_07496_ ) );
AND2_X1 _15607_ ( .A1(_07496_ ), .A2(_06425_ ), .ZN(_07497_ ) );
OR3_X1 _15608_ ( .A1(_06549_ ), .A2(_06940_ ), .A3(_07497_ ), .ZN(_07498_ ) );
NAND3_X1 _15609_ ( .A1(_06582_ ), .A2(_06296_ ), .A3(_06299_ ), .ZN(_07499_ ) );
NOR2_X1 _15610_ ( .A1(_07499_ ), .A2(_06581_ ), .ZN(_07500_ ) );
OAI21_X1 _15611_ ( .A(_06249_ ), .B1(_07498_ ), .B2(_07500_ ), .ZN(_07501_ ) );
OAI21_X1 _15612_ ( .A(_03772_ ), .B1(_06946_ ), .B2(_06953_ ), .ZN(_07502_ ) );
INV_X1 _15613_ ( .A(_06955_ ), .ZN(_07503_ ) );
NAND2_X1 _15614_ ( .A1(_07502_ ), .A2(_07503_ ), .ZN(_07504_ ) );
AOI21_X1 _15615_ ( .A(_06659_ ), .B1(_07504_ ), .B2(_03778_ ), .ZN(_07505_ ) );
OAI21_X1 _15616_ ( .A(_07505_ ), .B1(_03778_ ), .B2(_07504_ ), .ZN(_07506_ ) );
NAND2_X1 _15617_ ( .A1(_06665_ ), .A2(_06842_ ), .ZN(_07507_ ) );
AOI21_X1 _15618_ ( .A(_06607_ ), .B1(_07324_ ), .B2(_07325_ ), .ZN(_07508_ ) );
AOI21_X1 _15619_ ( .A(_06620_ ), .B1(_06348_ ), .B2(_06353_ ), .ZN(_07509_ ) );
OR3_X1 _15620_ ( .A1(_07508_ ), .A2(_07509_ ), .A3(_06765_ ), .ZN(_07510_ ) );
NAND3_X1 _15621_ ( .A1(_07507_ ), .A2(_07510_ ), .A3(_06778_ ), .ZN(_07511_ ) );
NAND3_X1 _15622_ ( .A1(_07496_ ), .A2(_06630_ ), .A3(_06818_ ), .ZN(_07512_ ) );
NAND2_X1 _15623_ ( .A1(_07511_ ), .A2(_07512_ ), .ZN(_07513_ ) );
AND2_X1 _15624_ ( .A1(_07066_ ), .A2(_06918_ ), .ZN(_07514_ ) );
AOI22_X1 _15625_ ( .A1(_03778_ ), .A2(_06368_ ), .B1(_03776_ ), .B2(_06367_ ), .ZN(_07515_ ) );
OAI21_X1 _15626_ ( .A(_07515_ ), .B1(_03777_ ), .B2(_06565_ ), .ZN(_07516_ ) );
NOR3_X1 _15627_ ( .A1(_07513_ ), .A2(_07514_ ), .A3(_07516_ ), .ZN(_07517_ ) );
NAND3_X1 _15628_ ( .A1(_07501_ ), .A2(_07506_ ), .A3(_07517_ ), .ZN(_07518_ ) );
AOI21_X1 _15629_ ( .A(_07495_ ), .B1(_07518_ ), .B2(_07291_ ), .ZN(_07519_ ) );
OAI21_X1 _15630_ ( .A(_05867_ ), .B1(_04855_ ), .B2(_06391_ ), .ZN(_07520_ ) );
OAI21_X1 _15631_ ( .A(_07485_ ), .B1(_07519_ ), .B2(_07520_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
INV_X1 _15632_ ( .A(_06077_ ), .ZN(_07521_ ) );
OAI22_X1 _15633_ ( .A1(_04884_ ), .A2(_06118_ ), .B1(_02433_ ), .B2(_06383_ ), .ZN(_07522_ ) );
OAI21_X1 _15634_ ( .A(_06125_ ), .B1(_07487_ ), .B2(_07488_ ), .ZN(_07523_ ) );
AOI21_X1 _15635_ ( .A(_07523_ ), .B1(_07488_ ), .B2(_07487_ ), .ZN(_07524_ ) );
OAI21_X1 _15636_ ( .A(_06381_ ), .B1(_07522_ ), .B2(_07524_ ), .ZN(_07525_ ) );
NAND2_X1 _15637_ ( .A1(_07525_ ), .A2(_04161_ ), .ZN(_07526_ ) );
AND4_X1 _15638_ ( .A1(_07083_ ), .A2(_06278_ ), .A3(_06287_ ), .A4(_06293_ ), .ZN(_07527_ ) );
AND2_X1 _15639_ ( .A1(_06699_ ), .A2(_06668_ ), .ZN(_07528_ ) );
AND2_X1 _15640_ ( .A1(_07528_ ), .A2(_06530_ ), .ZN(_07529_ ) );
OR2_X1 _15641_ ( .A1(_07527_ ), .A2(_07529_ ), .ZN(_07530_ ) );
OAI21_X1 _15642_ ( .A(_06249_ ), .B1(_06549_ ), .B2(_07530_ ), .ZN(_07531_ ) );
OR3_X1 _15643_ ( .A1(_06946_ ), .A2(_03772_ ), .A3(_06953_ ), .ZN(_07532_ ) );
NAND3_X1 _15644_ ( .A1(_07532_ ), .A2(_06561_ ), .A3(_07502_ ), .ZN(_07533_ ) );
OR3_X1 _15645_ ( .A1(_03771_ ), .A2(_06168_ ), .A3(_06488_ ), .ZN(_07534_ ) );
AOI21_X1 _15646_ ( .A(_06620_ ), .B1(_06456_ ), .B2(_06459_ ), .ZN(_07535_ ) );
AOI21_X1 _15647_ ( .A(_06618_ ), .B1(_07398_ ), .B2(_07399_ ), .ZN(_07536_ ) );
OAI21_X1 _15648_ ( .A(_06668_ ), .B1(_07535_ ), .B2(_07536_ ), .ZN(_07537_ ) );
NAND2_X1 _15649_ ( .A1(_07537_ ), .A2(_06777_ ), .ZN(_07538_ ) );
AOI21_X1 _15650_ ( .A(_06609_ ), .B1(_06711_ ), .B2(_06712_ ), .ZN(_07539_ ) );
NOR2_X1 _15651_ ( .A1(_07538_ ), .A2(_07539_ ), .ZN(_07540_ ) );
AOI21_X1 _15652_ ( .A(_07540_ ), .B1(_07529_ ), .B2(_06181_ ), .ZN(_07541_ ) );
AOI21_X1 _15653_ ( .A(_06565_ ), .B1(_03771_ ), .B2(_06168_ ), .ZN(_07542_ ) );
AOI21_X1 _15654_ ( .A(_07542_ ), .B1(_03772_ ), .B2(_06567_ ), .ZN(_07543_ ) );
NAND3_X1 _15655_ ( .A1(_07095_ ), .A2(_06918_ ), .A3(_07096_ ), .ZN(_07544_ ) );
AND4_X1 _15656_ ( .A1(_07534_ ), .A2(_07541_ ), .A3(_07543_ ), .A4(_07544_ ), .ZN(_07545_ ) );
NAND3_X1 _15657_ ( .A1(_07531_ ), .A2(_07533_ ), .A3(_07545_ ), .ZN(_07546_ ) );
AOI21_X1 _15658_ ( .A(_07526_ ), .B1(_07546_ ), .B2(_07291_ ), .ZN(_07547_ ) );
OAI21_X1 _15659_ ( .A(_05867_ ), .B1(_04882_ ), .B2(_06391_ ), .ZN(_07548_ ) );
OAI21_X1 _15660_ ( .A(_07521_ ), .B1(_07547_ ), .B2(_07548_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
OAI21_X1 _15661_ ( .A(_05916_ ), .B1(_04898_ ), .B2(_04904_ ), .ZN(_07549_ ) );
AND3_X1 _15662_ ( .A1(_06121_ ), .A2(_03085_ ), .A3(_03109_ ), .ZN(_07550_ ) );
OR2_X1 _15663_ ( .A1(_07550_ ), .A2(_04064_ ), .ZN(_07551_ ) );
AND2_X1 _15664_ ( .A1(_07551_ ), .A2(_03034_ ), .ZN(_07552_ ) );
OR3_X1 _15665_ ( .A1(_07552_ ), .A2(_03059_ ), .A3(_04058_ ), .ZN(_07553_ ) );
OAI21_X1 _15666_ ( .A(_03059_ ), .B1(_07552_ ), .B2(_04058_ ), .ZN(_07554_ ) );
NAND3_X1 _15667_ ( .A1(_07553_ ), .A2(_06501_ ), .A3(_07554_ ), .ZN(_07555_ ) );
AOI22_X1 _15668_ ( .A1(_04895_ ), .A2(_06116_ ), .B1(\ID_EX_imm [23] ), .B2(_06382_ ), .ZN(_07556_ ) );
AOI21_X1 _15669_ ( .A(_06573_ ), .B1(_07555_ ), .B2(_07556_ ), .ZN(_07557_ ) );
OR2_X1 _15670_ ( .A1(_07557_ ), .A2(_01650_ ), .ZN(_07558_ ) );
NOR2_X1 _15671_ ( .A1(_06549_ ), .A2(_06940_ ), .ZN(_07559_ ) );
INV_X1 _15672_ ( .A(_07559_ ), .ZN(_07560_ ) );
AND2_X1 _15673_ ( .A1(_07140_ ), .A2(_06530_ ), .ZN(_07561_ ) );
OAI21_X1 _15674_ ( .A(_06248_ ), .B1(_07560_ ), .B2(_07561_ ), .ZN(_07562_ ) );
NAND3_X1 _15675_ ( .A1(_07140_ ), .A2(_06630_ ), .A3(_06181_ ), .ZN(_07563_ ) );
NAND2_X1 _15676_ ( .A1(_07562_ ), .A2(_07563_ ), .ZN(_07564_ ) );
NAND3_X1 _15677_ ( .A1(_06774_ ), .A2(_06775_ ), .A3(_06765_ ), .ZN(_07565_ ) );
NAND2_X1 _15678_ ( .A1(_07448_ ), .A2(_06422_ ), .ZN(_07566_ ) );
NAND3_X1 _15679_ ( .A1(_06522_ ), .A2(_06523_ ), .A3(_06154_ ), .ZN(_07567_ ) );
NAND2_X1 _15680_ ( .A1(_07566_ ), .A2(_07567_ ), .ZN(_07568_ ) );
OAI211_X1 _15681_ ( .A(_06530_ ), .B(_07565_ ), .C1(_07568_ ), .C2(_06842_ ), .ZN(_07569_ ) );
OAI211_X1 _15682_ ( .A(_06600_ ), .B(_06669_ ), .C1(_06771_ ), .C2(_06772_ ), .ZN(_07570_ ) );
AOI21_X1 _15683_ ( .A(_06305_ ), .B1(_07569_ ), .B2(_07570_ ), .ZN(_07571_ ) );
NOR3_X1 _15684_ ( .A1(_03788_ ), .A2(_03789_ ), .A3(_03987_ ), .ZN(_07572_ ) );
NOR3_X1 _15685_ ( .A1(_03787_ ), .A2(_03058_ ), .A3(_06488_ ), .ZN(_07573_ ) );
NOR2_X1 _15686_ ( .A1(_03789_ ), .A2(_06135_ ), .ZN(_07574_ ) );
OR2_X1 _15687_ ( .A1(_07573_ ), .A2(_07574_ ), .ZN(_07575_ ) );
NOR4_X1 _15688_ ( .A1(_07564_ ), .A2(_07571_ ), .A3(_07572_ ), .A4(_07575_ ), .ZN(_07576_ ) );
OR3_X1 _15689_ ( .A1(_06238_ ), .A2(_06239_ ), .A3(_06241_ ), .ZN(_07577_ ) );
INV_X1 _15690_ ( .A(_06949_ ), .ZN(_07578_ ) );
AOI21_X1 _15691_ ( .A(_03784_ ), .B1(_07577_ ), .B2(_07578_ ), .ZN(_07579_ ) );
NOR2_X1 _15692_ ( .A1(_03782_ ), .A2(_03033_ ), .ZN(_07580_ ) );
NOR3_X1 _15693_ ( .A1(_07579_ ), .A2(_03962_ ), .A3(_07580_ ), .ZN(_07581_ ) );
OAI21_X1 _15694_ ( .A(_03962_ ), .B1(_07579_ ), .B2(_07580_ ), .ZN(_07582_ ) );
NAND2_X1 _15695_ ( .A1(_07582_ ), .A2(_06561_ ), .ZN(_07583_ ) );
OAI21_X1 _15696_ ( .A(_07576_ ), .B1(_07581_ ), .B2(_07583_ ), .ZN(_07584_ ) );
AOI21_X1 _15697_ ( .A(_07558_ ), .B1(_07584_ ), .B2(_07291_ ), .ZN(_07585_ ) );
OAI21_X1 _15698_ ( .A(_05867_ ), .B1(_04908_ ), .B2(_06391_ ), .ZN(_07586_ ) );
OAI21_X1 _15699_ ( .A(_07549_ ), .B1(_07585_ ), .B2(_07586_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _15700_ ( .A1(_04917_ ), .A2(_05879_ ), .A3(_04918_ ), .ZN(_07587_ ) );
AOI21_X1 _15701_ ( .A(_06386_ ), .B1(_07551_ ), .B2(_03034_ ), .ZN(_07588_ ) );
OAI21_X1 _15702_ ( .A(_07588_ ), .B1(_03034_ ), .B2(_07551_ ), .ZN(_07589_ ) );
AOI22_X1 _15703_ ( .A1(_04924_ ), .A2(_06116_ ), .B1(\ID_EX_imm [22] ), .B2(_06382_ ), .ZN(_07590_ ) );
AOI21_X1 _15704_ ( .A(_06132_ ), .B1(_07589_ ), .B2(_07590_ ), .ZN(_07591_ ) );
OR2_X1 _15705_ ( .A1(_07591_ ), .A2(_01650_ ), .ZN(_07592_ ) );
AND3_X1 _15706_ ( .A1(_06793_ ), .A2(_06301_ ), .A3(_06293_ ), .ZN(_07593_ ) );
AND2_X1 _15707_ ( .A1(_07154_ ), .A2(_06530_ ), .ZN(_07594_ ) );
OR3_X1 _15708_ ( .A1(_06549_ ), .A2(_07593_ ), .A3(_07594_ ), .ZN(_07595_ ) );
NAND2_X1 _15709_ ( .A1(_07595_ ), .A2(_06249_ ), .ZN(_07596_ ) );
AND3_X1 _15710_ ( .A1(_07577_ ), .A2(_03784_ ), .A3(_07578_ ), .ZN(_07597_ ) );
OR3_X1 _15711_ ( .A1(_07597_ ), .A2(_07579_ ), .A3(_06659_ ), .ZN(_07598_ ) );
NAND3_X1 _15712_ ( .A1(_07154_ ), .A2(_06630_ ), .A3(_06818_ ), .ZN(_07599_ ) );
AND3_X1 _15713_ ( .A1(_06925_ ), .A2(_06668_ ), .A3(_06926_ ), .ZN(_07600_ ) );
AND3_X1 _15714_ ( .A1(_06813_ ), .A2(_06364_ ), .A3(_06814_ ), .ZN(_07601_ ) );
OAI21_X1 _15715_ ( .A(_06667_ ), .B1(_07600_ ), .B2(_07601_ ), .ZN(_07602_ ) );
OAI21_X1 _15716_ ( .A(_06600_ ), .B1(_06811_ ), .B2(_06842_ ), .ZN(_07603_ ) );
NAND3_X1 _15717_ ( .A1(_07602_ ), .A2(_04070_ ), .A3(_07603_ ), .ZN(_07604_ ) );
NAND3_X1 _15718_ ( .A1(_03963_ ), .A2(_01793_ ), .A3(_07034_ ), .ZN(_07605_ ) );
AOI21_X1 _15719_ ( .A(_06135_ ), .B1(_03782_ ), .B2(_03033_ ), .ZN(_07606_ ) );
AOI21_X1 _15720_ ( .A(_07606_ ), .B1(_03783_ ), .B2(_06368_ ), .ZN(_07607_ ) );
AND4_X1 _15721_ ( .A1(_07599_ ), .A2(_07604_ ), .A3(_07605_ ), .A4(_07607_ ), .ZN(_07608_ ) );
NAND3_X1 _15722_ ( .A1(_07596_ ), .A2(_07598_ ), .A3(_07608_ ), .ZN(_07609_ ) );
AOI21_X1 _15723_ ( .A(_07592_ ), .B1(_07609_ ), .B2(_07291_ ), .ZN(_07610_ ) );
NAND2_X1 _15724_ ( .A1(_04921_ ), .A2(_06685_ ), .ZN(_07611_ ) );
NAND2_X1 _15725_ ( .A1(_07611_ ), .A2(_05888_ ), .ZN(_07612_ ) );
OAI21_X1 _15726_ ( .A(_07587_ ), .B1(_07610_ ), .B2(_07612_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
OR2_X1 _15727_ ( .A1(_04981_ ), .A2(_06117_ ), .ZN(_07613_ ) );
AOI21_X1 _15728_ ( .A(_04031_ ), .B1(_06909_ ), .B2(_03550_ ), .ZN(_07614_ ) );
XNOR2_X1 _15729_ ( .A(_07614_ ), .B(_03572_ ), .ZN(_07615_ ) );
AOI22_X1 _15730_ ( .A1(_07615_ ), .A2(_06125_ ), .B1(\ID_EX_imm [31] ), .B2(_06382_ ), .ZN(_07616_ ) );
AOI21_X1 _15731_ ( .A(_06132_ ), .B1(_07613_ ), .B2(_07616_ ), .ZN(_07617_ ) );
NOR2_X1 _15732_ ( .A1(_06965_ ), .A2(_03744_ ), .ZN(_07618_ ) );
AOI21_X1 _15733_ ( .A(_06634_ ), .B1(_07618_ ), .B2(_03977_ ), .ZN(_07619_ ) );
OAI21_X1 _15734_ ( .A(_07619_ ), .B1(_03977_ ), .B2(_07618_ ), .ZN(_07620_ ) );
AND2_X1 _15735_ ( .A1(_06769_ ), .A2(_06322_ ), .ZN(_07621_ ) );
OAI21_X1 _15736_ ( .A(_06247_ ), .B1(_06290_ ), .B2(_07621_ ), .ZN(_07622_ ) );
NAND3_X1 _15737_ ( .A1(_06773_ ), .A2(_06776_ ), .A3(_06918_ ), .ZN(_07623_ ) );
OAI21_X1 _15738_ ( .A(_06144_ ), .B1(_06396_ ), .B2(_04029_ ), .ZN(_07624_ ) );
MUX2_X1 _15739_ ( .A(_07320_ ), .B(_07624_ ), .S(_06146_ ), .Z(_07625_ ) );
MUX2_X1 _15740_ ( .A(_07445_ ), .B(_07625_ ), .S(_06316_ ), .Z(_07626_ ) );
MUX2_X1 _15741_ ( .A(_07568_ ), .B(_07626_ ), .S(_06546_ ), .Z(_07627_ ) );
NAND2_X1 _15742_ ( .A1(_07627_ ), .A2(_06777_ ), .ZN(_07628_ ) );
AND3_X1 _15743_ ( .A1(_06769_ ), .A2(_06177_ ), .A3(_06180_ ), .ZN(_07629_ ) );
AND3_X1 _15744_ ( .A1(_06271_ ), .A2(_02571_ ), .A3(_03723_ ), .ZN(_07630_ ) );
OAI21_X1 _15745_ ( .A(_04075_ ), .B1(_06271_ ), .B2(_02571_ ), .ZN(_07631_ ) );
OAI21_X1 _15746_ ( .A(_07631_ ), .B1(_03977_ ), .B2(_03987_ ), .ZN(_07632_ ) );
NOR3_X1 _15747_ ( .A1(_07629_ ), .A2(_07630_ ), .A3(_07632_ ), .ZN(_07633_ ) );
AND4_X1 _15748_ ( .A1(_07622_ ), .A2(_07623_ ), .A3(_07628_ ), .A4(_07633_ ), .ZN(_07634_ ) );
AOI21_X1 _15749_ ( .A(_06375_ ), .B1(_07620_ ), .B2(_07634_ ), .ZN(_07635_ ) );
OAI21_X1 _15750_ ( .A(_01654_ ), .B1(_07617_ ), .B2(_07635_ ), .ZN(_07636_ ) );
OAI21_X1 _15751_ ( .A(_07636_ ), .B1(_04161_ ), .B2(_04986_ ), .ZN(_07637_ ) );
MUX2_X1 _15752_ ( .A(_06107_ ), .B(_07637_ ), .S(_05867_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_D ) );
AND3_X1 _15753_ ( .A1(_01217_ ), .A2(EXU_valid_LSU ), .A3(\mylsu.state [0] ), .ZN(\myexu.state_$_ANDNOT__A_Y ) );
INV_X1 _15754_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_07638_ ) );
AOI21_X1 _15755_ ( .A(_07638_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
INV_X1 _15756_ ( .A(\myifu.state [1] ), .ZN(_07639_ ) );
NOR3_X1 _15757_ ( .A1(_05544_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_07639_ ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__B_Y ) );
NOR2_X1 _15758_ ( .A1(_05186_ ), .A2(_05241_ ), .ZN(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OAI22_X1 _15759_ ( .A1(_05544_ ), .A2(_05187_ ), .B1(_01643_ ), .B2(IDU_ready_IFU ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
INV_X1 _15760_ ( .A(loaduse_clear ), .ZN(_07640_ ) );
NAND2_X1 _15761_ ( .A1(_07640_ ), .A2(\myidu.state [2] ), .ZN(_07641_ ) );
OAI21_X1 _15762_ ( .A(_07641_ ), .B1(_05733_ ), .B2(_01643_ ), .ZN(_07642_ ) );
NOR2_X1 _15763_ ( .A1(_05367_ ), .A2(_07639_ ), .ZN(_07643_ ) );
INV_X1 _15764_ ( .A(_07643_ ), .ZN(_07644_ ) );
AOI221_X4 _15765_ ( .A(_07642_ ), .B1(IDU_ready_IFU ), .B2(_07644_ ), .C1(_05186_ ), .C2(_07638_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
INV_X1 _15766_ ( .A(_05313_ ), .ZN(_07645_ ) );
NOR2_X1 _15767_ ( .A1(_05265_ ), .A2(_07645_ ), .ZN(_07646_ ) );
INV_X1 _15768_ ( .A(_05145_ ), .ZN(_07647_ ) );
NAND3_X1 _15769_ ( .A1(_05310_ ), .A2(_07646_ ), .A3(_07647_ ), .ZN(_07648_ ) );
AND2_X2 _15770_ ( .A1(_05179_ ), .A2(_05081_ ), .ZN(_07649_ ) );
INV_X1 _15771_ ( .A(_07649_ ), .ZN(_07650_ ) );
OAI21_X1 _15772_ ( .A(_05294_ ), .B1(_07648_ ), .B2(_07650_ ), .ZN(_07651_ ) );
OAI211_X1 _15773_ ( .A(_05243_ ), .B(_07651_ ), .C1(_05286_ ), .C2(_05301_ ), .ZN(_07652_ ) );
NAND3_X1 _15774_ ( .A1(_01051_ ), .A2(IDU_ready_IFU ), .A3(\myifu.state [1] ), .ZN(_07653_ ) );
AOI21_X1 _15775_ ( .A(_07653_ ), .B1(_05238_ ), .B2(check_quest ), .ZN(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
NAND2_X1 _15776_ ( .A1(_07652_ ), .A2(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .ZN(_00297_ ) );
NAND3_X1 _15777_ ( .A1(_01052_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_00298_ ) );
OAI211_X1 _15778_ ( .A(_00297_ ), .B(_00298_ ), .C1(_01643_ ), .C2(_05007_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _15779_ ( .A(_01052_ ), .B(IDU_ready_IFU ), .C1(_05544_ ), .C2(_07639_ ), .ZN(_00299_ ) );
NAND3_X1 _15780_ ( .A1(_00299_ ), .A2(_01329_ ), .A3(_01645_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _15781_ ( .A1(_05367_ ), .A2(_05294_ ), .A3(_07653_ ), .ZN(_00300_ ) );
OAI211_X1 _15782_ ( .A(_05243_ ), .B(_00300_ ), .C1(_05286_ ), .C2(_05301_ ), .ZN(_00301_ ) );
OAI21_X1 _15783_ ( .A(_00301_ ), .B1(fanout_net_5 ), .B2(_07641_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR4_X1 _15784_ ( .A1(_02574_ ), .A2(_01656_ ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_B ), .A4(_05714_ ), .ZN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OAI21_X1 _15785_ ( .A(_07653_ ), .B1(_01633_ ), .B2(\myifu.state [1] ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
INV_X1 _15786_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00302_ ) );
NAND2_X1 _15787_ ( .A1(_00302_ ), .A2(\IF_ID_pc [2] ), .ZN(_00303_ ) );
NAND2_X1 _15788_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00304_ ) );
NAND2_X2 _15789_ ( .A1(_00303_ ), .A2(_00304_ ), .ZN(_00305_ ) );
BUF_X4 _15790_ ( .A(_00305_ ), .Z(_00306_ ) );
MUX2_X1 _15791_ ( .A(\myifu.myicache.data[6][21] ), .B(\myifu.myicache.data[7][21] ), .S(_00306_ ), .Z(_00307_ ) );
BUF_X4 _15792_ ( .A(_00305_ ), .Z(_00308_ ) );
BUF_X4 _15793_ ( .A(_00308_ ), .Z(_00309_ ) );
MUX2_X1 _15794_ ( .A(\myifu.myicache.data[4][21] ), .B(\myifu.myicache.data[5][21] ), .S(_00309_ ), .Z(_00310_ ) );
BUF_X4 _15795_ ( .A(_05406_ ), .Z(_00311_ ) );
MUX2_X1 _15796_ ( .A(_00307_ ), .B(_00310_ ), .S(_00311_ ), .Z(_00312_ ) );
BUF_X4 _15797_ ( .A(_00308_ ), .Z(_00313_ ) );
MUX2_X1 _15798_ ( .A(\myifu.myicache.data[2][21] ), .B(\myifu.myicache.data[3][21] ), .S(_00313_ ), .Z(_00314_ ) );
BUF_X2 _15799_ ( .A(_00305_ ), .Z(_00315_ ) );
MUX2_X1 _15800_ ( .A(\myifu.myicache.data[0][21] ), .B(\myifu.myicache.data[1][21] ), .S(_00315_ ), .Z(_00316_ ) );
MUX2_X1 _15801_ ( .A(_00314_ ), .B(_00316_ ), .S(_05627_ ), .Z(_00317_ ) );
MUX2_X1 _15802_ ( .A(_00312_ ), .B(_00317_ ), .S(_05623_ ), .Z(_00318_ ) );
MUX2_X1 _15803_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_05779_ ), .Z(_00319_ ) );
AND3_X1 _15804_ ( .A1(_05686_ ), .A2(_05689_ ), .A3(_00319_ ), .ZN(_00320_ ) );
AOI21_X1 _15805_ ( .A(\io_master_rdata [21] ), .B1(_05686_ ), .B2(_05689_ ), .ZN(_00321_ ) );
NOR3_X1 _15806_ ( .A1(_00320_ ), .A2(_00321_ ), .A3(_01618_ ), .ZN(\myifu.data_in [21] ) );
XNOR2_X1 _15807_ ( .A(\IF_ID_pc [2] ), .B(\myifu.tmp_offset [2] ), .ZN(_00322_ ) );
AND2_X1 _15808_ ( .A1(_05397_ ), .A2(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .ZN(_00323_ ) );
AND2_X2 _15809_ ( .A1(_00322_ ), .A2(_00323_ ), .ZN(_00324_ ) );
BUF_X4 _15810_ ( .A(_00324_ ), .Z(_00325_ ) );
MUX2_X1 _15811_ ( .A(\IF_ID_inst [21] ), .B(\myifu.data_in [21] ), .S(_00325_ ), .Z(_00326_ ) );
MUX2_X1 _15812_ ( .A(\IF_ID_inst [21] ), .B(_00326_ ), .S(_05695_ ), .Z(_00327_ ) );
MUX2_X1 _15813_ ( .A(_00318_ ), .B(_00327_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _15814_ ( .A(\myifu.myicache.data[6][20] ), .B(\myifu.myicache.data[7][20] ), .S(_00306_ ), .Z(_00328_ ) );
MUX2_X1 _15815_ ( .A(\myifu.myicache.data[4][20] ), .B(\myifu.myicache.data[5][20] ), .S(_00309_ ), .Z(_00329_ ) );
MUX2_X1 _15816_ ( .A(_00328_ ), .B(_00329_ ), .S(_00311_ ), .Z(_00330_ ) );
MUX2_X1 _15817_ ( .A(\myifu.myicache.data[2][20] ), .B(\myifu.myicache.data[3][20] ), .S(_00309_ ), .Z(_00331_ ) );
MUX2_X1 _15818_ ( .A(\myifu.myicache.data[0][20] ), .B(\myifu.myicache.data[1][20] ), .S(_00315_ ), .Z(_00332_ ) );
MUX2_X1 _15819_ ( .A(_00331_ ), .B(_00332_ ), .S(_05627_ ), .Z(_00333_ ) );
MUX2_X1 _15820_ ( .A(_00330_ ), .B(_00333_ ), .S(_05623_ ), .Z(_00334_ ) );
OR2_X1 _15821_ ( .A1(_05697_ ), .A2(\io_master_rdata [20] ), .ZN(_00335_ ) );
CLKBUF_X2 _15822_ ( .A(_05777_ ), .Z(_00336_ ) );
OR3_X1 _15823_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00337_ ) );
OAI211_X1 _15824_ ( .A(_05697_ ), .B(_00337_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05779_ ), .ZN(_00338_ ) );
AND3_X1 _15825_ ( .A1(_00335_ ), .A2(_00338_ ), .A3(_05731_ ), .ZN(\myifu.data_in [20] ) );
MUX2_X1 _15826_ ( .A(\IF_ID_inst [20] ), .B(\myifu.data_in [20] ), .S(_00325_ ), .Z(_00339_ ) );
MUX2_X1 _15827_ ( .A(\IF_ID_inst [20] ), .B(_00339_ ), .S(_05695_ ), .Z(_00340_ ) );
MUX2_X1 _15828_ ( .A(_00334_ ), .B(_00340_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _15829_ ( .A(\myifu.myicache.data[6][19] ), .B(\myifu.myicache.data[7][19] ), .S(_00306_ ), .Z(_00341_ ) );
MUX2_X1 _15830_ ( .A(\myifu.myicache.data[4][19] ), .B(\myifu.myicache.data[5][19] ), .S(_00309_ ), .Z(_00342_ ) );
BUF_X4 _15831_ ( .A(_05406_ ), .Z(_00343_ ) );
MUX2_X1 _15832_ ( .A(_00341_ ), .B(_00342_ ), .S(_00343_ ), .Z(_00344_ ) );
MUX2_X1 _15833_ ( .A(\myifu.myicache.data[2][19] ), .B(\myifu.myicache.data[3][19] ), .S(_00309_ ), .Z(_00345_ ) );
MUX2_X1 _15834_ ( .A(\myifu.myicache.data[0][19] ), .B(\myifu.myicache.data[1][19] ), .S(_00315_ ), .Z(_00346_ ) );
MUX2_X1 _15835_ ( .A(_00345_ ), .B(_00346_ ), .S(_05627_ ), .Z(_00347_ ) );
MUX2_X1 _15836_ ( .A(_00344_ ), .B(_00347_ ), .S(_05623_ ), .Z(_00348_ ) );
CLKBUF_X2 _15837_ ( .A(_05698_ ), .Z(_00349_ ) );
OR2_X1 _15838_ ( .A1(_00349_ ), .A2(\io_master_rdata [19] ), .ZN(_00350_ ) );
BUF_X4 _15839_ ( .A(_05698_ ), .Z(_00351_ ) );
CLKBUF_X2 _15840_ ( .A(_05729_ ), .Z(_00352_ ) );
CLKBUF_X2 _15841_ ( .A(_00336_ ), .Z(_00353_ ) );
OR3_X1 _15842_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00354_ ) );
OAI211_X1 _15843_ ( .A(_00351_ ), .B(_00354_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00355_ ) );
AND3_X1 _15844_ ( .A1(_00350_ ), .A2(_00355_ ), .A3(_05731_ ), .ZN(\myifu.data_in [19] ) );
MUX2_X1 _15845_ ( .A(\IF_ID_inst [19] ), .B(\myifu.data_in [19] ), .S(_00325_ ), .Z(_00356_ ) );
MUX2_X1 _15846_ ( .A(\IF_ID_inst [19] ), .B(_00356_ ), .S(_05695_ ), .Z(_00357_ ) );
MUX2_X1 _15847_ ( .A(_00348_ ), .B(_00357_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _15848_ ( .A(\myifu.myicache.data[6][18] ), .B(\myifu.myicache.data[7][18] ), .S(_00306_ ), .Z(_00358_ ) );
MUX2_X1 _15849_ ( .A(\myifu.myicache.data[4][18] ), .B(\myifu.myicache.data[5][18] ), .S(_00309_ ), .Z(_00359_ ) );
MUX2_X1 _15850_ ( .A(_00358_ ), .B(_00359_ ), .S(_00343_ ), .Z(_00360_ ) );
MUX2_X1 _15851_ ( .A(\myifu.myicache.data[2][18] ), .B(\myifu.myicache.data[3][18] ), .S(_00309_ ), .Z(_00361_ ) );
BUF_X4 _15852_ ( .A(_00308_ ), .Z(_00362_ ) );
MUX2_X1 _15853_ ( .A(\myifu.myicache.data[0][18] ), .B(\myifu.myicache.data[1][18] ), .S(_00362_ ), .Z(_00363_ ) );
MUX2_X1 _15854_ ( .A(_00361_ ), .B(_00363_ ), .S(_05627_ ), .Z(_00364_ ) );
MUX2_X1 _15855_ ( .A(_00360_ ), .B(_00364_ ), .S(_05623_ ), .Z(_00365_ ) );
OR2_X1 _15856_ ( .A1(_00349_ ), .A2(\io_master_rdata [18] ), .ZN(_00366_ ) );
OR3_X1 _15857_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00367_ ) );
BUF_X4 _15858_ ( .A(_05779_ ), .Z(_00368_ ) );
OAI211_X1 _15859_ ( .A(_00351_ ), .B(_00367_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00369_ ) );
AND3_X1 _15860_ ( .A1(_00366_ ), .A2(_00369_ ), .A3(_05731_ ), .ZN(\myifu.data_in [18] ) );
MUX2_X1 _15861_ ( .A(\IF_ID_inst [18] ), .B(\myifu.data_in [18] ), .S(_00325_ ), .Z(_00370_ ) );
MUX2_X1 _15862_ ( .A(\IF_ID_inst [18] ), .B(_00370_ ), .S(_05695_ ), .Z(_00371_ ) );
MUX2_X1 _15863_ ( .A(_00365_ ), .B(_00371_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _15864_ ( .A(\myifu.myicache.data[6][17] ), .B(\myifu.myicache.data[7][17] ), .S(_00306_ ), .Z(_00372_ ) );
MUX2_X1 _15865_ ( .A(\myifu.myicache.data[4][17] ), .B(\myifu.myicache.data[5][17] ), .S(_00309_ ), .Z(_00373_ ) );
MUX2_X1 _15866_ ( .A(_00372_ ), .B(_00373_ ), .S(_00343_ ), .Z(_00374_ ) );
MUX2_X1 _15867_ ( .A(\myifu.myicache.data[2][17] ), .B(\myifu.myicache.data[3][17] ), .S(_00309_ ), .Z(_00375_ ) );
MUX2_X1 _15868_ ( .A(\myifu.myicache.data[0][17] ), .B(\myifu.myicache.data[1][17] ), .S(_00362_ ), .Z(_00376_ ) );
BUF_X4 _15869_ ( .A(_05406_ ), .Z(_00377_ ) );
MUX2_X1 _15870_ ( .A(_00375_ ), .B(_00376_ ), .S(_00377_ ), .Z(_00378_ ) );
BUF_X4 _15871_ ( .A(_05622_ ), .Z(_00379_ ) );
BUF_X4 _15872_ ( .A(_00379_ ), .Z(_00380_ ) );
MUX2_X1 _15873_ ( .A(_00374_ ), .B(_00378_ ), .S(_00380_ ), .Z(_00381_ ) );
OR2_X1 _15874_ ( .A1(_00349_ ), .A2(\io_master_rdata [17] ), .ZN(_00382_ ) );
CLKBUF_X2 _15875_ ( .A(_00336_ ), .Z(_00383_ ) );
OR3_X1 _15876_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00384_ ) );
OAI211_X1 _15877_ ( .A(_00351_ ), .B(_00384_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00385_ ) );
AND3_X1 _15878_ ( .A1(_00382_ ), .A2(_00385_ ), .A3(_05731_ ), .ZN(\myifu.data_in [17] ) );
MUX2_X1 _15879_ ( .A(\IF_ID_inst [17] ), .B(\myifu.data_in [17] ), .S(_00325_ ), .Z(_00386_ ) );
MUX2_X1 _15880_ ( .A(\IF_ID_inst [17] ), .B(_00386_ ), .S(_05695_ ), .Z(_00387_ ) );
MUX2_X1 _15881_ ( .A(_00381_ ), .B(_00387_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _15882_ ( .A(\myifu.myicache.data[6][16] ), .B(\myifu.myicache.data[7][16] ), .S(_00306_ ), .Z(_00388_ ) );
BUF_X4 _15883_ ( .A(_00308_ ), .Z(_00389_ ) );
MUX2_X1 _15884_ ( .A(\myifu.myicache.data[4][16] ), .B(\myifu.myicache.data[5][16] ), .S(_00389_ ), .Z(_00390_ ) );
MUX2_X1 _15885_ ( .A(_00388_ ), .B(_00390_ ), .S(_00343_ ), .Z(_00391_ ) );
MUX2_X1 _15886_ ( .A(\myifu.myicache.data[2][16] ), .B(\myifu.myicache.data[3][16] ), .S(_00309_ ), .Z(_00392_ ) );
MUX2_X1 _15887_ ( .A(\myifu.myicache.data[0][16] ), .B(\myifu.myicache.data[1][16] ), .S(_00362_ ), .Z(_00393_ ) );
MUX2_X1 _15888_ ( .A(_00392_ ), .B(_00393_ ), .S(_00377_ ), .Z(_00394_ ) );
MUX2_X1 _15889_ ( .A(_00391_ ), .B(_00394_ ), .S(_00380_ ), .Z(_00395_ ) );
OR2_X1 _15890_ ( .A1(_00349_ ), .A2(\io_master_rdata [16] ), .ZN(_00396_ ) );
OR3_X1 _15891_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00397_ ) );
OAI211_X1 _15892_ ( .A(_00351_ ), .B(_00397_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00398_ ) );
AND3_X1 _15893_ ( .A1(_00396_ ), .A2(_00398_ ), .A3(_05731_ ), .ZN(\myifu.data_in [16] ) );
MUX2_X1 _15894_ ( .A(\IF_ID_inst [16] ), .B(\myifu.data_in [16] ), .S(_00325_ ), .Z(_00399_ ) );
MUX2_X1 _15895_ ( .A(\IF_ID_inst [16] ), .B(_00399_ ), .S(_05695_ ), .Z(_00400_ ) );
MUX2_X1 _15896_ ( .A(_00395_ ), .B(_00400_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _15897_ ( .A(\myifu.myicache.data[6][15] ), .B(\myifu.myicache.data[7][15] ), .S(_00306_ ), .Z(_00401_ ) );
MUX2_X1 _15898_ ( .A(\myifu.myicache.data[4][15] ), .B(\myifu.myicache.data[5][15] ), .S(_00389_ ), .Z(_00402_ ) );
MUX2_X1 _15899_ ( .A(_00401_ ), .B(_00402_ ), .S(_00343_ ), .Z(_00403_ ) );
MUX2_X1 _15900_ ( .A(\myifu.myicache.data[2][15] ), .B(\myifu.myicache.data[3][15] ), .S(_00389_ ), .Z(_00404_ ) );
MUX2_X1 _15901_ ( .A(\myifu.myicache.data[0][15] ), .B(\myifu.myicache.data[1][15] ), .S(_00362_ ), .Z(_00405_ ) );
MUX2_X1 _15902_ ( .A(_00404_ ), .B(_00405_ ), .S(_00377_ ), .Z(_00406_ ) );
MUX2_X1 _15903_ ( .A(_00403_ ), .B(_00406_ ), .S(_00380_ ), .Z(_00407_ ) );
OR3_X1 _15904_ ( .A1(_01533_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00408_ ) );
OAI211_X1 _15905_ ( .A(_05697_ ), .B(_00408_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05778_ ), .ZN(_00409_ ) );
OAI21_X1 _15906_ ( .A(_00409_ ), .B1(_05697_ ), .B2(\io_master_rdata [15] ), .ZN(_00410_ ) );
NOR2_X1 _15907_ ( .A1(_00410_ ), .A2(_05755_ ), .ZN(\myifu.data_in [15] ) );
MUX2_X1 _15908_ ( .A(\IF_ID_inst [15] ), .B(\myifu.data_in [15] ), .S(_00325_ ), .Z(_00411_ ) );
MUX2_X1 _15909_ ( .A(\IF_ID_inst [15] ), .B(_00411_ ), .S(_05695_ ), .Z(_00412_ ) );
MUX2_X1 _15910_ ( .A(_00407_ ), .B(_00412_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_16_D ) );
BUF_X4 _15911_ ( .A(_00305_ ), .Z(_00413_ ) );
MUX2_X1 _15912_ ( .A(\myifu.myicache.data[6][14] ), .B(\myifu.myicache.data[7][14] ), .S(_00413_ ), .Z(_00414_ ) );
MUX2_X1 _15913_ ( .A(\myifu.myicache.data[4][14] ), .B(\myifu.myicache.data[5][14] ), .S(_00389_ ), .Z(_00415_ ) );
MUX2_X1 _15914_ ( .A(_00414_ ), .B(_00415_ ), .S(_00343_ ), .Z(_00416_ ) );
MUX2_X1 _15915_ ( .A(\myifu.myicache.data[2][14] ), .B(\myifu.myicache.data[3][14] ), .S(_00389_ ), .Z(_00417_ ) );
MUX2_X1 _15916_ ( .A(\myifu.myicache.data[0][14] ), .B(\myifu.myicache.data[1][14] ), .S(_00362_ ), .Z(_00418_ ) );
MUX2_X1 _15917_ ( .A(_00417_ ), .B(_00418_ ), .S(_00377_ ), .Z(_00419_ ) );
MUX2_X1 _15918_ ( .A(_00416_ ), .B(_00419_ ), .S(_00380_ ), .Z(_00420_ ) );
OR3_X1 _15919_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00421_ ) );
OAI211_X1 _15920_ ( .A(_05698_ ), .B(_00421_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05779_ ), .ZN(_00422_ ) );
BUF_X2 _15921_ ( .A(_05698_ ), .Z(_00423_ ) );
OAI21_X1 _15922_ ( .A(_00422_ ), .B1(_00423_ ), .B2(\io_master_rdata [14] ), .ZN(_00424_ ) );
NOR2_X1 _15923_ ( .A1(_00424_ ), .A2(_05755_ ), .ZN(\myifu.data_in [14] ) );
MUX2_X1 _15924_ ( .A(\IF_ID_inst [14] ), .B(\myifu.data_in [14] ), .S(_00325_ ), .Z(_00425_ ) );
MUX2_X1 _15925_ ( .A(\IF_ID_inst [14] ), .B(_00425_ ), .S(_05695_ ), .Z(_00426_ ) );
MUX2_X1 _15926_ ( .A(_00420_ ), .B(_00426_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _15927_ ( .A(\myifu.myicache.data[6][13] ), .B(\myifu.myicache.data[7][13] ), .S(_00413_ ), .Z(_00427_ ) );
MUX2_X1 _15928_ ( .A(\myifu.myicache.data[4][13] ), .B(\myifu.myicache.data[5][13] ), .S(_00389_ ), .Z(_00428_ ) );
MUX2_X1 _15929_ ( .A(_00427_ ), .B(_00428_ ), .S(_00343_ ), .Z(_00429_ ) );
MUX2_X1 _15930_ ( .A(\myifu.myicache.data[2][13] ), .B(\myifu.myicache.data[3][13] ), .S(_00389_ ), .Z(_00430_ ) );
MUX2_X1 _15931_ ( .A(\myifu.myicache.data[0][13] ), .B(\myifu.myicache.data[1][13] ), .S(_00362_ ), .Z(_00431_ ) );
MUX2_X1 _15932_ ( .A(_00430_ ), .B(_00431_ ), .S(_00377_ ), .Z(_00432_ ) );
MUX2_X1 _15933_ ( .A(_00429_ ), .B(_00432_ ), .S(_00380_ ), .Z(_00433_ ) );
OR2_X1 _15934_ ( .A1(_00349_ ), .A2(\io_master_rdata [13] ), .ZN(_00434_ ) );
OR3_X1 _15935_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00435_ ) );
OAI211_X1 _15936_ ( .A(_00423_ ), .B(_00435_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00436_ ) );
AND3_X1 _15937_ ( .A1(_00434_ ), .A2(_00436_ ), .A3(_05731_ ), .ZN(\myifu.data_in [13] ) );
MUX2_X1 _15938_ ( .A(\IF_ID_inst [13] ), .B(\myifu.data_in [13] ), .S(_00325_ ), .Z(_00437_ ) );
MUX2_X1 _15939_ ( .A(\IF_ID_inst [13] ), .B(_00437_ ), .S(_05695_ ), .Z(_00438_ ) );
MUX2_X1 _15940_ ( .A(_00433_ ), .B(_00438_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _15941_ ( .A(\myifu.myicache.data[6][12] ), .B(\myifu.myicache.data[7][12] ), .S(_00413_ ), .Z(_00439_ ) );
MUX2_X1 _15942_ ( .A(\myifu.myicache.data[4][12] ), .B(\myifu.myicache.data[5][12] ), .S(_00389_ ), .Z(_00440_ ) );
MUX2_X1 _15943_ ( .A(_00439_ ), .B(_00440_ ), .S(_00343_ ), .Z(_00441_ ) );
MUX2_X1 _15944_ ( .A(\myifu.myicache.data[2][12] ), .B(\myifu.myicache.data[3][12] ), .S(_00389_ ), .Z(_00442_ ) );
MUX2_X1 _15945_ ( .A(\myifu.myicache.data[0][12] ), .B(\myifu.myicache.data[1][12] ), .S(_00362_ ), .Z(_00443_ ) );
MUX2_X1 _15946_ ( .A(_00442_ ), .B(_00443_ ), .S(_00377_ ), .Z(_00444_ ) );
MUX2_X1 _15947_ ( .A(_00441_ ), .B(_00444_ ), .S(_00380_ ), .Z(_00445_ ) );
OR2_X1 _15948_ ( .A1(_00349_ ), .A2(\io_master_rdata [12] ), .ZN(_00446_ ) );
OR3_X1 _15949_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00447_ ) );
OAI211_X1 _15950_ ( .A(_00351_ ), .B(_00447_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00448_ ) );
CLKBUF_X2 _15951_ ( .A(_05730_ ), .Z(_00449_ ) );
AND3_X1 _15952_ ( .A1(_00446_ ), .A2(_00448_ ), .A3(_00449_ ), .ZN(\myifu.data_in [12] ) );
MUX2_X1 _15953_ ( .A(\IF_ID_inst [12] ), .B(\myifu.data_in [12] ), .S(_00325_ ), .Z(_00450_ ) );
BUF_X4 _15954_ ( .A(_05694_ ), .Z(_00451_ ) );
MUX2_X1 _15955_ ( .A(\IF_ID_inst [12] ), .B(_00450_ ), .S(_00451_ ), .Z(_00452_ ) );
MUX2_X1 _15956_ ( .A(_00445_ ), .B(_00452_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_19_D ) );
MUX2_X1 _15957_ ( .A(\myifu.myicache.data[6][30] ), .B(\myifu.myicache.data[7][30] ), .S(_00413_ ), .Z(_00453_ ) );
BUF_X4 _15958_ ( .A(_00305_ ), .Z(_00454_ ) );
MUX2_X1 _15959_ ( .A(\myifu.myicache.data[4][30] ), .B(\myifu.myicache.data[5][30] ), .S(_00454_ ), .Z(_00455_ ) );
MUX2_X1 _15960_ ( .A(_00453_ ), .B(_00455_ ), .S(_00343_ ), .Z(_00456_ ) );
MUX2_X1 _15961_ ( .A(\myifu.myicache.data[2][30] ), .B(\myifu.myicache.data[3][30] ), .S(_00389_ ), .Z(_00457_ ) );
MUX2_X1 _15962_ ( .A(\myifu.myicache.data[0][30] ), .B(\myifu.myicache.data[1][30] ), .S(_00362_ ), .Z(_00458_ ) );
MUX2_X1 _15963_ ( .A(_00457_ ), .B(_00458_ ), .S(_00377_ ), .Z(_00459_ ) );
MUX2_X1 _15964_ ( .A(_00456_ ), .B(_00459_ ), .S(_00380_ ), .Z(_00460_ ) );
OR3_X1 _15965_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00461_ ) );
OAI21_X1 _15966_ ( .A(_00461_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_05779_ ), .ZN(_00462_ ) );
MUX2_X1 _15967_ ( .A(\io_master_rdata [30] ), .B(_00462_ ), .S(_04994_ ), .Z(_00463_ ) );
AND2_X1 _15968_ ( .A1(_00463_ ), .A2(_05731_ ), .ZN(\myifu.data_in [30] ) );
BUF_X4 _15969_ ( .A(_00324_ ), .Z(_00464_ ) );
MUX2_X1 _15970_ ( .A(\IF_ID_inst [30] ), .B(\myifu.data_in [30] ), .S(_00464_ ), .Z(_00465_ ) );
MUX2_X1 _15971_ ( .A(\IF_ID_inst [30] ), .B(_00465_ ), .S(_00451_ ), .Z(_00466_ ) );
MUX2_X1 _15972_ ( .A(_00460_ ), .B(_00466_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _15973_ ( .A(\myifu.myicache.data[6][11] ), .B(\myifu.myicache.data[7][11] ), .S(_00413_ ), .Z(_00467_ ) );
MUX2_X1 _15974_ ( .A(\myifu.myicache.data[4][11] ), .B(\myifu.myicache.data[5][11] ), .S(_00454_ ), .Z(_00468_ ) );
MUX2_X1 _15975_ ( .A(_00467_ ), .B(_00468_ ), .S(_00343_ ), .Z(_00469_ ) );
MUX2_X1 _15976_ ( .A(\myifu.myicache.data[2][11] ), .B(\myifu.myicache.data[3][11] ), .S(_00454_ ), .Z(_00470_ ) );
MUX2_X1 _15977_ ( .A(\myifu.myicache.data[0][11] ), .B(\myifu.myicache.data[1][11] ), .S(_00362_ ), .Z(_00471_ ) );
MUX2_X1 _15978_ ( .A(_00470_ ), .B(_00471_ ), .S(_00377_ ), .Z(_00472_ ) );
MUX2_X1 _15979_ ( .A(_00469_ ), .B(_00472_ ), .S(_00380_ ), .Z(_00473_ ) );
OR2_X1 _15980_ ( .A1(_00423_ ), .A2(\io_master_rdata [11] ), .ZN(_00474_ ) );
OR3_X1 _15981_ ( .A1(_05730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00475_ ) );
OAI211_X1 _15982_ ( .A(_00351_ ), .B(_00475_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00476_ ) );
AND3_X1 _15983_ ( .A1(_00474_ ), .A2(_00476_ ), .A3(_00449_ ), .ZN(\myifu.data_in [11] ) );
MUX2_X1 _15984_ ( .A(\IF_ID_inst [11] ), .B(\myifu.data_in [11] ), .S(_00464_ ), .Z(_00477_ ) );
MUX2_X1 _15985_ ( .A(\IF_ID_inst [11] ), .B(_00477_ ), .S(_00451_ ), .Z(_00478_ ) );
MUX2_X1 _15986_ ( .A(_00473_ ), .B(_00478_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _15987_ ( .A(\myifu.myicache.data[6][10] ), .B(\myifu.myicache.data[7][10] ), .S(_00413_ ), .Z(_00479_ ) );
MUX2_X1 _15988_ ( .A(\myifu.myicache.data[4][10] ), .B(\myifu.myicache.data[5][10] ), .S(_00454_ ), .Z(_00480_ ) );
BUF_X4 _15989_ ( .A(_05406_ ), .Z(_00481_ ) );
MUX2_X1 _15990_ ( .A(_00479_ ), .B(_00480_ ), .S(_00481_ ), .Z(_00482_ ) );
MUX2_X1 _15991_ ( .A(\myifu.myicache.data[2][10] ), .B(\myifu.myicache.data[3][10] ), .S(_00454_ ), .Z(_00483_ ) );
MUX2_X1 _15992_ ( .A(\myifu.myicache.data[0][10] ), .B(\myifu.myicache.data[1][10] ), .S(_00362_ ), .Z(_00484_ ) );
MUX2_X1 _15993_ ( .A(_00483_ ), .B(_00484_ ), .S(_00377_ ), .Z(_00485_ ) );
MUX2_X1 _15994_ ( .A(_00482_ ), .B(_00485_ ), .S(_00380_ ), .Z(_00486_ ) );
OR2_X1 _15995_ ( .A1(_00349_ ), .A2(\io_master_rdata [10] ), .ZN(_00487_ ) );
OR3_X1 _15996_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00488_ ) );
OAI211_X1 _15997_ ( .A(_00423_ ), .B(_00488_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00489_ ) );
AND3_X1 _15998_ ( .A1(_00487_ ), .A2(_00489_ ), .A3(_00449_ ), .ZN(\myifu.data_in [10] ) );
MUX2_X1 _15999_ ( .A(\IF_ID_inst [10] ), .B(\myifu.data_in [10] ), .S(_00464_ ), .Z(_00490_ ) );
MUX2_X1 _16000_ ( .A(\IF_ID_inst [10] ), .B(_00490_ ), .S(_00451_ ), .Z(_00491_ ) );
MUX2_X1 _16001_ ( .A(_00486_ ), .B(_00491_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _16002_ ( .A(\myifu.myicache.data[6][9] ), .B(\myifu.myicache.data[7][9] ), .S(_00413_ ), .Z(_00492_ ) );
MUX2_X1 _16003_ ( .A(\myifu.myicache.data[4][9] ), .B(\myifu.myicache.data[5][9] ), .S(_00454_ ), .Z(_00493_ ) );
MUX2_X1 _16004_ ( .A(_00492_ ), .B(_00493_ ), .S(_00481_ ), .Z(_00494_ ) );
MUX2_X1 _16005_ ( .A(\myifu.myicache.data[2][9] ), .B(\myifu.myicache.data[3][9] ), .S(_00454_ ), .Z(_00495_ ) );
BUF_X4 _16006_ ( .A(_00308_ ), .Z(_00496_ ) );
MUX2_X1 _16007_ ( .A(\myifu.myicache.data[0][9] ), .B(\myifu.myicache.data[1][9] ), .S(_00496_ ), .Z(_00497_ ) );
MUX2_X1 _16008_ ( .A(_00495_ ), .B(_00497_ ), .S(_00377_ ), .Z(_00498_ ) );
MUX2_X1 _16009_ ( .A(_00494_ ), .B(_00498_ ), .S(_00380_ ), .Z(_00499_ ) );
OR2_X1 _16010_ ( .A1(_00423_ ), .A2(\io_master_rdata [9] ), .ZN(_00500_ ) );
OR3_X1 _16011_ ( .A1(_05730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00501_ ) );
OAI211_X1 _16012_ ( .A(_00351_ ), .B(_00501_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00502_ ) );
AND3_X1 _16013_ ( .A1(_00500_ ), .A2(_00502_ ), .A3(_00449_ ), .ZN(\myifu.data_in [9] ) );
MUX2_X1 _16014_ ( .A(\IF_ID_inst [9] ), .B(\myifu.data_in [9] ), .S(_00464_ ), .Z(_00503_ ) );
MUX2_X1 _16015_ ( .A(\IF_ID_inst [9] ), .B(_00503_ ), .S(_00451_ ), .Z(_00504_ ) );
MUX2_X1 _16016_ ( .A(_00499_ ), .B(_00504_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _16017_ ( .A(\myifu.myicache.data[6][8] ), .B(\myifu.myicache.data[7][8] ), .S(_00413_ ), .Z(_00505_ ) );
MUX2_X1 _16018_ ( .A(\myifu.myicache.data[4][8] ), .B(\myifu.myicache.data[5][8] ), .S(_00454_ ), .Z(_00506_ ) );
MUX2_X1 _16019_ ( .A(_00505_ ), .B(_00506_ ), .S(_00481_ ), .Z(_00507_ ) );
MUX2_X1 _16020_ ( .A(\myifu.myicache.data[2][8] ), .B(\myifu.myicache.data[3][8] ), .S(_00454_ ), .Z(_00508_ ) );
MUX2_X1 _16021_ ( .A(\myifu.myicache.data[0][8] ), .B(\myifu.myicache.data[1][8] ), .S(_00496_ ), .Z(_00509_ ) );
BUF_X4 _16022_ ( .A(_05406_ ), .Z(_00510_ ) );
MUX2_X1 _16023_ ( .A(_00508_ ), .B(_00509_ ), .S(_00510_ ), .Z(_00511_ ) );
BUF_X4 _16024_ ( .A(_00379_ ), .Z(_00512_ ) );
MUX2_X1 _16025_ ( .A(_00507_ ), .B(_00511_ ), .S(_00512_ ), .Z(_00513_ ) );
OR2_X1 _16026_ ( .A1(_00423_ ), .A2(\io_master_rdata [8] ), .ZN(_00514_ ) );
OR3_X1 _16027_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00515_ ) );
OAI211_X1 _16028_ ( .A(_00351_ ), .B(_00515_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00516_ ) );
AND3_X1 _16029_ ( .A1(_00514_ ), .A2(_00516_ ), .A3(_00449_ ), .ZN(\myifu.data_in [8] ) );
MUX2_X1 _16030_ ( .A(\IF_ID_inst [8] ), .B(\myifu.data_in [8] ), .S(_00464_ ), .Z(_00517_ ) );
MUX2_X1 _16031_ ( .A(\IF_ID_inst [8] ), .B(_00517_ ), .S(_00451_ ), .Z(_00518_ ) );
MUX2_X1 _16032_ ( .A(_00513_ ), .B(_00518_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _16033_ ( .A(\myifu.myicache.data[6][7] ), .B(\myifu.myicache.data[7][7] ), .S(_00413_ ), .Z(_00519_ ) );
BUF_X4 _16034_ ( .A(_00305_ ), .Z(_00520_ ) );
MUX2_X1 _16035_ ( .A(\myifu.myicache.data[4][7] ), .B(\myifu.myicache.data[5][7] ), .S(_00520_ ), .Z(_00521_ ) );
MUX2_X1 _16036_ ( .A(_00519_ ), .B(_00521_ ), .S(_00481_ ), .Z(_00522_ ) );
MUX2_X1 _16037_ ( .A(\myifu.myicache.data[2][7] ), .B(\myifu.myicache.data[3][7] ), .S(_00454_ ), .Z(_00523_ ) );
MUX2_X1 _16038_ ( .A(\myifu.myicache.data[0][7] ), .B(\myifu.myicache.data[1][7] ), .S(_00496_ ), .Z(_00524_ ) );
MUX2_X1 _16039_ ( .A(_00523_ ), .B(_00524_ ), .S(_00510_ ), .Z(_00525_ ) );
MUX2_X1 _16040_ ( .A(_00522_ ), .B(_00525_ ), .S(_00512_ ), .Z(_00526_ ) );
OR2_X2 _16041_ ( .A1(_05696_ ), .A2(\io_master_rdata [7] ), .ZN(_00527_ ) );
OR3_X1 _16042_ ( .A1(_01533_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05777_ ), .ZN(_00528_ ) );
OAI211_X1 _16043_ ( .A(_05696_ ), .B(_00528_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05778_ ), .ZN(_00529_ ) );
AND3_X1 _16044_ ( .A1(_00527_ ), .A2(_00529_ ), .A3(_00449_ ), .ZN(\myifu.data_in [7] ) );
MUX2_X1 _16045_ ( .A(\IF_ID_inst [7] ), .B(\myifu.data_in [7] ), .S(_00464_ ), .Z(_00530_ ) );
MUX2_X1 _16046_ ( .A(\IF_ID_inst [7] ), .B(_00530_ ), .S(_00451_ ), .Z(_00531_ ) );
MUX2_X1 _16047_ ( .A(_00526_ ), .B(_00531_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _16048_ ( .A(\myifu.myicache.data[6][6] ), .B(\myifu.myicache.data[7][6] ), .S(_00413_ ), .Z(_00532_ ) );
MUX2_X1 _16049_ ( .A(\myifu.myicache.data[4][6] ), .B(\myifu.myicache.data[5][6] ), .S(_00520_ ), .Z(_00533_ ) );
MUX2_X1 _16050_ ( .A(_00532_ ), .B(_00533_ ), .S(_00481_ ), .Z(_00534_ ) );
MUX2_X1 _16051_ ( .A(\myifu.myicache.data[2][6] ), .B(\myifu.myicache.data[3][6] ), .S(_00520_ ), .Z(_00535_ ) );
MUX2_X1 _16052_ ( .A(\myifu.myicache.data[0][6] ), .B(\myifu.myicache.data[1][6] ), .S(_00496_ ), .Z(_00536_ ) );
MUX2_X1 _16053_ ( .A(_00535_ ), .B(_00536_ ), .S(_00510_ ), .Z(_00537_ ) );
MUX2_X1 _16054_ ( .A(_00534_ ), .B(_00537_ ), .S(_00512_ ), .Z(_00538_ ) );
OR3_X1 _16055_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00539_ ) );
OAI211_X1 _16056_ ( .A(_05697_ ), .B(_00539_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05779_ ), .ZN(_00540_ ) );
OAI21_X1 _16057_ ( .A(_00540_ ), .B1(_05698_ ), .B2(\io_master_rdata [6] ), .ZN(_00541_ ) );
BUF_X4 _16058_ ( .A(_01618_ ), .Z(_00542_ ) );
NOR2_X1 _16059_ ( .A1(_00541_ ), .A2(_00542_ ), .ZN(\myifu.data_in [6] ) );
MUX2_X1 _16060_ ( .A(\IF_ID_inst [6] ), .B(\myifu.data_in [6] ), .S(_00464_ ), .Z(_00543_ ) );
MUX2_X1 _16061_ ( .A(\IF_ID_inst [6] ), .B(_00543_ ), .S(_00451_ ), .Z(_00544_ ) );
MUX2_X1 _16062_ ( .A(_00538_ ), .B(_00544_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_25_D ) );
BUF_X4 _16063_ ( .A(_00305_ ), .Z(_00545_ ) );
MUX2_X1 _16064_ ( .A(\myifu.myicache.data[6][5] ), .B(\myifu.myicache.data[7][5] ), .S(_00545_ ), .Z(_00546_ ) );
MUX2_X1 _16065_ ( .A(\myifu.myicache.data[4][5] ), .B(\myifu.myicache.data[5][5] ), .S(_00520_ ), .Z(_00547_ ) );
MUX2_X1 _16066_ ( .A(_00546_ ), .B(_00547_ ), .S(_00481_ ), .Z(_00548_ ) );
MUX2_X1 _16067_ ( .A(\myifu.myicache.data[2][5] ), .B(\myifu.myicache.data[3][5] ), .S(_00520_ ), .Z(_00549_ ) );
MUX2_X1 _16068_ ( .A(\myifu.myicache.data[0][5] ), .B(\myifu.myicache.data[1][5] ), .S(_00496_ ), .Z(_00550_ ) );
MUX2_X1 _16069_ ( .A(_00549_ ), .B(_00550_ ), .S(_00510_ ), .Z(_00551_ ) );
MUX2_X1 _16070_ ( .A(_00548_ ), .B(_00551_ ), .S(_00512_ ), .Z(_00552_ ) );
OR3_X1 _16071_ ( .A1(_05730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00553_ ) );
OAI211_X1 _16072_ ( .A(_00351_ ), .B(_00553_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00554_ ) );
OAI21_X1 _16073_ ( .A(_00554_ ), .B1(_05699_ ), .B2(\io_master_rdata [5] ), .ZN(_00555_ ) );
NOR2_X1 _16074_ ( .A1(_00555_ ), .A2(_00542_ ), .ZN(\myifu.data_in [5] ) );
MUX2_X1 _16075_ ( .A(\IF_ID_inst [5] ), .B(\myifu.data_in [5] ), .S(_00464_ ), .Z(_00556_ ) );
MUX2_X1 _16076_ ( .A(\IF_ID_inst [5] ), .B(_00556_ ), .S(_00451_ ), .Z(_00557_ ) );
MUX2_X1 _16077_ ( .A(_00552_ ), .B(_00557_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _16078_ ( .A(\myifu.myicache.data[6][4] ), .B(\myifu.myicache.data[7][4] ), .S(_00545_ ), .Z(_00558_ ) );
MUX2_X1 _16079_ ( .A(\myifu.myicache.data[4][4] ), .B(\myifu.myicache.data[5][4] ), .S(_00520_ ), .Z(_00559_ ) );
MUX2_X1 _16080_ ( .A(_00558_ ), .B(_00559_ ), .S(_00481_ ), .Z(_00560_ ) );
MUX2_X1 _16081_ ( .A(\myifu.myicache.data[2][4] ), .B(\myifu.myicache.data[3][4] ), .S(_00520_ ), .Z(_00561_ ) );
MUX2_X1 _16082_ ( .A(\myifu.myicache.data[0][4] ), .B(\myifu.myicache.data[1][4] ), .S(_00496_ ), .Z(_00562_ ) );
MUX2_X1 _16083_ ( .A(_00561_ ), .B(_00562_ ), .S(_00510_ ), .Z(_00563_ ) );
MUX2_X1 _16084_ ( .A(_00560_ ), .B(_00563_ ), .S(_00512_ ), .Z(_00564_ ) );
OR3_X1 _16085_ ( .A1(_01533_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00565_ ) );
OAI211_X1 _16086_ ( .A(_05697_ ), .B(_00565_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05778_ ), .ZN(_00566_ ) );
OAI21_X1 _16087_ ( .A(_00566_ ), .B1(_05697_ ), .B2(\io_master_rdata [4] ), .ZN(_00567_ ) );
NOR2_X1 _16088_ ( .A1(_00567_ ), .A2(_00542_ ), .ZN(\myifu.data_in [4] ) );
MUX2_X1 _16089_ ( .A(\IF_ID_inst [4] ), .B(\myifu.data_in [4] ), .S(_00464_ ), .Z(_00568_ ) );
MUX2_X1 _16090_ ( .A(\IF_ID_inst [4] ), .B(_00568_ ), .S(_00451_ ), .Z(_00569_ ) );
MUX2_X1 _16091_ ( .A(_00564_ ), .B(_00569_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _16092_ ( .A(\myifu.myicache.data[6][3] ), .B(\myifu.myicache.data[7][3] ), .S(_00545_ ), .Z(_00570_ ) );
MUX2_X1 _16093_ ( .A(\myifu.myicache.data[4][3] ), .B(\myifu.myicache.data[5][3] ), .S(_00520_ ), .Z(_00571_ ) );
MUX2_X1 _16094_ ( .A(_00570_ ), .B(_00571_ ), .S(_00481_ ), .Z(_00572_ ) );
MUX2_X1 _16095_ ( .A(\myifu.myicache.data[2][3] ), .B(\myifu.myicache.data[3][3] ), .S(_00520_ ), .Z(_00573_ ) );
MUX2_X1 _16096_ ( .A(\myifu.myicache.data[0][3] ), .B(\myifu.myicache.data[1][3] ), .S(_00496_ ), .Z(_00574_ ) );
MUX2_X1 _16097_ ( .A(_00573_ ), .B(_00574_ ), .S(_00510_ ), .Z(_00575_ ) );
MUX2_X1 _16098_ ( .A(_00572_ ), .B(_00575_ ), .S(_00512_ ), .Z(_00576_ ) );
OR3_X1 _16099_ ( .A1(_05730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00577_ ) );
OAI211_X1 _16100_ ( .A(_05699_ ), .B(_00577_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00578_ ) );
OAI21_X1 _16101_ ( .A(_00578_ ), .B1(_05699_ ), .B2(\io_master_rdata [3] ), .ZN(_00579_ ) );
NOR2_X1 _16102_ ( .A1(_00579_ ), .A2(_00542_ ), .ZN(\myifu.data_in [3] ) );
MUX2_X1 _16103_ ( .A(\IF_ID_inst [3] ), .B(\myifu.data_in [3] ), .S(_00464_ ), .Z(_00580_ ) );
BUF_X4 _16104_ ( .A(_05694_ ), .Z(_00581_ ) );
MUX2_X1 _16105_ ( .A(\IF_ID_inst [3] ), .B(_00580_ ), .S(_00581_ ), .Z(_00582_ ) );
MUX2_X1 _16106_ ( .A(_00576_ ), .B(_00582_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_28_D ) );
MUX2_X1 _16107_ ( .A(\myifu.myicache.data[6][2] ), .B(\myifu.myicache.data[7][2] ), .S(_00545_ ), .Z(_00583_ ) );
BUF_X4 _16108_ ( .A(_00305_ ), .Z(_00584_ ) );
MUX2_X1 _16109_ ( .A(\myifu.myicache.data[4][2] ), .B(\myifu.myicache.data[5][2] ), .S(_00584_ ), .Z(_00585_ ) );
MUX2_X1 _16110_ ( .A(_00583_ ), .B(_00585_ ), .S(_00481_ ), .Z(_00586_ ) );
MUX2_X1 _16111_ ( .A(\myifu.myicache.data[2][2] ), .B(\myifu.myicache.data[3][2] ), .S(_00520_ ), .Z(_00587_ ) );
MUX2_X1 _16112_ ( .A(\myifu.myicache.data[0][2] ), .B(\myifu.myicache.data[1][2] ), .S(_00496_ ), .Z(_00588_ ) );
MUX2_X1 _16113_ ( .A(_00587_ ), .B(_00588_ ), .S(_00510_ ), .Z(_00589_ ) );
MUX2_X1 _16114_ ( .A(_00586_ ), .B(_00589_ ), .S(_00512_ ), .Z(_00590_ ) );
OR3_X1 _16115_ ( .A1(_05730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00591_ ) );
OAI211_X1 _16116_ ( .A(_05699_ ), .B(_00591_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00592_ ) );
OAI21_X1 _16117_ ( .A(_00592_ ), .B1(_05699_ ), .B2(\io_master_rdata [2] ), .ZN(_00593_ ) );
NOR2_X1 _16118_ ( .A1(_00593_ ), .A2(_00542_ ), .ZN(\myifu.data_in [2] ) );
BUF_X4 _16119_ ( .A(_00324_ ), .Z(_00594_ ) );
MUX2_X1 _16120_ ( .A(\IF_ID_inst [2] ), .B(\myifu.data_in [2] ), .S(_00594_ ), .Z(_00595_ ) );
MUX2_X1 _16121_ ( .A(\IF_ID_inst [2] ), .B(_00595_ ), .S(_00581_ ), .Z(_00596_ ) );
MUX2_X1 _16122_ ( .A(_00590_ ), .B(_00596_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _16123_ ( .A(\myifu.myicache.data[6][29] ), .B(\myifu.myicache.data[7][29] ), .S(_00545_ ), .Z(_00597_ ) );
MUX2_X1 _16124_ ( .A(\myifu.myicache.data[4][29] ), .B(\myifu.myicache.data[5][29] ), .S(_00584_ ), .Z(_00598_ ) );
MUX2_X1 _16125_ ( .A(_00597_ ), .B(_00598_ ), .S(_00481_ ), .Z(_00599_ ) );
MUX2_X1 _16126_ ( .A(\myifu.myicache.data[2][29] ), .B(\myifu.myicache.data[3][29] ), .S(_00584_ ), .Z(_00600_ ) );
MUX2_X1 _16127_ ( .A(\myifu.myicache.data[0][29] ), .B(\myifu.myicache.data[1][29] ), .S(_00496_ ), .Z(_00601_ ) );
MUX2_X1 _16128_ ( .A(_00600_ ), .B(_00601_ ), .S(_00510_ ), .Z(_00602_ ) );
MUX2_X1 _16129_ ( .A(_00599_ ), .B(_00602_ ), .S(_00512_ ), .Z(_00603_ ) );
OR2_X1 _16130_ ( .A1(_00349_ ), .A2(\io_master_rdata [29] ), .ZN(_00604_ ) );
OR3_X1 _16131_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00605_ ) );
OAI211_X1 _16132_ ( .A(_00423_ ), .B(_00605_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00606_ ) );
AND3_X1 _16133_ ( .A1(_00604_ ), .A2(_00606_ ), .A3(_00449_ ), .ZN(\myifu.data_in [29] ) );
MUX2_X1 _16134_ ( .A(\IF_ID_inst [29] ), .B(\myifu.data_in [29] ), .S(_00594_ ), .Z(_00607_ ) );
MUX2_X1 _16135_ ( .A(\IF_ID_inst [29] ), .B(_00607_ ), .S(_00581_ ), .Z(_00608_ ) );
MUX2_X1 _16136_ ( .A(_00603_ ), .B(_00608_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _16137_ ( .A(\myifu.myicache.data[6][1] ), .B(\myifu.myicache.data[7][1] ), .S(_00545_ ), .Z(_00609_ ) );
MUX2_X1 _16138_ ( .A(\myifu.myicache.data[4][1] ), .B(\myifu.myicache.data[5][1] ), .S(_00584_ ), .Z(_00610_ ) );
BUF_X4 _16139_ ( .A(_05406_ ), .Z(_00611_ ) );
MUX2_X1 _16140_ ( .A(_00609_ ), .B(_00610_ ), .S(_00611_ ), .Z(_00612_ ) );
MUX2_X1 _16141_ ( .A(\myifu.myicache.data[2][1] ), .B(\myifu.myicache.data[3][1] ), .S(_00584_ ), .Z(_00613_ ) );
MUX2_X1 _16142_ ( .A(\myifu.myicache.data[0][1] ), .B(\myifu.myicache.data[1][1] ), .S(_00496_ ), .Z(_00614_ ) );
MUX2_X1 _16143_ ( .A(_00613_ ), .B(_00614_ ), .S(_00510_ ), .Z(_00615_ ) );
MUX2_X1 _16144_ ( .A(_00612_ ), .B(_00615_ ), .S(_00512_ ), .Z(_00616_ ) );
OR3_X1 _16145_ ( .A1(_05730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00353_ ), .ZN(_00617_ ) );
OAI211_X1 _16146_ ( .A(_05699_ ), .B(_00617_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00618_ ) );
OAI21_X1 _16147_ ( .A(_00618_ ), .B1(_05699_ ), .B2(\io_master_rdata [1] ), .ZN(_00619_ ) );
NOR2_X1 _16148_ ( .A1(_00619_ ), .A2(_00542_ ), .ZN(\myifu.data_in [1] ) );
MUX2_X1 _16149_ ( .A(\IF_ID_inst [1] ), .B(\myifu.data_in [1] ), .S(_00594_ ), .Z(_00620_ ) );
MUX2_X1 _16150_ ( .A(\IF_ID_inst [1] ), .B(_00620_ ), .S(_00581_ ), .Z(_00621_ ) );
MUX2_X1 _16151_ ( .A(_00616_ ), .B(_00621_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _16152_ ( .A(\myifu.myicache.data[6][0] ), .B(\myifu.myicache.data[7][0] ), .S(_00545_ ), .Z(_00622_ ) );
MUX2_X1 _16153_ ( .A(\myifu.myicache.data[4][0] ), .B(\myifu.myicache.data[5][0] ), .S(_00584_ ), .Z(_00623_ ) );
MUX2_X1 _16154_ ( .A(_00622_ ), .B(_00623_ ), .S(_00611_ ), .Z(_00624_ ) );
MUX2_X1 _16155_ ( .A(\myifu.myicache.data[2][0] ), .B(\myifu.myicache.data[3][0] ), .S(_00584_ ), .Z(_00625_ ) );
MUX2_X1 _16156_ ( .A(\myifu.myicache.data[0][0] ), .B(\myifu.myicache.data[1][0] ), .S(_00313_ ), .Z(_00626_ ) );
MUX2_X1 _16157_ ( .A(_00625_ ), .B(_00626_ ), .S(_00510_ ), .Z(_00627_ ) );
MUX2_X1 _16158_ ( .A(_00624_ ), .B(_00627_ ), .S(_00512_ ), .Z(_00628_ ) );
OR3_X1 _16159_ ( .A1(_05730_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00353_ ), .ZN(_00629_ ) );
OAI211_X1 _16160_ ( .A(_00351_ ), .B(_00629_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00630_ ) );
OAI21_X1 _16161_ ( .A(_00630_ ), .B1(_05699_ ), .B2(\io_master_rdata [0] ), .ZN(_00631_ ) );
NOR2_X1 _16162_ ( .A1(_00631_ ), .A2(_00542_ ), .ZN(\myifu.data_in [0] ) );
MUX2_X1 _16163_ ( .A(\IF_ID_inst [0] ), .B(\myifu.data_in [0] ), .S(_00594_ ), .Z(_00632_ ) );
MUX2_X1 _16164_ ( .A(\IF_ID_inst [0] ), .B(_00632_ ), .S(_00581_ ), .Z(_00633_ ) );
MUX2_X1 _16165_ ( .A(_00628_ ), .B(_00633_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _16166_ ( .A(\myifu.myicache.data[6][28] ), .B(\myifu.myicache.data[7][28] ), .S(_00545_ ), .Z(_00634_ ) );
MUX2_X1 _16167_ ( .A(\myifu.myicache.data[4][28] ), .B(\myifu.myicache.data[5][28] ), .S(_00584_ ), .Z(_00635_ ) );
MUX2_X1 _16168_ ( .A(_00634_ ), .B(_00635_ ), .S(_00611_ ), .Z(_00636_ ) );
MUX2_X1 _16169_ ( .A(\myifu.myicache.data[2][28] ), .B(\myifu.myicache.data[3][28] ), .S(_00584_ ), .Z(_00637_ ) );
MUX2_X1 _16170_ ( .A(\myifu.myicache.data[0][28] ), .B(\myifu.myicache.data[1][28] ), .S(_00313_ ), .Z(_00638_ ) );
MUX2_X1 _16171_ ( .A(_00637_ ), .B(_00638_ ), .S(_00311_ ), .Z(_00639_ ) );
MUX2_X1 _16172_ ( .A(_00636_ ), .B(_00639_ ), .S(_00379_ ), .Z(_00640_ ) );
OR2_X1 _16173_ ( .A1(_05697_ ), .A2(\io_master_rdata [28] ), .ZN(_00641_ ) );
OR3_X1 _16174_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00642_ ) );
OAI211_X1 _16175_ ( .A(_05698_ ), .B(_00642_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05779_ ), .ZN(_00643_ ) );
AND3_X1 _16176_ ( .A1(_00641_ ), .A2(_00643_ ), .A3(_00449_ ), .ZN(\myifu.data_in [28] ) );
MUX2_X1 _16177_ ( .A(\IF_ID_inst [28] ), .B(\myifu.data_in [28] ), .S(_00594_ ), .Z(_00644_ ) );
MUX2_X1 _16178_ ( .A(\IF_ID_inst [28] ), .B(_00644_ ), .S(_00581_ ), .Z(_00645_ ) );
MUX2_X1 _16179_ ( .A(_00640_ ), .B(_00645_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _16180_ ( .A(\myifu.myicache.data[6][27] ), .B(\myifu.myicache.data[7][27] ), .S(_00545_ ), .Z(_00646_ ) );
BUF_X4 _16181_ ( .A(_00305_ ), .Z(_00647_ ) );
MUX2_X1 _16182_ ( .A(\myifu.myicache.data[4][27] ), .B(\myifu.myicache.data[5][27] ), .S(_00647_ ), .Z(_00648_ ) );
MUX2_X1 _16183_ ( .A(_00646_ ), .B(_00648_ ), .S(_00611_ ), .Z(_00649_ ) );
MUX2_X1 _16184_ ( .A(\myifu.myicache.data[2][27] ), .B(\myifu.myicache.data[3][27] ), .S(_00584_ ), .Z(_00650_ ) );
MUX2_X1 _16185_ ( .A(\myifu.myicache.data[0][27] ), .B(\myifu.myicache.data[1][27] ), .S(_00313_ ), .Z(_00651_ ) );
MUX2_X1 _16186_ ( .A(_00650_ ), .B(_00651_ ), .S(_00311_ ), .Z(_00652_ ) );
MUX2_X1 _16187_ ( .A(_00649_ ), .B(_00652_ ), .S(_00379_ ), .Z(_00653_ ) );
OR2_X1 _16188_ ( .A1(_00349_ ), .A2(\io_master_rdata [27] ), .ZN(_00654_ ) );
OR3_X1 _16189_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00655_ ) );
OAI211_X1 _16190_ ( .A(_00423_ ), .B(_00655_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00656_ ) );
AND3_X1 _16191_ ( .A1(_00654_ ), .A2(_00656_ ), .A3(_00449_ ), .ZN(\myifu.data_in [27] ) );
MUX2_X1 _16192_ ( .A(\IF_ID_inst [27] ), .B(\myifu.data_in [27] ), .S(_00594_ ), .Z(_00657_ ) );
MUX2_X1 _16193_ ( .A(\IF_ID_inst [27] ), .B(_00657_ ), .S(_00581_ ), .Z(_00658_ ) );
MUX2_X1 _16194_ ( .A(_00653_ ), .B(_00658_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _16195_ ( .A(\myifu.myicache.data[6][26] ), .B(\myifu.myicache.data[7][26] ), .S(_00545_ ), .Z(_00659_ ) );
MUX2_X1 _16196_ ( .A(\myifu.myicache.data[4][26] ), .B(\myifu.myicache.data[5][26] ), .S(_00647_ ), .Z(_00660_ ) );
MUX2_X1 _16197_ ( .A(_00659_ ), .B(_00660_ ), .S(_00611_ ), .Z(_00661_ ) );
MUX2_X1 _16198_ ( .A(\myifu.myicache.data[2][26] ), .B(\myifu.myicache.data[3][26] ), .S(_00647_ ), .Z(_00662_ ) );
MUX2_X1 _16199_ ( .A(\myifu.myicache.data[0][26] ), .B(\myifu.myicache.data[1][26] ), .S(_00313_ ), .Z(_00663_ ) );
MUX2_X1 _16200_ ( .A(_00662_ ), .B(_00663_ ), .S(_00311_ ), .Z(_00664_ ) );
MUX2_X1 _16201_ ( .A(_00661_ ), .B(_00664_ ), .S(_00379_ ), .Z(_00665_ ) );
OR2_X1 _16202_ ( .A1(_05698_ ), .A2(\io_master_rdata [26] ), .ZN(_00666_ ) );
OR3_X1 _16203_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00667_ ) );
OAI211_X1 _16204_ ( .A(_00423_ ), .B(_00667_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00668_ ) );
AND3_X1 _16205_ ( .A1(_00666_ ), .A2(_00668_ ), .A3(_00449_ ), .ZN(\myifu.data_in [26] ) );
MUX2_X1 _16206_ ( .A(\IF_ID_inst [26] ), .B(\myifu.data_in [26] ), .S(_00594_ ), .Z(_00669_ ) );
MUX2_X1 _16207_ ( .A(\IF_ID_inst [26] ), .B(_00669_ ), .S(_00581_ ), .Z(_00670_ ) );
MUX2_X1 _16208_ ( .A(_00665_ ), .B(_00670_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _16209_ ( .A(\myifu.myicache.data[6][25] ), .B(\myifu.myicache.data[7][25] ), .S(_00308_ ), .Z(_00671_ ) );
MUX2_X1 _16210_ ( .A(\myifu.myicache.data[4][25] ), .B(\myifu.myicache.data[5][25] ), .S(_00647_ ), .Z(_00672_ ) );
MUX2_X1 _16211_ ( .A(_00671_ ), .B(_00672_ ), .S(_00611_ ), .Z(_00673_ ) );
MUX2_X1 _16212_ ( .A(\myifu.myicache.data[2][25] ), .B(\myifu.myicache.data[3][25] ), .S(_00647_ ), .Z(_00674_ ) );
MUX2_X1 _16213_ ( .A(\myifu.myicache.data[0][25] ), .B(\myifu.myicache.data[1][25] ), .S(_00313_ ), .Z(_00675_ ) );
MUX2_X1 _16214_ ( .A(_00674_ ), .B(_00675_ ), .S(_00311_ ), .Z(_00676_ ) );
MUX2_X1 _16215_ ( .A(_00673_ ), .B(_00676_ ), .S(_00379_ ), .Z(_00677_ ) );
MUX2_X1 _16216_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_05779_ ), .Z(_00678_ ) );
OR3_X1 _16217_ ( .A1(_05673_ ), .A2(_05676_ ), .A3(_00678_ ), .ZN(_00679_ ) );
OAI21_X1 _16218_ ( .A(\io_master_rdata [25] ), .B1(_05673_ ), .B2(_05676_ ), .ZN(_00680_ ) );
AOI21_X1 _16219_ ( .A(_00542_ ), .B1(_00679_ ), .B2(_00680_ ), .ZN(\myifu.data_in [25] ) );
MUX2_X1 _16220_ ( .A(\IF_ID_inst [25] ), .B(\myifu.data_in [25] ), .S(_00594_ ), .Z(_00681_ ) );
MUX2_X1 _16221_ ( .A(\IF_ID_inst [25] ), .B(_00681_ ), .S(_00581_ ), .Z(_00682_ ) );
MUX2_X1 _16222_ ( .A(_00677_ ), .B(_00682_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _16223_ ( .A(\myifu.myicache.data[6][24] ), .B(\myifu.myicache.data[7][24] ), .S(_00308_ ), .Z(_00683_ ) );
MUX2_X1 _16224_ ( .A(\myifu.myicache.data[4][24] ), .B(\myifu.myicache.data[5][24] ), .S(_00647_ ), .Z(_00684_ ) );
MUX2_X1 _16225_ ( .A(_00683_ ), .B(_00684_ ), .S(_00611_ ), .Z(_00685_ ) );
MUX2_X1 _16226_ ( .A(\myifu.myicache.data[2][24] ), .B(\myifu.myicache.data[3][24] ), .S(_00647_ ), .Z(_00686_ ) );
MUX2_X1 _16227_ ( .A(\myifu.myicache.data[0][24] ), .B(\myifu.myicache.data[1][24] ), .S(_00313_ ), .Z(_00687_ ) );
MUX2_X1 _16228_ ( .A(_00686_ ), .B(_00687_ ), .S(_00311_ ), .Z(_00688_ ) );
MUX2_X1 _16229_ ( .A(_00685_ ), .B(_00688_ ), .S(_00379_ ), .Z(_00689_ ) );
OR2_X1 _16230_ ( .A1(_00349_ ), .A2(\io_master_rdata [24] ), .ZN(_00690_ ) );
OR3_X1 _16231_ ( .A1(_00352_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00383_ ), .ZN(_00691_ ) );
OAI211_X1 _16232_ ( .A(_00423_ ), .B(_00691_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00368_ ), .ZN(_00692_ ) );
AND3_X1 _16233_ ( .A1(_00690_ ), .A2(_00692_ ), .A3(_05730_ ), .ZN(\myifu.data_in [24] ) );
MUX2_X1 _16234_ ( .A(\IF_ID_inst [24] ), .B(\myifu.data_in [24] ), .S(_00594_ ), .Z(_00693_ ) );
MUX2_X1 _16235_ ( .A(\IF_ID_inst [24] ), .B(_00693_ ), .S(_00581_ ), .Z(_00694_ ) );
MUX2_X1 _16236_ ( .A(_00689_ ), .B(_00694_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _16237_ ( .A(\myifu.myicache.data[6][23] ), .B(\myifu.myicache.data[7][23] ), .S(_00308_ ), .Z(_00695_ ) );
MUX2_X1 _16238_ ( .A(\myifu.myicache.data[4][23] ), .B(\myifu.myicache.data[5][23] ), .S(_00647_ ), .Z(_00696_ ) );
MUX2_X1 _16239_ ( .A(_00695_ ), .B(_00696_ ), .S(_00611_ ), .Z(_00697_ ) );
MUX2_X1 _16240_ ( .A(\myifu.myicache.data[2][23] ), .B(\myifu.myicache.data[3][23] ), .S(_00647_ ), .Z(_00698_ ) );
MUX2_X1 _16241_ ( .A(\myifu.myicache.data[0][23] ), .B(\myifu.myicache.data[1][23] ), .S(_00313_ ), .Z(_00699_ ) );
MUX2_X1 _16242_ ( .A(_00698_ ), .B(_00699_ ), .S(_00311_ ), .Z(_00700_ ) );
MUX2_X1 _16243_ ( .A(_00697_ ), .B(_00700_ ), .S(_00379_ ), .Z(_00701_ ) );
OR3_X1 _16244_ ( .A1(_01533_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05777_ ), .ZN(_00702_ ) );
OAI211_X1 _16245_ ( .A(_05696_ ), .B(_00702_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05778_ ), .ZN(_00703_ ) );
OAI21_X2 _16246_ ( .A(_00703_ ), .B1(_05697_ ), .B2(\io_master_rdata [23] ), .ZN(_00704_ ) );
NOR2_X1 _16247_ ( .A1(_00704_ ), .A2(_00542_ ), .ZN(\myifu.data_in [23] ) );
MUX2_X1 _16248_ ( .A(\IF_ID_inst [23] ), .B(\myifu.data_in [23] ), .S(_00594_ ), .Z(_00705_ ) );
MUX2_X1 _16249_ ( .A(\IF_ID_inst [23] ), .B(_00705_ ), .S(_05694_ ), .Z(_00706_ ) );
MUX2_X1 _16250_ ( .A(_00701_ ), .B(_00706_ ), .S(fanout_net_39 ), .Z(\myifu.inst_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _16251_ ( .A(\myifu.myicache.data[6][22] ), .B(\myifu.myicache.data[7][22] ), .S(_00308_ ), .Z(_00707_ ) );
MUX2_X1 _16252_ ( .A(\myifu.myicache.data[4][22] ), .B(\myifu.myicache.data[5][22] ), .S(_00306_ ), .Z(_00708_ ) );
MUX2_X1 _16253_ ( .A(_00707_ ), .B(_00708_ ), .S(_00611_ ), .Z(_00709_ ) );
MUX2_X1 _16254_ ( .A(\myifu.myicache.data[2][22] ), .B(\myifu.myicache.data[3][22] ), .S(_00647_ ), .Z(_00710_ ) );
MUX2_X1 _16255_ ( .A(\myifu.myicache.data[0][22] ), .B(\myifu.myicache.data[1][22] ), .S(_00313_ ), .Z(_00711_ ) );
MUX2_X1 _16256_ ( .A(_00710_ ), .B(_00711_ ), .S(_00311_ ), .Z(_00712_ ) );
MUX2_X1 _16257_ ( .A(_00709_ ), .B(_00712_ ), .S(_00379_ ), .Z(_00713_ ) );
OR3_X1 _16258_ ( .A1(_05729_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00714_ ) );
OAI211_X1 _16259_ ( .A(_05698_ ), .B(_00714_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05779_ ), .ZN(_00715_ ) );
OAI21_X1 _16260_ ( .A(_00715_ ), .B1(\io_master_rdata [22] ), .B2(_05698_ ), .ZN(_00716_ ) );
NOR2_X1 _16261_ ( .A1(_00716_ ), .A2(_00542_ ), .ZN(\myifu.data_in [22] ) );
MUX2_X1 _16262_ ( .A(\IF_ID_inst [22] ), .B(\myifu.data_in [22] ), .S(_00324_ ), .Z(_00717_ ) );
MUX2_X1 _16263_ ( .A(\IF_ID_inst [22] ), .B(_00717_ ), .S(_05694_ ), .Z(_00718_ ) );
MUX2_X1 _16264_ ( .A(_00713_ ), .B(_00718_ ), .S(\myifu.state [2] ), .Z(\myifu.inst_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _16265_ ( .A(\myifu.myicache.data[6][31] ), .B(\myifu.myicache.data[7][31] ), .S(_00308_ ), .Z(_00719_ ) );
MUX2_X1 _16266_ ( .A(\myifu.myicache.data[4][31] ), .B(\myifu.myicache.data[5][31] ), .S(_00306_ ), .Z(_00720_ ) );
MUX2_X1 _16267_ ( .A(_00719_ ), .B(_00720_ ), .S(_00611_ ), .Z(_00721_ ) );
MUX2_X1 _16268_ ( .A(\myifu.myicache.data[2][31] ), .B(\myifu.myicache.data[3][31] ), .S(_00306_ ), .Z(_00722_ ) );
MUX2_X1 _16269_ ( .A(\myifu.myicache.data[0][31] ), .B(\myifu.myicache.data[1][31] ), .S(_00313_ ), .Z(_00723_ ) );
MUX2_X1 _16270_ ( .A(_00722_ ), .B(_00723_ ), .S(_00311_ ), .Z(_00724_ ) );
MUX2_X1 _16271_ ( .A(_00721_ ), .B(_00724_ ), .S(_00379_ ), .Z(_00725_ ) );
OR3_X1 _16272_ ( .A1(_01533_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00336_ ), .ZN(_00726_ ) );
OAI21_X1 _16273_ ( .A(_00726_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_05778_ ), .ZN(_00727_ ) );
MUX2_X1 _16274_ ( .A(\io_master_rdata [31] ), .B(_00727_ ), .S(_04994_ ), .Z(_00728_ ) );
AND2_X1 _16275_ ( .A1(_00728_ ), .A2(_05731_ ), .ZN(\myifu.data_in [31] ) );
MUX2_X1 _16276_ ( .A(\IF_ID_inst [31] ), .B(\myifu.data_in [31] ), .S(_00324_ ), .Z(_00729_ ) );
MUX2_X1 _16277_ ( .A(\IF_ID_inst [31] ), .B(_00729_ ), .S(_05694_ ), .Z(_00730_ ) );
MUX2_X1 _16278_ ( .A(_00725_ ), .B(_00730_ ), .S(\myifu.state [2] ), .Z(\myifu.inst_$_DFFE_PP__Q_D ) );
INV_X1 _16279_ ( .A(_00239_ ), .ZN(_00731_ ) );
NAND2_X1 _16280_ ( .A1(_00731_ ), .A2(_01624_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16281_ ( .A1(_05623_ ), .A2(\IF_ID_pc [3] ), .ZN(_00732_ ) );
OAI21_X1 _16282_ ( .A(_01624_ ), .B1(_00732_ ), .B2(_00302_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16283_ ( .A1(_05627_ ), .A2(\IF_ID_pc [4] ), .ZN(_00733_ ) );
OAI21_X1 _16284_ ( .A(_01624_ ), .B1(_00733_ ), .B2(_00302_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16285_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .ZN(_00734_ ) );
OAI21_X1 _16286_ ( .A(_01624_ ), .B1(_00734_ ), .B2(_00302_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
AOI221_X4 _16287_ ( .A(_05395_ ), .B1(\IF_ID_inst [16] ), .B2(_05023_ ), .C1(_07650_ ), .C2(\IF_ID_inst [8] ), .ZN(_00735_ ) );
INV_X1 _16288_ ( .A(_05263_ ), .ZN(_00736_ ) );
OAI22_X1 _16289_ ( .A1(_05146_ ), .A2(_05327_ ), .B1(_00736_ ), .B2(_05126_ ), .ZN(_00737_ ) );
NOR2_X1 _16290_ ( .A1(_05139_ ), .A2(_05140_ ), .ZN(_00738_ ) );
INV_X1 _16291_ ( .A(_00738_ ), .ZN(_00739_ ) );
AND3_X1 _16292_ ( .A1(_00737_ ), .A2(_07647_ ), .A3(_00739_ ), .ZN(_00740_ ) );
NOR3_X1 _16293_ ( .A1(_05251_ ), .A2(_05023_ ), .A3(_05254_ ), .ZN(_00741_ ) );
INV_X1 _16294_ ( .A(_05047_ ), .ZN(_00742_ ) );
AND2_X1 _16295_ ( .A1(_00742_ ), .A2(_05330_ ), .ZN(_00743_ ) );
NAND3_X1 _16296_ ( .A1(_00740_ ), .A2(_00741_ ), .A3(_00743_ ), .ZN(_00744_ ) );
NOR2_X1 _16297_ ( .A1(_05109_ ), .A2(_05117_ ), .ZN(_00745_ ) );
NAND3_X1 _16298_ ( .A1(_05179_ ), .A2(_05081_ ), .A3(_00745_ ), .ZN(_00746_ ) );
NOR2_X1 _16299_ ( .A1(_00744_ ), .A2(_00746_ ), .ZN(_00747_ ) );
INV_X1 _16300_ ( .A(_00747_ ), .ZN(_00748_ ) );
OAI21_X1 _16301_ ( .A(_00735_ ), .B1(_00748_ ), .B2(_05020_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
NAND4_X1 _16302_ ( .A1(_05296_ ), .A2(_05161_ ), .A3(_05182_ ), .A4(_05173_ ), .ZN(_00749_ ) );
NAND3_X1 _16303_ ( .A1(_05258_ ), .A2(_05183_ ), .A3(_05156_ ), .ZN(_00750_ ) );
OAI21_X1 _16304_ ( .A(_05466_ ), .B1(_00749_ ), .B2(_00750_ ), .ZN(_00751_ ) );
BUF_X4 _16305_ ( .A(_00751_ ), .Z(_00752_ ) );
AND2_X1 _16306_ ( .A1(_05109_ ), .A2(\IF_ID_inst [31] ), .ZN(_00753_ ) );
INV_X1 _16307_ ( .A(_00753_ ), .ZN(_00754_ ) );
BUF_X4 _16308_ ( .A(_00754_ ), .Z(_00755_ ) );
AND3_X1 _16309_ ( .A1(_05179_ ), .A2(_05081_ ), .A3(_05118_ ), .ZN(_00756_ ) );
OAI211_X1 _16310_ ( .A(_00752_ ), .B(_00755_ ), .C1(_05390_ ), .C2(_00756_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
OR2_X1 _16311_ ( .A1(_07649_ ), .A2(_05390_ ), .ZN(_00757_ ) );
BUF_X4 _16312_ ( .A(_00757_ ), .Z(_00758_ ) );
NAND3_X1 _16313_ ( .A1(_05115_ ), .A2(\IF_ID_inst [30] ), .A3(_05116_ ), .ZN(_00759_ ) );
NAND4_X1 _16314_ ( .A1(_00758_ ), .A2(_00755_ ), .A3(_00752_ ), .A4(_00759_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
AND2_X2 _16315_ ( .A1(_00757_ ), .A2(_00751_ ), .ZN(_00760_ ) );
OAI211_X1 _16316_ ( .A(_00760_ ), .B(_00755_ ), .C1(_05020_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
NAND3_X1 _16317_ ( .A1(_05115_ ), .A2(\IF_ID_inst [20] ), .A3(_05116_ ), .ZN(_00761_ ) );
NAND4_X1 _16318_ ( .A1(_00758_ ), .A2(_00755_ ), .A3(_00752_ ), .A4(_00761_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
OAI211_X1 _16319_ ( .A(_00758_ ), .B(_00752_ ), .C1(_05106_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI211_X1 _16320_ ( .A(_00758_ ), .B(_00752_ ), .C1(_05120_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI211_X1 _16321_ ( .A(_00758_ ), .B(_00752_ ), .C1(_05121_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI211_X1 _16322_ ( .A(_00758_ ), .B(_00752_ ), .C1(_05245_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI211_X1 _16323_ ( .A(_00758_ ), .B(_00752_ ), .C1(_05030_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI211_X1 _16324_ ( .A(_00758_ ), .B(_00752_ ), .C1(_05130_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI211_X1 _16325_ ( .A(_00758_ ), .B(_00751_ ), .C1(_05073_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI211_X1 _16326_ ( .A(_00758_ ), .B(_00751_ ), .C1(_05013_ ), .C2(_00745_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16327_ ( .A(_00760_ ), .B(_00755_ ), .C1(_05025_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
NAND3_X1 _16328_ ( .A1(_05078_ ), .A2(\IF_ID_inst [7] ), .A3(_05079_ ), .ZN(_00762_ ) );
OR2_X1 _16329_ ( .A1(_05179_ ), .A2(_05390_ ), .ZN(_00763_ ) );
NAND4_X1 _16330_ ( .A1(_00752_ ), .A2(_05436_ ), .A3(_00762_ ), .A4(_00763_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
NAND2_X1 _16331_ ( .A1(_07650_ ), .A2(\IF_ID_inst [30] ), .ZN(_00764_ ) );
OAI211_X1 _16332_ ( .A(_00764_ ), .B(_05445_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .C2(_05300_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
OAI221_X1 _16333_ ( .A(_05440_ ), .B1(_05025_ ), .B2(_07649_ ), .C1(_05300_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
OAI221_X1 _16334_ ( .A(_05426_ ), .B1(_05026_ ), .B2(_07649_ ), .C1(_05300_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
INV_X1 _16335_ ( .A(\IF_ID_inst [27] ), .ZN(_00765_ ) );
OAI221_X1 _16336_ ( .A(_05381_ ), .B1(_00765_ ), .B2(_07649_ ), .C1(_05300_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16337_ ( .A(\IF_ID_inst [26] ), .ZN(_00766_ ) );
OAI221_X1 _16338_ ( .A(_05416_ ), .B1(_00766_ ), .B2(_07649_ ), .C1(_05300_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16339_ ( .A(\IF_ID_inst [25] ), .ZN(_00767_ ) );
OAI221_X1 _16340_ ( .A(_05412_ ), .B1(_00767_ ), .B2(_07649_ ), .C1(_05300_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16341_ ( .A(_00760_ ), .B(_00755_ ), .C1(_05026_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16342_ ( .A(_00760_ ), .B(_00755_ ), .C1(_00765_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16343_ ( .A(_00760_ ), .B(_00755_ ), .C1(_00766_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16344_ ( .A(_00760_ ), .B(_00755_ ), .C1(_00767_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16345_ ( .A(_00760_ ), .B(_00755_ ), .C1(_05049_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16346_ ( .A(_00760_ ), .B(_00754_ ), .C1(_05050_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16347_ ( .A(_00760_ ), .B(_00754_ ), .C1(_05269_ ), .C2(_05335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
AOI21_X1 _16348_ ( .A(_05385_ ), .B1(_05023_ ), .B2(\IF_ID_inst [19] ), .ZN(_00768_ ) );
OAI221_X1 _16349_ ( .A(_00768_ ), .B1(_05029_ ), .B2(_07649_ ), .C1(_00748_ ), .C2(_05049_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
AOI21_X1 _16350_ ( .A(_05392_ ), .B1(_07650_ ), .B2(\IF_ID_inst [10] ), .ZN(_00769_ ) );
OAI221_X1 _16351_ ( .A(_00769_ ), .B1(_05120_ ), .B2(_05021_ ), .C1(_00748_ ), .C2(_05050_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
NAND2_X1 _16352_ ( .A1(_07650_ ), .A2(\IF_ID_inst [9] ), .ZN(_00770_ ) );
NOR2_X1 _16353_ ( .A1(_00747_ ), .A2(_05109_ ), .ZN(_00771_ ) );
OAI221_X1 _16354_ ( .A(_00770_ ), .B1(_05121_ ), .B2(_05021_ ), .C1(_00771_ ), .C2(_05269_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16355_ ( .A1(_05179_ ), .A2(_05093_ ), .ZN(_00772_ ) );
OAI221_X1 _16356_ ( .A(_00772_ ), .B1(_05030_ ), .B2(_05021_ ), .C1(_00748_ ), .C2(_05024_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
NAND2_X1 _16357_ ( .A1(_05225_ ), .A2(_05236_ ), .ZN(_00773_ ) );
INV_X1 _16358_ ( .A(_05208_ ), .ZN(_00774_ ) );
OAI211_X1 _16359_ ( .A(check_quest ), .B(\myifu.pc_$_SDFFE_PP1P__Q_E ), .C1(_00773_ ), .C2(_00774_ ), .ZN(_00775_ ) );
INV_X1 _16360_ ( .A(_00775_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
OR3_X1 _16361_ ( .A1(_07639_ ), .A2(reset ), .A3(IDU_ready_IFU ), .ZN(_00776_ ) );
NAND4_X1 _16362_ ( .A1(_01527_ ), .A2(_01450_ ), .A3(_01410_ ), .A4(_01634_ ), .ZN(_00777_ ) );
NAND2_X1 _16363_ ( .A1(_01051_ ), .A2(\myifu.state [2] ), .ZN(_00778_ ) );
OAI211_X1 _16364_ ( .A(_00776_ ), .B(_00777_ ), .C1(_05700_ ), .C2(_00778_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
AOI21_X1 _16365_ ( .A(_01626_ ), .B1(_04995_ ), .B2(_05731_ ), .ZN(_00779_ ) );
AND3_X1 _16366_ ( .A1(_01051_ ), .A2(\myidu.stall_quest_fencei ), .A3(\myifu.state [0] ), .ZN(_00780_ ) );
OR4_X1 _16367_ ( .A1(reset ), .A2(_00779_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A4(_00780_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _16368_ ( .A1(_05186_ ), .A2(reset ), .A3(_05241_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_Y ) );
OAI21_X1 _16369_ ( .A(_05239_ ), .B1(_05048_ ), .B2(_05067_ ), .ZN(_00781_ ) );
INV_X1 _16370_ ( .A(_00781_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_ORNOT__A_Y_$_NAND__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16371_ ( .A1(_05186_ ), .A2(_05241_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_2_B_$_NOR__Y_B_$_OR__Y_B_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND3_X1 _16372_ ( .A1(_05700_ ), .A2(_01246_ ), .A3(\myifu.state [2] ), .ZN(_00782_ ) );
NAND3_X1 _16373_ ( .A1(_04995_ ), .A2(\io_master_arburst [0] ), .A3(_01625_ ), .ZN(_00783_ ) );
NAND2_X1 _16374_ ( .A1(_00782_ ), .A2(_00783_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _16375_ ( .A1(_05683_ ), .A2(_05692_ ), .A3(\myifu.state [2] ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _16376_ ( .A1(_05623_ ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00315_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND3_X1 _16377_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05728_ ), .A3(_00315_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _16378_ ( .A1(\IF_ID_pc [4] ), .A2(_05727_ ), .A3(_05627_ ), .A4(_00315_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
INV_X1 _16379_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_00784_ ) );
NOR3_X1 _16380_ ( .A1(_00784_ ), .A2(_00315_ ), .A3(_00734_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
AND4_X1 _16381_ ( .A1(\IF_ID_pc [4] ), .A2(_05727_ ), .A3(\IF_ID_pc [3] ), .A4(_00315_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
NOR3_X1 _16382_ ( .A1(_00784_ ), .A2(_00733_ ), .A3(_00315_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
NOR3_X1 _16383_ ( .A1(_00784_ ), .A2(_00732_ ), .A3(_00315_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _16384_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05728_ ), .A3(_00303_ ), .A4(_00304_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
AND3_X1 _16385_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_05627_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
AND3_X1 _16386_ ( .A1(_01624_ ), .A2(_05728_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
AND3_X1 _16387_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
AND3_X1 _16388_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05623_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
INV_X1 _16389_ ( .A(\myidu.stall_quest_fencei ), .ZN(_00785_ ) );
NAND4_X1 _16390_ ( .A1(_04995_ ), .A2(_00785_ ), .A3(_01548_ ), .A4(\io_master_arburst [0] ), .ZN(_00786_ ) );
OR2_X1 _16391_ ( .A1(\myifu.wen_$_SDFFE_PP0P__Q_D ), .A2(\myifu.state [0] ), .ZN(_00787_ ) );
AOI22_X1 _16392_ ( .A1(_05700_ ), .A2(_01549_ ), .B1(_00786_ ), .B2(_00787_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
AOI221_X4 _16393_ ( .A(_01548_ ), .B1(\myidu.stall_quest_fencei ), .B2(\myifu.state [0] ), .C1(_01633_ ), .C2(_00778_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ) );
OAI22_X1 _16394_ ( .A1(_01679_ ), .A2(\EX_LS_flag [1] ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_flag [0] ), .ZN(_00788_ ) );
AOI211_X1 _16395_ ( .A(reset ), .B(_05794_ ), .C1(_05720_ ), .C2(_00788_ ), .ZN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_Y ) );
MUX2_X1 _16396_ ( .A(_05702_ ), .B(_05733_ ), .S(\mylsu.state [0] ), .Z(_00789_ ) );
NOR2_X1 _16397_ ( .A1(_05802_ ), .A2(_00789_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _16398_ ( .A1(_05802_ ), .A2(reset ), .A3(_00789_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ORNOT__B_Y_$_ANDNOT__B_Y ) );
AND2_X1 _16399_ ( .A1(_04997_ ), .A2(_05006_ ), .ZN(_00790_ ) );
NAND4_X1 _16400_ ( .A1(_04995_ ), .A2(\mylsu.state [0] ), .A3(\io_master_arid [1] ), .A4(_00790_ ), .ZN(_00791_ ) );
OAI21_X1 _16401_ ( .A(_00791_ ), .B1(_05723_ ), .B2(_05800_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND2_X1 _16402_ ( .A1(io_master_awready ), .A2(io_master_wready ), .ZN(_00792_ ) );
NOR3_X1 _16403_ ( .A1(_05719_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A3(_00792_ ), .ZN(_00793_ ) );
AND2_X1 _16404_ ( .A1(_00793_ ), .A2(_04999_ ), .ZN(_00794_ ) );
NAND4_X1 _16405_ ( .A1(_00794_ ), .A2(_01242_ ), .A3(io_master_awready ), .A4(\mylsu.state [0] ), .ZN(_00795_ ) );
NAND3_X1 _16406_ ( .A1(_01217_ ), .A2(_05790_ ), .A3(\mylsu.state [2] ), .ZN(_00796_ ) );
NAND2_X1 _16407_ ( .A1(_00795_ ), .A2(_00796_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _16408_ ( .A1(_04999_ ), .A2(\mylsu.state [0] ), .A3(_00792_ ), .ZN(_00797_ ) );
NOR3_X1 _16409_ ( .A1(_00797_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A3(_05719_ ), .ZN(_00798_ ) );
OAI21_X1 _16410_ ( .A(_01148_ ), .B1(_00798_ ), .B2(_05808_ ), .ZN(_00799_ ) );
NAND3_X1 _16411_ ( .A1(_01148_ ), .A2(io_master_wready ), .A3(\mylsu.state [2] ), .ZN(_00800_ ) );
NAND3_X1 _16412_ ( .A1(_01242_ ), .A2(io_master_awready ), .A3(\mylsu.state [4] ), .ZN(_00801_ ) );
NAND3_X1 _16413_ ( .A1(_00799_ ), .A2(_00800_ ), .A3(_00801_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
NOR3_X1 _16414_ ( .A1(_05003_ ), .A2(reset ), .A3(EXU_valid_LSU ), .ZN(_00802_ ) );
INV_X1 _16415_ ( .A(_00790_ ), .ZN(_00803_ ) );
AOI21_X1 _16416_ ( .A(_00803_ ), .B1(_04995_ ), .B2(\io_master_arid [1] ), .ZN(_00804_ ) );
AOI21_X1 _16417_ ( .A(_00802_ ), .B1(_00804_ ), .B2(\mylsu.state [0] ), .ZN(_00805_ ) );
NAND3_X1 _16418_ ( .A1(_05799_ ), .A2(_05692_ ), .A3(_00279_ ), .ZN(_00806_ ) );
AOI22_X1 _16419_ ( .A1(_05807_ ), .A2(\mylsu.state [1] ), .B1(_05719_ ), .B2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_00807_ ) );
AND3_X1 _16420_ ( .A1(_00806_ ), .A2(_01147_ ), .A3(_00807_ ), .ZN(_00808_ ) );
INV_X1 _16421_ ( .A(_00794_ ), .ZN(_00809_ ) );
NAND2_X1 _16422_ ( .A1(_01051_ ), .A2(_05000_ ), .ZN(_00810_ ) );
OR4_X1 _16423_ ( .A1(io_master_wready ), .A2(_00809_ ), .A3(_05003_ ), .A4(_00810_ ), .ZN(_00811_ ) );
NOR4_X1 _16424_ ( .A1(_04997_ ), .A2(_04999_ ), .A3(reset ), .A4(_05733_ ), .ZN(_00812_ ) );
NAND3_X1 _16425_ ( .A1(_00812_ ), .A2(\mylsu.state [0] ), .A3(_05720_ ), .ZN(_00813_ ) );
NAND4_X1 _16426_ ( .A1(_00805_ ), .A2(_00808_ ), .A3(_00811_ ), .A4(_00813_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NOR4_X1 _16427_ ( .A1(_00810_ ), .A2(_01674_ ), .A3(_05790_ ), .A4(\EX_LS_flag [2] ), .ZN(_00814_ ) );
NAND3_X1 _16428_ ( .A1(_00793_ ), .A2(\mylsu.state [0] ), .A3(_00814_ ), .ZN(_00815_ ) );
OAI21_X1 _16429_ ( .A(_00815_ ), .B1(_05004_ ), .B2(_00810_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
AND2_X2 _16430_ ( .A1(_05704_ ), .A2(_05707_ ), .ZN(_00816_ ) );
BUF_X4 _16431_ ( .A(_00816_ ), .Z(_00817_ ) );
MUX2_X1 _16432_ ( .A(\EX_LS_pc [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _16433_ ( .A(\EX_LS_pc [20] ), .B(\EX_LS_result_csreg_mem [20] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _16434_ ( .A(\EX_LS_pc [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _16435_ ( .A(\EX_LS_pc [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _16436_ ( .A(\EX_LS_pc [17] ), .B(\EX_LS_result_csreg_mem [17] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _16437_ ( .A(\EX_LS_pc [16] ), .B(\EX_LS_result_csreg_mem [16] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _16438_ ( .A(\EX_LS_pc [15] ), .B(\EX_LS_result_csreg_mem [15] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _16439_ ( .A(\EX_LS_pc [14] ), .B(\EX_LS_result_csreg_mem [14] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _16440_ ( .A(\EX_LS_pc [13] ), .B(\EX_LS_result_csreg_mem [13] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _16441_ ( .A(\EX_LS_pc [12] ), .B(\EX_LS_result_csreg_mem [12] ), .S(_00817_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
BUF_X4 _16442_ ( .A(_00816_ ), .Z(_00818_ ) );
MUX2_X1 _16443_ ( .A(\EX_LS_pc [30] ), .B(\EX_LS_result_csreg_mem [30] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _16444_ ( .A(\EX_LS_pc [11] ), .B(\EX_LS_result_csreg_mem [11] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _16445_ ( .A(\EX_LS_pc [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _16446_ ( .A(\EX_LS_pc [9] ), .B(\EX_LS_result_csreg_mem [9] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _16447_ ( .A(\EX_LS_pc [8] ), .B(\EX_LS_result_csreg_mem [8] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _16448_ ( .A(\EX_LS_pc [7] ), .B(\EX_LS_result_csreg_mem [7] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _16449_ ( .A(\EX_LS_pc [6] ), .B(\EX_LS_result_csreg_mem [6] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _16450_ ( .A(\EX_LS_pc [5] ), .B(\EX_LS_result_csreg_mem [5] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _16451_ ( .A(\EX_LS_pc [4] ), .B(\EX_LS_result_csreg_mem [4] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _16452_ ( .A(\EX_LS_pc [3] ), .B(\EX_LS_result_csreg_mem [3] ), .S(_00818_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
BUF_X4 _16453_ ( .A(_00816_ ), .Z(_00819_ ) );
MUX2_X1 _16454_ ( .A(\EX_LS_pc [2] ), .B(\EX_LS_result_csreg_mem [2] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _16455_ ( .A(\EX_LS_pc [29] ), .B(\EX_LS_result_csreg_mem [29] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _16456_ ( .A(\EX_LS_pc [1] ), .B(\EX_LS_result_csreg_mem [1] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _16457_ ( .A(\EX_LS_pc [0] ), .B(\EX_LS_result_csreg_mem [0] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _16458_ ( .A(\EX_LS_pc [28] ), .B(\EX_LS_result_csreg_mem [28] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _16459_ ( .A(\EX_LS_pc [27] ), .B(\EX_LS_result_csreg_mem [27] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _16460_ ( .A(\EX_LS_pc [26] ), .B(\EX_LS_result_csreg_mem [26] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _16461_ ( .A(\EX_LS_pc [25] ), .B(\EX_LS_result_csreg_mem [25] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _16462_ ( .A(\EX_LS_pc [24] ), .B(\EX_LS_result_csreg_mem [24] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _16463_ ( .A(\EX_LS_pc [23] ), .B(\EX_LS_result_csreg_mem [23] ), .S(_00819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _16464_ ( .A(\EX_LS_pc [22] ), .B(\EX_LS_result_csreg_mem [22] ), .S(_00816_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _16465_ ( .A(\EX_LS_pc [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_00816_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _16466_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_00820_ ) );
INV_X1 _16467_ ( .A(_00820_ ), .ZN(_00821_ ) );
NOR2_X1 _16468_ ( .A1(_05739_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_00822_ ) );
INV_X1 _16469_ ( .A(_00822_ ), .ZN(_00823_ ) );
NOR3_X1 _16470_ ( .A1(_00704_ ), .A2(_05735_ ), .A3(_00823_ ), .ZN(_00824_ ) );
NOR3_X1 _16471_ ( .A1(_00410_ ), .A2(\mylsu.araddr_tmp [1] ), .A3(_05735_ ), .ZN(_00825_ ) );
OAI21_X1 _16472_ ( .A(_00821_ ), .B1(_00824_ ), .B2(_00825_ ), .ZN(_00826_ ) );
AND3_X1 _16473_ ( .A1(_00527_ ), .A2(_00529_ ), .A3(_01540_ ), .ZN(_00827_ ) );
NAND2_X1 _16474_ ( .A1(_00827_ ), .A2(_00820_ ), .ZN(_00828_ ) );
NAND4_X1 _16475_ ( .A1(_00728_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_01622_ ), .ZN(_00829_ ) );
NAND3_X1 _16476_ ( .A1(_00826_ ), .A2(_00828_ ), .A3(_00829_ ), .ZN(_00830_ ) );
NOR2_X1 _16477_ ( .A1(\mylsu.typ_tmp [0] ), .A2(\mylsu.typ_tmp [1] ), .ZN(_00831_ ) );
AND2_X1 _16478_ ( .A1(_00831_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_00832_ ) );
BUF_X4 _16479_ ( .A(_00832_ ), .Z(_00833_ ) );
NAND2_X2 _16480_ ( .A1(_00830_ ), .A2(_00833_ ), .ZN(_00834_ ) );
AND2_X2 _16481_ ( .A1(_00834_ ), .A2(\mylsu.state [3] ), .ZN(_00835_ ) );
BUF_X4 _16482_ ( .A(_00835_ ), .Z(_00836_ ) );
NAND3_X1 _16483_ ( .A1(_00728_ ), .A2(_01540_ ), .A3(_00821_ ), .ZN(_00837_ ) );
OR3_X1 _16484_ ( .A1(_00410_ ), .A2(_05735_ ), .A3(_00821_ ), .ZN(_00838_ ) );
NAND2_X1 _16485_ ( .A1(_00837_ ), .A2(_00838_ ), .ZN(_00839_ ) );
AND2_X2 _16486_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_00840_ ) );
INV_X1 _16487_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_00841_ ) );
AND2_X1 _16488_ ( .A1(_00840_ ), .A2(_00841_ ), .ZN(_00842_ ) );
INV_X1 _16489_ ( .A(_00842_ ), .ZN(_00843_ ) );
NOR2_X1 _16490_ ( .A1(_00839_ ), .A2(_00843_ ), .ZN(_00844_ ) );
OR2_X1 _16491_ ( .A1(_00841_ ), .A2(\mylsu.typ_tmp [1] ), .ZN(_00845_ ) );
NOR2_X1 _16492_ ( .A1(_00845_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_00846_ ) );
NOR2_X1 _16493_ ( .A1(_00846_ ), .A2(_00833_ ), .ZN(_00847_ ) );
INV_X1 _16494_ ( .A(_00847_ ), .ZN(_00848_ ) );
NOR2_X1 _16495_ ( .A1(_00844_ ), .A2(_00848_ ), .ZN(_00849_ ) );
BUF_X4 _16496_ ( .A(_00849_ ), .Z(_00850_ ) );
AND2_X1 _16497_ ( .A1(_00840_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_00851_ ) );
BUF_X2 _16498_ ( .A(_00851_ ), .Z(_00852_ ) );
NOR4_X1 _16499_ ( .A1(_00320_ ), .A2(_00321_ ), .A3(_05737_ ), .A4(_00852_ ), .ZN(_00853_ ) );
BUF_X4 _16500_ ( .A(_00842_ ), .Z(_00854_ ) );
BUF_X4 _16501_ ( .A(_00854_ ), .Z(_00855_ ) );
OAI21_X1 _16502_ ( .A(_00850_ ), .B1(_00853_ ), .B2(_00855_ ), .ZN(_00856_ ) );
BUF_X4 _16503_ ( .A(_05801_ ), .Z(_00857_ ) );
AOI22_X1 _16504_ ( .A1(_00836_ ), .A2(_00856_ ), .B1(_00857_ ), .B2(_03086_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
NAND3_X1 _16505_ ( .A1(_00335_ ), .A2(_00338_ ), .A3(\io_master_arid [1] ), .ZN(_00858_ ) );
NOR2_X1 _16506_ ( .A1(_00858_ ), .A2(_00852_ ), .ZN(_00859_ ) );
OAI21_X1 _16507_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_00859_ ), .ZN(_00860_ ) );
AOI22_X1 _16508_ ( .A1(_00836_ ), .A2(_00860_ ), .B1(_00857_ ), .B2(_03081_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _16509_ ( .A1(_00350_ ), .A2(_00355_ ), .A3(_01623_ ), .ZN(_00861_ ) );
NOR2_X1 _16510_ ( .A1(_00861_ ), .A2(_00852_ ), .ZN(_00862_ ) );
OAI21_X1 _16511_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_00862_ ), .ZN(_00863_ ) );
NAND2_X1 _16512_ ( .A1(_00863_ ), .A2(_00834_ ), .ZN(_00864_ ) );
MUX2_X1 _16513_ ( .A(\EX_LS_result_reg [19] ), .B(_00864_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _16514_ ( .A1(_00366_ ), .A2(_00369_ ), .A3(_01622_ ), .ZN(_00865_ ) );
NOR2_X1 _16515_ ( .A1(_00865_ ), .A2(_00852_ ), .ZN(_00866_ ) );
OAI21_X1 _16516_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_00866_ ), .ZN(_00867_ ) );
NAND2_X1 _16517_ ( .A1(_00867_ ), .A2(_00834_ ), .ZN(_00868_ ) );
MUX2_X1 _16518_ ( .A(\EX_LS_result_reg [18] ), .B(_00868_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _16519_ ( .A1(_00382_ ), .A2(_00385_ ), .A3(_01622_ ), .ZN(_00869_ ) );
NOR2_X1 _16520_ ( .A1(_00869_ ), .A2(_00852_ ), .ZN(_00870_ ) );
OAI21_X1 _16521_ ( .A(_00849_ ), .B1(_00854_ ), .B2(_00870_ ), .ZN(_00871_ ) );
NAND2_X1 _16522_ ( .A1(_00871_ ), .A2(_00834_ ), .ZN(_00872_ ) );
MUX2_X1 _16523_ ( .A(\EX_LS_result_reg [17] ), .B(_00872_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _16524_ ( .A1(_00396_ ), .A2(_00398_ ), .A3(_01623_ ), .ZN(_00873_ ) );
NOR2_X1 _16525_ ( .A1(_00873_ ), .A2(_00852_ ), .ZN(_00874_ ) );
OAI21_X1 _16526_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_00874_ ), .ZN(_00875_ ) );
AOI22_X1 _16527_ ( .A1(_00836_ ), .A2(_00875_ ), .B1(_00857_ ), .B2(_02925_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
NOR4_X1 _16528_ ( .A1(_00410_ ), .A2(_05737_ ), .A3(_00840_ ), .A4(_00848_ ), .ZN(_00876_ ) );
AOI21_X1 _16529_ ( .A(_00876_ ), .B1(_00839_ ), .B2(_00840_ ), .ZN(_00877_ ) );
AOI22_X1 _16530_ ( .A1(_00836_ ), .A2(_00877_ ), .B1(_00857_ ), .B2(_03138_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
AND2_X1 _16531_ ( .A1(_00830_ ), .A2(_00833_ ), .ZN(_00878_ ) );
NOR2_X1 _16532_ ( .A1(_00424_ ), .A2(_05736_ ), .ZN(_00879_ ) );
INV_X1 _16533_ ( .A(_00840_ ), .ZN(_00880_ ) );
NOR2_X1 _16534_ ( .A1(_00880_ ), .A2(_00820_ ), .ZN(_00881_ ) );
OAI21_X1 _16535_ ( .A(_00847_ ), .B1(_00879_ ), .B2(_00881_ ), .ZN(_00882_ ) );
AND2_X1 _16536_ ( .A1(_00463_ ), .A2(_01622_ ), .ZN(_00883_ ) );
INV_X1 _16537_ ( .A(_00883_ ), .ZN(_00884_ ) );
AOI21_X1 _16538_ ( .A(_00882_ ), .B1(_00881_ ), .B2(_00884_ ), .ZN(_00885_ ) );
OR2_X1 _16539_ ( .A1(_00878_ ), .A2(_00885_ ), .ZN(_00886_ ) );
MUX2_X1 _16540_ ( .A(\EX_LS_result_reg [14] ), .B(_00886_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
NAND4_X1 _16541_ ( .A1(_00604_ ), .A2(_00606_ ), .A3(\io_master_arid [1] ), .A4(_00881_ ), .ZN(_00887_ ) );
NOR2_X1 _16542_ ( .A1(_05736_ ), .A2(_00881_ ), .ZN(_00888_ ) );
AND2_X1 _16543_ ( .A1(_00888_ ), .A2(_00847_ ), .ZN(_00889_ ) );
NAND3_X1 _16544_ ( .A1(_00434_ ), .A2(_00436_ ), .A3(_00889_ ), .ZN(_00890_ ) );
AND2_X1 _16545_ ( .A1(_00887_ ), .A2(_00890_ ), .ZN(_00891_ ) );
AOI22_X1 _16546_ ( .A1(_00836_ ), .A2(_00891_ ), .B1(_00857_ ), .B2(_03190_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
NAND4_X1 _16547_ ( .A1(_00641_ ), .A2(_00643_ ), .A3(\io_master_arid [1] ), .A4(_00881_ ), .ZN(_00892_ ) );
NAND3_X1 _16548_ ( .A1(_00446_ ), .A2(_00448_ ), .A3(_00889_ ), .ZN(_00893_ ) );
AND2_X1 _16549_ ( .A1(_00892_ ), .A2(_00893_ ), .ZN(_00894_ ) );
AOI22_X1 _16550_ ( .A1(_00836_ ), .A2(_00894_ ), .B1(_00857_ ), .B2(_03165_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
AND3_X1 _16551_ ( .A1(_00463_ ), .A2(_01623_ ), .A3(_00880_ ), .ZN(_00895_ ) );
OAI21_X1 _16552_ ( .A(_00849_ ), .B1(_00854_ ), .B2(_00895_ ), .ZN(_00896_ ) );
NAND2_X1 _16553_ ( .A1(_00896_ ), .A2(_00834_ ), .ZN(_00897_ ) );
MUX2_X1 _16554_ ( .A(\EX_LS_result_reg [30] ), .B(_00897_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
AND4_X1 _16555_ ( .A1(\io_master_arid [1] ), .A2(_00654_ ), .A3(_00656_ ), .A4(_00881_ ), .ZN(_00898_ ) );
AND3_X1 _16556_ ( .A1(_00474_ ), .A2(_00476_ ), .A3(_00888_ ), .ZN(_00899_ ) );
OAI21_X1 _16557_ ( .A(_00847_ ), .B1(_00898_ ), .B2(_00899_ ), .ZN(_00900_ ) );
AOI22_X1 _16558_ ( .A1(_00836_ ), .A2(_00900_ ), .B1(_00857_ ), .B2(_03218_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
NAND4_X1 _16559_ ( .A1(_00666_ ), .A2(_00668_ ), .A3(\io_master_arid [1] ), .A4(_00881_ ), .ZN(_00901_ ) );
NAND3_X1 _16560_ ( .A1(_00487_ ), .A2(_00489_ ), .A3(_00889_ ), .ZN(_00902_ ) );
AND2_X1 _16561_ ( .A1(_00901_ ), .A2(_00902_ ), .ZN(_00903_ ) );
AOI22_X1 _16562_ ( .A1(_00836_ ), .A2(_00903_ ), .B1(_00857_ ), .B2(_03243_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
AND3_X1 _16563_ ( .A1(_00500_ ), .A2(_00502_ ), .A3(_00889_ ), .ZN(_00904_ ) );
AND2_X1 _16564_ ( .A1(_00679_ ), .A2(_00680_ ), .ZN(_00905_ ) );
NOR2_X1 _16565_ ( .A1(_00905_ ), .A2(_05737_ ), .ZN(_00906_ ) );
AOI21_X1 _16566_ ( .A(_00904_ ), .B1(_00906_ ), .B2(_00881_ ), .ZN(_00907_ ) );
AOI22_X1 _16567_ ( .A1(_00836_ ), .A2(_00907_ ), .B1(_00857_ ), .B2(_03269_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
AND4_X1 _16568_ ( .A1(\io_master_arid [1] ), .A2(_00690_ ), .A3(_00692_ ), .A4(_00881_ ), .ZN(_00908_ ) );
AND3_X1 _16569_ ( .A1(_00514_ ), .A2(_00516_ ), .A3(_00888_ ), .ZN(_00909_ ) );
OAI21_X1 _16570_ ( .A(_00847_ ), .B1(_00908_ ), .B2(_00909_ ), .ZN(_00910_ ) );
AOI22_X1 _16571_ ( .A1(_00836_ ), .A2(_00910_ ), .B1(_00857_ ), .B2(_03314_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
OR3_X2 _16572_ ( .A1(_00704_ ), .A2(_05735_ ), .A3(_00820_ ), .ZN(_00911_ ) );
NAND2_X1 _16573_ ( .A1(_00911_ ), .A2(_00828_ ), .ZN(_00912_ ) );
MUX2_X1 _16574_ ( .A(_00827_ ), .B(_00912_ ), .S(_00851_ ), .Z(_00913_ ) );
MUX2_X1 _16575_ ( .A(_00912_ ), .B(_00913_ ), .S(_00843_ ), .Z(_00914_ ) );
MUX2_X1 _16576_ ( .A(_00914_ ), .B(_00830_ ), .S(_00846_ ), .Z(_00915_ ) );
MUX2_X1 _16577_ ( .A(_00915_ ), .B(_00830_ ), .S(_00833_ ), .Z(_00916_ ) );
MUX2_X1 _16578_ ( .A(\EX_LS_result_reg [7] ), .B(_00916_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
AND3_X1 _16579_ ( .A1(_00463_ ), .A2(_01622_ ), .A3(_00823_ ), .ZN(_00917_ ) );
NOR3_X1 _16580_ ( .A1(_00716_ ), .A2(_05736_ ), .A3(_00823_ ), .ZN(_00918_ ) );
OAI22_X1 _16581_ ( .A1(_00917_ ), .A2(_00918_ ), .B1(_05741_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_00919_ ) );
NOR2_X1 _16582_ ( .A1(_05741_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_00920_ ) );
NAND2_X1 _16583_ ( .A1(_00879_ ), .A2(_00920_ ), .ZN(_00921_ ) );
AOI21_X1 _16584_ ( .A(_00820_ ), .B1(_00919_ ), .B2(_00921_ ), .ZN(_00922_ ) );
NOR3_X1 _16585_ ( .A1(_00541_ ), .A2(_05735_ ), .A3(_00821_ ), .ZN(_00923_ ) );
OAI21_X1 _16586_ ( .A(_00833_ ), .B1(_00922_ ), .B2(_00923_ ), .ZN(_00924_ ) );
OAI21_X1 _16587_ ( .A(_00846_ ), .B1(_00922_ ), .B2(_00923_ ), .ZN(_00925_ ) );
NOR3_X1 _16588_ ( .A1(_00716_ ), .A2(_05736_ ), .A3(_00820_ ), .ZN(_00926_ ) );
OAI21_X1 _16589_ ( .A(_00852_ ), .B1(_00926_ ), .B2(_00923_ ), .ZN(_00927_ ) );
OR3_X1 _16590_ ( .A1(_00541_ ), .A2(_05736_ ), .A3(_00852_ ), .ZN(_00928_ ) );
AOI21_X1 _16591_ ( .A(_00854_ ), .B1(_00927_ ), .B2(_00928_ ), .ZN(_00929_ ) );
INV_X1 _16592_ ( .A(_00926_ ), .ZN(_00930_ ) );
INV_X1 _16593_ ( .A(_00923_ ), .ZN(_00931_ ) );
AOI21_X1 _16594_ ( .A(_00843_ ), .B1(_00930_ ), .B2(_00931_ ), .ZN(_00932_ ) );
OAI22_X1 _16595_ ( .A1(_00929_ ), .A2(_00932_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_00845_ ), .ZN(_00933_ ) );
AND2_X1 _16596_ ( .A1(_00925_ ), .A2(_00933_ ), .ZN(_00934_ ) );
OAI21_X1 _16597_ ( .A(_00924_ ), .B1(_00934_ ), .B2(_00833_ ), .ZN(_00935_ ) );
MUX2_X1 _16598_ ( .A(\EX_LS_result_reg [6] ), .B(_00935_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _16599_ ( .A1(_05801_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_00936_ ) );
NOR3_X1 _16600_ ( .A1(_00846_ ), .A2(_00840_ ), .A3(_00833_ ), .ZN(_00937_ ) );
NOR2_X1 _16601_ ( .A1(_00937_ ), .A2(_00820_ ), .ZN(_00938_ ) );
INV_X1 _16602_ ( .A(_00938_ ), .ZN(_00939_ ) );
AOI211_X1 _16603_ ( .A(_05702_ ), .B(_05737_ ), .C1(_00555_ ), .C2(_00939_ ), .ZN(_00940_ ) );
NOR2_X1 _16604_ ( .A1(_00847_ ), .A2(_05741_ ), .ZN(_00941_ ) );
INV_X1 _16605_ ( .A(_00941_ ), .ZN(_00942_ ) );
AND2_X1 _16606_ ( .A1(_00942_ ), .A2(_00938_ ), .ZN(_00943_ ) );
OAI21_X1 _16607_ ( .A(_00943_ ), .B1(_00320_ ), .B2(_00321_ ), .ZN(_00944_ ) );
NAND2_X1 _16608_ ( .A1(_00940_ ), .A2(_00944_ ), .ZN(_00945_ ) );
NAND3_X1 _16609_ ( .A1(_00604_ ), .A2(_00606_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_00946_ ) );
NAND3_X1 _16610_ ( .A1(_00434_ ), .A2(_00436_ ), .A3(_05739_ ), .ZN(_00947_ ) );
AND3_X1 _16611_ ( .A1(_00946_ ), .A2(_00947_ ), .A3(_00941_ ), .ZN(_00948_ ) );
OAI21_X1 _16612_ ( .A(_00936_ ), .B1(_00945_ ), .B2(_00948_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
AND4_X1 _16613_ ( .A1(_01622_ ), .A2(_00641_ ), .A3(_00643_ ), .A4(_00823_ ), .ZN(_00949_ ) );
AND4_X1 _16614_ ( .A1(_01540_ ), .A2(_00335_ ), .A3(_00338_ ), .A4(_00822_ ), .ZN(_00950_ ) );
OAI22_X1 _16615_ ( .A1(_00949_ ), .A2(_00950_ ), .B1(_05741_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_00951_ ) );
NAND4_X1 _16616_ ( .A1(_00446_ ), .A2(_00448_ ), .A3(_01622_ ), .A4(_00920_ ), .ZN(_00952_ ) );
AOI21_X1 _16617_ ( .A(_00820_ ), .B1(_00951_ ), .B2(_00952_ ), .ZN(_00953_ ) );
NOR3_X1 _16618_ ( .A1(_00567_ ), .A2(_05735_ ), .A3(_00821_ ), .ZN(_00954_ ) );
OAI21_X1 _16619_ ( .A(_00833_ ), .B1(_00953_ ), .B2(_00954_ ), .ZN(_00955_ ) );
AND4_X1 _16620_ ( .A1(_01540_ ), .A2(_00335_ ), .A3(_00338_ ), .A4(_00821_ ), .ZN(_00956_ ) );
OR2_X1 _16621_ ( .A1(_00954_ ), .A2(_00956_ ), .ZN(_00957_ ) );
AND2_X1 _16622_ ( .A1(_00957_ ), .A2(_00854_ ), .ZN(_00958_ ) );
OAI21_X1 _16623_ ( .A(_00852_ ), .B1(_00954_ ), .B2(_00956_ ), .ZN(_00959_ ) );
OR3_X1 _16624_ ( .A1(_00567_ ), .A2(_05736_ ), .A3(_00852_ ), .ZN(_00960_ ) );
AOI21_X1 _16625_ ( .A(_00854_ ), .B1(_00959_ ), .B2(_00960_ ), .ZN(_00961_ ) );
OAI22_X1 _16626_ ( .A1(_00958_ ), .A2(_00961_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_00845_ ), .ZN(_00962_ ) );
OAI21_X1 _16627_ ( .A(_00846_ ), .B1(_00953_ ), .B2(_00954_ ), .ZN(_00963_ ) );
AND2_X1 _16628_ ( .A1(_00962_ ), .A2(_00963_ ), .ZN(_00964_ ) );
OAI21_X1 _16629_ ( .A(_00955_ ), .B1(_00964_ ), .B2(_00833_ ), .ZN(_00965_ ) );
MUX2_X1 _16630_ ( .A(\EX_LS_result_reg [4] ), .B(_00965_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _16631_ ( .A1(_05801_ ), .A2(\EX_LS_result_reg [3] ), .ZN(_00966_ ) );
AND2_X1 _16632_ ( .A1(_00579_ ), .A2(_00939_ ), .ZN(_00967_ ) );
INV_X1 _16633_ ( .A(_00943_ ), .ZN(_00968_ ) );
AOI21_X1 _16634_ ( .A(_00968_ ), .B1(_00350_ ), .B2(_00355_ ), .ZN(_00969_ ) );
OR4_X1 _16635_ ( .A1(_05801_ ), .A2(_00967_ ), .A3(_05737_ ), .A4(_00969_ ), .ZN(_00970_ ) );
NAND3_X1 _16636_ ( .A1(_00654_ ), .A2(_00656_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_00971_ ) );
NAND3_X1 _16637_ ( .A1(_00474_ ), .A2(_00476_ ), .A3(_05739_ ), .ZN(_00972_ ) );
AND3_X1 _16638_ ( .A1(_00971_ ), .A2(_00972_ ), .A3(_00941_ ), .ZN(_00973_ ) );
OAI21_X1 _16639_ ( .A(_00966_ ), .B1(_00970_ ), .B2(_00973_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
AND2_X1 _16640_ ( .A1(_00593_ ), .A2(_00939_ ), .ZN(_00974_ ) );
AOI21_X1 _16641_ ( .A(_00968_ ), .B1(_00366_ ), .B2(_00369_ ), .ZN(_00975_ ) );
OR4_X1 _16642_ ( .A1(_05702_ ), .A2(_00974_ ), .A3(_05737_ ), .A4(_00975_ ), .ZN(_00976_ ) );
NAND3_X1 _16643_ ( .A1(_00666_ ), .A2(_00668_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_00977_ ) );
NAND3_X1 _16644_ ( .A1(_00487_ ), .A2(_00489_ ), .A3(_05739_ ), .ZN(_00978_ ) );
AND3_X1 _16645_ ( .A1(_00977_ ), .A2(_00978_ ), .A3(_00941_ ), .ZN(_00979_ ) );
OAI22_X1 _16646_ ( .A1(_00976_ ), .A2(_00979_ ), .B1(\mylsu.state [3] ), .B2(_03694_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
AND4_X1 _16647_ ( .A1(_01622_ ), .A2(_00604_ ), .A3(_00606_ ), .A4(_00880_ ), .ZN(_00980_ ) );
OAI21_X1 _16648_ ( .A(_00849_ ), .B1(_00854_ ), .B2(_00980_ ), .ZN(_00981_ ) );
NAND2_X1 _16649_ ( .A1(_00981_ ), .A2(_00834_ ), .ZN(_00982_ ) );
MUX2_X1 _16650_ ( .A(\EX_LS_result_reg [29] ), .B(_00982_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
AND2_X1 _16651_ ( .A1(_00619_ ), .A2(_00939_ ), .ZN(_00983_ ) );
AOI21_X1 _16652_ ( .A(_00968_ ), .B1(_00382_ ), .B2(_00385_ ), .ZN(_00984_ ) );
OR4_X1 _16653_ ( .A1(_05702_ ), .A2(_00983_ ), .A3(_05737_ ), .A4(_00984_ ), .ZN(_00985_ ) );
NAND3_X1 _16654_ ( .A1(_00500_ ), .A2(_00502_ ), .A3(_05739_ ), .ZN(_00986_ ) );
NAND3_X1 _16655_ ( .A1(_05686_ ), .A2(_05689_ ), .A3(_00678_ ), .ZN(_00987_ ) );
OAI211_X1 _16656_ ( .A(\mylsu.araddr_tmp [1] ), .B(_00987_ ), .C1(_05699_ ), .C2(\io_master_rdata [25] ), .ZN(_00988_ ) );
AND3_X1 _16657_ ( .A1(_00986_ ), .A2(_00941_ ), .A3(_00988_ ), .ZN(_00989_ ) );
OAI22_X1 _16658_ ( .A1(_00985_ ), .A2(_00989_ ), .B1(\mylsu.state [3] ), .B2(_03621_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
AND2_X1 _16659_ ( .A1(_00631_ ), .A2(_00939_ ), .ZN(_00990_ ) );
AOI21_X1 _16660_ ( .A(_00968_ ), .B1(_00396_ ), .B2(_00398_ ), .ZN(_00991_ ) );
OR4_X1 _16661_ ( .A1(_05702_ ), .A2(_00990_ ), .A3(_05737_ ), .A4(_00991_ ), .ZN(_00992_ ) );
NAND3_X1 _16662_ ( .A1(_00690_ ), .A2(_00692_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_00993_ ) );
NAND3_X1 _16663_ ( .A1(_00514_ ), .A2(_00516_ ), .A3(_05739_ ), .ZN(_00994_ ) );
AND3_X1 _16664_ ( .A1(_00993_ ), .A2(_00994_ ), .A3(_00941_ ), .ZN(_00995_ ) );
OAI22_X1 _16665_ ( .A1(_00992_ ), .A2(_00995_ ), .B1(\mylsu.state [3] ), .B2(_03647_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
AND4_X1 _16666_ ( .A1(_01622_ ), .A2(_00641_ ), .A3(_00643_ ), .A4(_00880_ ), .ZN(_00996_ ) );
OAI21_X1 _16667_ ( .A(_00849_ ), .B1(_00854_ ), .B2(_00996_ ), .ZN(_00997_ ) );
NAND2_X1 _16668_ ( .A1(_00997_ ), .A2(_00834_ ), .ZN(_00998_ ) );
MUX2_X1 _16669_ ( .A(\EX_LS_result_reg [28] ), .B(_00998_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
AND4_X1 _16670_ ( .A1(_01623_ ), .A2(_00654_ ), .A3(_00656_ ), .A4(_00880_ ), .ZN(_00999_ ) );
OAI21_X1 _16671_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_00999_ ), .ZN(_01000_ ) );
AOI22_X1 _16672_ ( .A1(_00835_ ), .A2(_01000_ ), .B1(_05801_ ), .B2(_03499_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
AND4_X1 _16673_ ( .A1(_01623_ ), .A2(_00666_ ), .A3(_00668_ ), .A4(_00880_ ), .ZN(_01001_ ) );
OAI21_X1 _16674_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_01001_ ), .ZN(_01002_ ) );
AOI22_X1 _16675_ ( .A1(_00835_ ), .A2(_01002_ ), .B1(_05801_ ), .B2(_03523_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
AOI211_X1 _16676_ ( .A(_05736_ ), .B(_00840_ ), .C1(_00679_ ), .C2(_00680_ ), .ZN(_01003_ ) );
OAI21_X1 _16677_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_01003_ ), .ZN(_01004_ ) );
AOI22_X1 _16678_ ( .A1(_00835_ ), .A2(_01004_ ), .B1(_05801_ ), .B2(_03473_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
AND4_X1 _16679_ ( .A1(_01623_ ), .A2(_00690_ ), .A3(_00692_ ), .A4(_00880_ ), .ZN(_01005_ ) );
OAI21_X1 _16680_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_01005_ ), .ZN(_01006_ ) );
AOI22_X1 _16681_ ( .A1(_00835_ ), .A2(_01006_ ), .B1(_05801_ ), .B2(_03448_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _16682_ ( .A1(_00704_ ), .A2(_05737_ ), .A3(_00840_ ), .ZN(_01007_ ) );
OAI21_X1 _16683_ ( .A(_00850_ ), .B1(_00855_ ), .B2(_01007_ ), .ZN(_01008_ ) );
AOI22_X1 _16684_ ( .A1(_00835_ ), .A2(_01008_ ), .B1(_05801_ ), .B2(_03035_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _16685_ ( .A1(_00716_ ), .A2(_05736_ ), .A3(_00840_ ), .ZN(_01009_ ) );
OAI21_X1 _16686_ ( .A(_00849_ ), .B1(_00854_ ), .B2(_01009_ ), .ZN(_01010_ ) );
NAND2_X1 _16687_ ( .A1(_01010_ ), .A2(_00834_ ), .ZN(_01011_ ) );
MUX2_X1 _16688_ ( .A(\EX_LS_result_reg [22] ), .B(_01011_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _16689_ ( .A1(_00728_ ), .A2(_01623_ ), .A3(_00880_ ), .ZN(_01012_ ) );
OAI21_X1 _16690_ ( .A(_00849_ ), .B1(_00854_ ), .B2(_01012_ ), .ZN(_01013_ ) );
NAND2_X1 _16691_ ( .A1(_01013_ ), .A2(_00834_ ), .ZN(_01014_ ) );
MUX2_X1 _16692_ ( .A(\EX_LS_result_reg [31] ), .B(_01014_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR4_X1 _16693_ ( .A1(\LS_WB_waddr_csreg [1] ), .A2(\LS_WB_waddr_csreg [0] ), .A3(\LS_WB_waddr_csreg [3] ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_01015_ ) );
AND4_X1 _16694_ ( .A1(_05847_ ), .A2(_05856_ ), .A3(_05849_ ), .A4(_01015_ ), .ZN(\mycsreg.CSReg[0]_$_DFFE_PP__Q_E ) );
AND2_X1 _16695_ ( .A1(_05848_ ), .A2(_05850_ ), .ZN(_01016_ ) );
NAND4_X1 _16696_ ( .A1(_05858_ ), .A2(_01016_ ), .A3(\LS_WB_waddr_csreg [1] ), .A4(_05853_ ), .ZN(_01017_ ) );
AOI21_X1 _16697_ ( .A(reset ), .B1(_01017_ ), .B2(_01640_ ), .ZN(_01018_ ) );
AND2_X1 _16698_ ( .A1(_01018_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(\mycsreg.CSReg[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _16699_ ( .A1(_01217_ ), .A2(IDU_valid_EXU ), .A3(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__A_Y ) );
CLKBUF_X1 _16700_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _16701_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(\LS_WB_waddr_reg [1] ), .ZN(_01019_ ) );
INV_X1 _16702_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01020_ ) );
INV_X1 _16703_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01021_ ) );
NAND3_X1 _16704_ ( .A1(_01019_ ), .A2(_01020_ ), .A3(_01021_ ), .ZN(_01022_ ) );
AND2_X1 _16705_ ( .A1(_01050_ ), .A2(LS_WB_wen_reg ), .ZN(_01023_ ) );
NAND2_X1 _16706_ ( .A1(_01022_ ), .A2(_01023_ ), .ZN(_01024_ ) );
BUF_X4 _16707_ ( .A(_01024_ ), .Z(_01025_ ) );
INV_X1 _16708_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01026_ ) );
AOI21_X1 _16709_ ( .A(_01025_ ), .B1(_01020_ ), .B2(_01026_ ), .ZN(_01027_ ) );
INV_X1 _16710_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01028_ ) );
NOR2_X1 _16711_ ( .A1(_01024_ ), .A2(_01028_ ), .ZN(_01029_ ) );
NOR4_X1 _16712_ ( .A1(_01027_ ), .A2(_01029_ ), .A3(_01021_ ), .A4(_01025_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
NOR2_X1 _16713_ ( .A1(_01025_ ), .A2(_01026_ ), .ZN(_01030_ ) );
AND4_X1 _16714_ ( .A1(_01020_ ), .A2(_01030_ ), .A3(_01029_ ), .A4(_01021_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR2_X1 _16715_ ( .A1(_01024_ ), .A2(_01020_ ), .ZN(_01031_ ) );
AND4_X1 _16716_ ( .A1(_01026_ ), .A2(_01031_ ), .A3(_01029_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
AOI21_X1 _16717_ ( .A(_01025_ ), .B1(_01028_ ), .B2(_01021_ ), .ZN(_01032_ ) );
NOR4_X1 _16718_ ( .A1(_01032_ ), .A2(_01020_ ), .A3(_01026_ ), .A4(_01025_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
NOR2_X1 _16719_ ( .A1(_01025_ ), .A2(_01021_ ), .ZN(_01033_ ) );
AND4_X1 _16720_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01031_ ), .A3(_01033_ ), .A4(_01028_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
AND4_X1 _16721_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01031_ ), .A3(_01029_ ), .A4(_01021_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
NOR4_X1 _16722_ ( .A1(_01027_ ), .A2(_01033_ ), .A3(_01028_ ), .A4(_01025_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
NOR4_X1 _16723_ ( .A1(_01027_ ), .A2(_01028_ ), .A3(_01021_ ), .A4(_01025_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _16724_ ( .A1(_01032_ ), .A2(_01031_ ), .A3(_01026_ ), .A4(_01025_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _16725_ ( .A1(_01020_ ), .A2(_01030_ ), .A3(_01029_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
NOR4_X1 _16726_ ( .A1(_01032_ ), .A2(_01030_ ), .A3(_01020_ ), .A4(_01025_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _16727_ ( .A1(_01026_ ), .A2(_01031_ ), .A3(_01033_ ), .A4(_01028_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _16728_ ( .A1(_01026_ ), .A2(_01031_ ), .A3(_01029_ ), .A4(_01021_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _16729_ ( .A1(_01020_ ), .A2(_01030_ ), .A3(_01033_ ), .A4(_01028_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
AND4_X1 _16730_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01031_ ), .A3(_01033_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _16731_ ( .A1(_01531_ ), .A2(_01217_ ), .A3(_01538_ ), .ZN(_01034_ ) );
NAND2_X1 _16732_ ( .A1(_01034_ ), .A2(_01329_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _16733_ ( .A(reset ), .B(_01531_ ), .C1(_01532_ ), .C2(_05743_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _16734_ ( .A(_01022_ ), .Z(_01035_ ) );
CLKBUF_X2 _16735_ ( .A(_01023_ ), .Z(_01036_ ) );
AND3_X1 _16736_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _16737_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _16738_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _16739_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _16740_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _16741_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _16742_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _16743_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _16744_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _16745_ ( .A1(_01035_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01036_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _16746_ ( .A(_01022_ ), .Z(_01037_ ) );
CLKBUF_X2 _16747_ ( .A(_01023_ ), .Z(_01038_ ) );
AND3_X1 _16748_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _16749_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _16750_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _16751_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _16752_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _16753_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _16754_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _16755_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _16756_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _16757_ ( .A1(_01037_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01038_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _16758_ ( .A(_01022_ ), .Z(_01039_ ) );
CLKBUF_X2 _16759_ ( .A(_01023_ ), .Z(_01040_ ) );
AND3_X1 _16760_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _16761_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _16762_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _16763_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _16764_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _16765_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _16766_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _16767_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _16768_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _16769_ ( .A1(_01039_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01040_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _16770_ ( .A1(_01022_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01023_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _16771_ ( .A1(_01022_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01023_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_D ) );
AND3_X1 _16772_ ( .A1(_01217_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _16773_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01041_ ) );
AND2_X1 _16774_ ( .A1(_01041_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01042_ ) );
INV_X1 _16775_ ( .A(_01042_ ), .ZN(_01043_ ) );
NOR2_X1 _16776_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01044_ ) );
OAI211_X1 _16777_ ( .A(_01051_ ), .B(\mysc.state [0] ), .C1(_01043_ ), .C2(_01044_ ), .ZN(_01045_ ) );
INV_X1 _16778_ ( .A(_01045_ ), .ZN(_01046_ ) );
OR3_X1 _16779_ ( .A1(_01046_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _16780_ ( .A1(_01043_ ), .A2(reset ), .A3(_01044_ ), .ZN(_01047_ ) );
NAND2_X1 _16781_ ( .A1(_01047_ ), .A2(\mysc.state [0] ), .ZN(_01048_ ) );
OR3_X1 _16782_ ( .A1(_05726_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01049_ ) );
NAND2_X1 _16783_ ( .A1(_01048_ ), .A2(_01049_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _16784_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07654_ ) );
CLKGATE_X1 _16785_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07655_ ) );
CLKGATE_X1 _16786_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07656_ ) );
CLKGATE_X1 _16787_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07657_ ) );
CLKGATE_X1 _16788_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_07658_ ) );
CLKGATE_X1 _16789_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_07659_ ) );
CLKGATE_X1 _16790_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07660_ ) );
CLKGATE_X1 _16791_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07661_ ) );
CLKGATE_X1 _16792_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07662_ ) );
CLKGATE_X1 _16793_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07663_ ) );
CLKGATE_X1 _16794_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_07664_ ) );
CLKGATE_X1 _16795_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_07665_ ) );
CLKGATE_X1 _16796_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_07666_ ) );
CLKGATE_X1 _16797_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_07667_ ) );
CLKGATE_X1 _16798_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07668_ ) );
CLKGATE_X1 _16799_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_07669_ ) );
CLKGATE_X1 _16800_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_07670_ ) );
CLKGATE_X1 _16801_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__B_Y_$_NOR__A_Y ), .GCK(_07671_ ) );
CLKGATE_X1 _16802_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ORNOT__B_Y_$_ANDNOT__B_Y ), .GCK(_07672_ ) );
CLKGATE_X1 _16803_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_Y ), .GCK(_07673_ ) );
CLKGATE_X1 _16804_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ), .GCK(_07674_ ) );
CLKGATE_X1 _16805_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .GCK(_07675_ ) );
CLKGATE_X1 _16806_ ( .CK(clock ), .E(io_master_awready_$_NOR__A_Y_$_OR__A_Y_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_07676_ ) );
CLKGATE_X1 _16807_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__A_Y ), .GCK(_07677_ ) );
CLKGATE_X1 _16808_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_07678_ ) );
CLKGATE_X1 _16809_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_07679_ ) );
CLKGATE_X1 _16810_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_07680_ ) );
CLKGATE_X1 _16811_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_07681_ ) );
CLKGATE_X1 _16812_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_07682_ ) );
CLKGATE_X1 _16813_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_07683_ ) );
CLKGATE_X1 _16814_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_07684_ ) );
CLKGATE_X1 _16815_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_07685_ ) );
CLKGATE_X1 _16816_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_07686_ ) );
CLKGATE_X1 _16817_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_07687_ ) );
CLKGATE_X1 _16818_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_07688_ ) );
CLKGATE_X1 _16819_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_07689_ ) );
CLKGATE_X1 _16820_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07690_ ) );
CLKGATE_X1 _16821_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07691_ ) );
CLKGATE_X1 _16822_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07692_ ) );
CLKGATE_X1 _16823_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07693_ ) );
CLKGATE_X1 _16824_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07694_ ) );
CLKGATE_X1 _16825_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07695_ ) );
CLKGATE_X1 _16826_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07696_ ) );
CLKGATE_X1 _16827_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07697_ ) );
CLKGATE_X1 _16828_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07698_ ) );
CLKGATE_X1 _16829_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_07699_ ) );
CLKGATE_X1 _16830_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__B_Y ), .GCK(_07700_ ) );
CLKGATE_X1 _16831_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_07701_ ) );
CLKGATE_X1 _16832_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_07702_ ) );
CLKGATE_X1 _16833_ ( .CK(clock ), .E(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07703_ ) );
CLKGATE_X1 _16834_ ( .CK(clock ), .E(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_B_$_NOR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07704_ ) );
CLKGATE_X1 _16835_ ( .CK(clock ), .E(\myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_2_B_$_NOR__Y_B_$_OR__Y_B_$_OR__A_Y_$_OR__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07705_ ) );
CLKGATE_X1 _16836_ ( .CK(clock ), .E(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_07706_ ) );
CLKGATE_X1 _16837_ ( .CK(clock ), .E(\myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_Y ), .GCK(_07707_ ) );
CLKGATE_X1 _16838_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_07708_ ) );
CLKGATE_X1 _16839_ ( .CK(clock ), .E(\myifu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_ORNOT__A_Y_$_NAND__A_Y_$_ANDNOT__B_Y ), .GCK(_07709_ ) );
CLKGATE_X1 _16840_ ( .CK(clock ), .E(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07710_ ) );
CLKGATE_X1 _16841_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_07711_ ) );
CLKGATE_X1 _16842_ ( .CK(clock ), .E(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__A_Y ), .GCK(_07712_ ) );
CLKGATE_X1 _16843_ ( .CK(clock ), .E(\mycsreg.CSReg[3]_$_DFFE_PP__Q_E ), .GCK(_07713_ ) );
CLKGATE_X1 _16844_ ( .CK(clock ), .E(\mycsreg.CSReg[2]_$_DFFE_PP__Q_E ), .GCK(_07714_ ) );
CLKGATE_X1 _16845_ ( .CK(clock ), .E(\mycsreg.CSReg[1]_$_DFFE_PP__Q_E ), .GCK(_07715_ ) );
CLKGATE_X1 _16846_ ( .CK(clock ), .E(\mycsreg.CSReg[0]_$_DFFE_PP__Q_E ), .GCK(_07716_ ) );
LOGIC1_X1 _16847_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _16848_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_07940_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_07941_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_07942_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_07943_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_07944_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_07945_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_07946_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_07947_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_07948_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_07949_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_07950_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_07951_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_07952_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_07953_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_07954_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_07955_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_07956_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_07957_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_07958_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_07959_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_07960_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_07961_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_07962_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_07963_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_07964_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_07965_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_07966_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_07967_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_07968_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_07969_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_07970_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07716_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_07971_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07715_ ), .Q(\mtvec [31] ), .QN(_07972_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07715_ ), .Q(\mtvec [30] ), .QN(_07973_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07715_ ), .Q(\mtvec [21] ), .QN(_07974_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07715_ ), .Q(\mtvec [20] ), .QN(_07975_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07715_ ), .Q(\mtvec [19] ), .QN(_07976_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07715_ ), .Q(\mtvec [18] ), .QN(_07977_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07715_ ), .Q(\mtvec [17] ), .QN(_07978_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07715_ ), .Q(\mtvec [16] ), .QN(_07979_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07715_ ), .Q(\mtvec [15] ), .QN(_07980_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07715_ ), .Q(\mtvec [14] ), .QN(_07981_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07715_ ), .Q(\mtvec [13] ), .QN(_07982_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07715_ ), .Q(\mtvec [12] ), .QN(_07983_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07715_ ), .Q(\mtvec [29] ), .QN(_07984_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07715_ ), .Q(\mtvec [11] ), .QN(_07985_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07715_ ), .Q(\mtvec [10] ), .QN(_07986_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07715_ ), .Q(\mtvec [9] ), .QN(_07987_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07715_ ), .Q(\mtvec [8] ), .QN(_07988_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07715_ ), .Q(\mtvec [7] ), .QN(_07989_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07715_ ), .Q(\mtvec [6] ), .QN(_07990_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07715_ ), .Q(\mtvec [5] ), .QN(_07991_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07715_ ), .Q(\mtvec [4] ), .QN(_07992_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07715_ ), .Q(\mtvec [3] ), .QN(_07993_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07715_ ), .Q(\mtvec [2] ), .QN(_07994_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07715_ ), .Q(\mtvec [28] ), .QN(_07995_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07715_ ), .Q(\mtvec [1] ), .QN(_07996_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07715_ ), .Q(\mtvec [0] ), .QN(_07997_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07715_ ), .Q(\mtvec [27] ), .QN(_07998_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07715_ ), .Q(\mtvec [26] ), .QN(_07999_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07715_ ), .Q(\mtvec [25] ), .QN(_08000_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07715_ ), .Q(\mtvec [24] ), .QN(_08001_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07715_ ), .Q(\mtvec [23] ), .QN(_08002_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07715_ ), .Q(\mtvec [22] ), .QN(_08003_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07714_ ), .Q(\mepc [31] ), .QN(_08004_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07714_ ), .Q(\mepc [30] ), .QN(_08005_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07714_ ), .Q(\mepc [21] ), .QN(_08006_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07714_ ), .Q(\mepc [20] ), .QN(_08007_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07714_ ), .Q(\mepc [19] ), .QN(_08008_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07714_ ), .Q(\mepc [18] ), .QN(_08009_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07714_ ), .Q(\mepc [17] ), .QN(_08010_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07714_ ), .Q(\mepc [16] ), .QN(_08011_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07714_ ), .Q(\mepc [15] ), .QN(_08012_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07714_ ), .Q(\mepc [14] ), .QN(_08013_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07714_ ), .Q(\mepc [13] ), .QN(_08014_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07714_ ), .Q(\mepc [12] ), .QN(_08015_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07714_ ), .Q(\mepc [29] ), .QN(_08016_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07714_ ), .Q(\mepc [11] ), .QN(_08017_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07714_ ), .Q(\mepc [10] ), .QN(_08018_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07714_ ), .Q(\mepc [9] ), .QN(_08019_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07714_ ), .Q(\mepc [8] ), .QN(_08020_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07714_ ), .Q(\mepc [7] ), .QN(_08021_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07714_ ), .Q(\mepc [6] ), .QN(_08022_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07714_ ), .Q(\mepc [5] ), .QN(_08023_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07714_ ), .Q(\mepc [4] ), .QN(_08024_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07714_ ), .Q(\mepc [3] ), .QN(_08025_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07714_ ), .Q(\mepc [2] ), .QN(_08026_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07714_ ), .Q(\mepc [28] ), .QN(_08027_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07714_ ), .Q(\mepc [1] ), .QN(_08028_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07714_ ), .Q(\mepc [0] ), .QN(_08029_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07714_ ), .Q(\mepc [27] ), .QN(_08030_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07714_ ), .Q(\mepc [26] ), .QN(_08031_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07714_ ), .Q(\mepc [25] ), .QN(_08032_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07714_ ), .Q(\mepc [24] ), .QN(_08033_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07714_ ), .Q(\mepc [23] ), .QN(_08034_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07714_ ), .Q(\mepc [22] ), .QN(_08035_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08036_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08037_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_07939_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_07938_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_07937_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_07936_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_07935_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_07934_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_07933_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_07932_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_07931_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_07930_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_07929_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_07928_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_07927_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_07926_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_07925_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_07924_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_07923_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_07922_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_07921_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_07920_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_07919_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_07918_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_28 ( .D(_00086_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_07917_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00087_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_07916_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00088_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_07915_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00089_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_07914_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00090_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_07913_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00091_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_07912_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00092_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_07911_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00093_ ), .CK(_07713_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08038_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PP0__Q ( .D(_00094_ ), .CK(clock ), .Q(check_quest ), .QN(_08039_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_07910_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08040_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08041_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08042_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08043_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08044_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08045_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08046_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08047_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08048_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08049_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_07909_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00095_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_07908_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00096_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_07907_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00097_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_07906_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00098_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_07905_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00099_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_07904_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00100_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_07903_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00101_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_07902_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00102_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_07901_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00103_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_07900_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00104_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_07899_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00105_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_07898_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00106_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_07897_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00107_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_07896_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00108_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_07895_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00109_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_07894_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00110_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_07893_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00111_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_07892_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00112_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_07891_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00113_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_07890_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00114_ ), .CK(_07712_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_07889_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q ( .D(_00115_ ), .CK(_07711_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_07888_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_1 ( .D(_00116_ ), .CK(_07711_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_07887_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_2 ( .D(_00117_ ), .CK(_07711_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_07886_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_3 ( .D(_00118_ ), .CK(_07711_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_07885_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_4 ( .D(_00119_ ), .CK(_07711_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_07884_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q ( .D(_00120_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [30] ), .QN(_07883_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_1 ( .D(_00121_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [29] ), .QN(_07882_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_10 ( .D(_00122_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [20] ), .QN(_07881_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_11 ( .D(_00123_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [19] ), .QN(_07880_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_12 ( .D(_00124_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [18] ), .QN(_07879_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_13 ( .D(_00125_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [17] ), .QN(_07878_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_14 ( .D(_00126_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [16] ), .QN(_07877_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_15 ( .D(_00127_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [15] ), .QN(_07876_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_16 ( .D(_00128_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [14] ), .QN(_07875_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_17 ( .D(_00129_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [13] ), .QN(_07874_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_18 ( .D(_00130_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [12] ), .QN(_07873_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_19 ( .D(_00131_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [11] ), .QN(_07872_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_2 ( .D(_00132_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [28] ), .QN(_07871_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_20 ( .D(_00133_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [10] ), .QN(_07870_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_21 ( .D(_00134_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [9] ), .QN(_07869_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_22 ( .D(_00135_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [8] ), .QN(_07868_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_23 ( .D(_00136_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [7] ), .QN(_07867_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_24 ( .D(_00137_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [6] ), .QN(_07866_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_25 ( .D(_00138_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [5] ), .QN(_07865_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_26 ( .D(_00139_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [4] ), .QN(_07864_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_27 ( .D(_00140_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [3] ), .QN(_07863_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_28 ( .D(_00141_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [2] ), .QN(_07862_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_29 ( .D(_00142_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [1] ), .QN(_07861_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_3 ( .D(_00143_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [27] ), .QN(_07860_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_30 ( .D(_00144_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [0] ), .QN(_07859_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_4 ( .D(_00145_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [26] ), .QN(_07858_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_5 ( .D(_00146_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [25] ), .QN(_07857_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_6 ( .D(_00147_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [24] ), .QN(_07856_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_7 ( .D(_00148_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [23] ), .QN(_07855_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_8 ( .D(_00149_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [22] ), .QN(_07854_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_9 ( .D(_00150_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [21] ), .QN(_07853_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP1P__Q ( .D(_00151_ ), .CK(_07710_ ), .Q(\myexu.pc_jump [31] ), .QN(_07852_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q ( .D(_00152_ ), .CK(_07711_ ), .Q(\EX_LS_pc [31] ), .QN(_07851_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_1 ( .D(_00153_ ), .CK(_07711_ ), .Q(\EX_LS_pc [30] ), .QN(_07850_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_10 ( .D(_00154_ ), .CK(_07711_ ), .Q(\EX_LS_pc [21] ), .QN(_07849_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_11 ( .D(_00155_ ), .CK(_07711_ ), .Q(\EX_LS_pc [20] ), .QN(_07848_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_12 ( .D(_00156_ ), .CK(_07711_ ), .Q(\EX_LS_pc [19] ), .QN(_07847_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_13 ( .D(_00157_ ), .CK(_07711_ ), .Q(\EX_LS_pc [18] ), .QN(_07846_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_14 ( .D(_00158_ ), .CK(_07711_ ), .Q(\EX_LS_pc [17] ), .QN(_07845_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_15 ( .D(_00159_ ), .CK(_07711_ ), .Q(\EX_LS_pc [16] ), .QN(_07844_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_16 ( .D(_00160_ ), .CK(_07711_ ), .Q(\EX_LS_pc [15] ), .QN(_07843_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_17 ( .D(_00161_ ), .CK(_07711_ ), .Q(\EX_LS_pc [14] ), .QN(_07842_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_18 ( .D(_00162_ ), .CK(_07711_ ), .Q(\EX_LS_pc [13] ), .QN(_07841_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_19 ( .D(_00163_ ), .CK(_07711_ ), .Q(\EX_LS_pc [12] ), .QN(_07840_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_2 ( .D(_00164_ ), .CK(_07711_ ), .Q(\EX_LS_pc [29] ), .QN(_07839_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_20 ( .D(_00165_ ), .CK(_07711_ ), .Q(\EX_LS_pc [11] ), .QN(_07838_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_21 ( .D(_00166_ ), .CK(_07711_ ), .Q(\EX_LS_pc [10] ), .QN(_07837_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_22 ( .D(_00167_ ), .CK(_07711_ ), .Q(\EX_LS_pc [9] ), .QN(_07836_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_23 ( .D(_00168_ ), .CK(_07711_ ), .Q(\EX_LS_pc [8] ), .QN(_07835_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_24 ( .D(_00169_ ), .CK(_07711_ ), .Q(\EX_LS_pc [7] ), .QN(_07834_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_25 ( .D(_00170_ ), .CK(_07711_ ), .Q(\EX_LS_pc [6] ), .QN(_07833_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_26 ( .D(_00171_ ), .CK(_07711_ ), .Q(\EX_LS_pc [5] ), .QN(_07832_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_27 ( .D(_00172_ ), .CK(_07711_ ), .Q(\EX_LS_pc [4] ), .QN(_07831_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_28 ( .D(_00173_ ), .CK(_07711_ ), .Q(\EX_LS_pc [3] ), .QN(_07830_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_29 ( .D(_00174_ ), .CK(_07711_ ), .Q(\EX_LS_pc [2] ), .QN(_07829_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_3 ( .D(_00175_ ), .CK(_07711_ ), .Q(\EX_LS_pc [28] ), .QN(_07828_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_30 ( .D(_00176_ ), .CK(_07711_ ), .Q(\EX_LS_pc [1] ), .QN(_07827_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_31 ( .D(_00177_ ), .CK(_07711_ ), .Q(\EX_LS_pc [0] ), .QN(_07826_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_4 ( .D(_00178_ ), .CK(_07711_ ), .Q(\EX_LS_pc [27] ), .QN(_07825_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_5 ( .D(_00179_ ), .CK(_07711_ ), .Q(\EX_LS_pc [26] ), .QN(_07824_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_6 ( .D(_00180_ ), .CK(_07711_ ), .Q(\EX_LS_pc [25] ), .QN(_07823_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_7 ( .D(_00181_ ), .CK(_07711_ ), .Q(\EX_LS_pc [24] ), .QN(_07822_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_8 ( .D(_00182_ ), .CK(_07711_ ), .Q(\EX_LS_pc [23] ), .QN(_07821_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_9 ( .D(_00183_ ), .CK(_07711_ ), .Q(\EX_LS_pc [22] ), .QN(_08050_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08051_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08052_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08053_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08054_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08055_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08056_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08057_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08058_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08059_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08060_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08061_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08062_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08063_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08064_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08065_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08066_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08067_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08068_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08069_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08070_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08071_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08072_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08073_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08074_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08075_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08076_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08077_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08078_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08079_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08080_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08081_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07712_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08082_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_07712_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PP0__Q ( .D(_00185_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q ( .D(_00184_ ), .CK(_07711_ ), .Q(\EX_LS_flag [2] ), .QN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E_$_ANDNOT__A_B_$_OR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_MUX__Y_A_$_ANDNOT__B_1_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_1 ( .D(_00186_ ), .CK(_07711_ ), .Q(\EX_LS_flag [1] ), .QN(_07820_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_2 ( .D(_00187_ ), .CK(_07711_ ), .Q(\EX_LS_flag [0] ), .QN(_07819_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_3 ( .D(_00188_ ), .CK(_07711_ ), .Q(\EX_LS_typ [4] ), .QN(_07818_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_4 ( .D(_00189_ ), .CK(_07711_ ), .Q(\EX_LS_typ [3] ), .QN(_07817_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_5 ( .D(_00190_ ), .CK(_07711_ ), .Q(\EX_LS_typ [2] ), .QN(_07816_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_6 ( .D(_00191_ ), .CK(_07711_ ), .Q(\EX_LS_typ [1] ), .QN(_07815_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_7 ( .D(_00192_ ), .CK(_07711_ ), .Q(\EX_LS_typ [0] ), .QN(_07814_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00193_ ), .CK(_07709_ ), .Q(\ID_EX_csr [11] ), .QN(_07813_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00194_ ), .CK(_07709_ ), .Q(\ID_EX_csr [10] ), .QN(_07812_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00195_ ), .CK(_07709_ ), .Q(\ID_EX_csr [1] ), .QN(_07811_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00196_ ), .CK(_07709_ ), .Q(\ID_EX_csr [0] ), .QN(_07810_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00197_ ), .CK(_07709_ ), .Q(\ID_EX_csr [9] ), .QN(_07809_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00198_ ), .CK(_07709_ ), .Q(\ID_EX_csr [8] ), .QN(_07808_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00199_ ), .CK(_07709_ ), .Q(\ID_EX_csr [7] ), .QN(_07807_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00200_ ), .CK(_07709_ ), .Q(\ID_EX_csr [6] ), .QN(_07806_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00201_ ), .CK(_07709_ ), .Q(\ID_EX_csr [5] ), .QN(_07805_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00202_ ), .CK(_07709_ ), .Q(\ID_EX_csr [4] ), .QN(_07804_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00203_ ), .CK(_07709_ ), .Q(\ID_EX_csr [3] ), .QN(_07803_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00204_ ), .CK(_07709_ ), .Q(\ID_EX_csr [2] ), .QN(_07802_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00205_ ), .CK(_07708_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_07707_ ), .Q(\ID_EX_imm [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_07707_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_07707_ ), .Q(\ID_EX_imm [21] ), .QN(_08083_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_07707_ ), .Q(\ID_EX_imm [20] ), .QN(_08084_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_07707_ ), .Q(\ID_EX_imm [19] ), .QN(_08085_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_07707_ ), .Q(\ID_EX_imm [18] ), .QN(_08086_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_07707_ ), .Q(\ID_EX_imm [17] ), .QN(_08087_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_07707_ ), .Q(\ID_EX_imm [16] ), .QN(_08088_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_07707_ ), .Q(\ID_EX_imm [15] ), .QN(_08089_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_07707_ ), .Q(\ID_EX_imm [14] ), .QN(_08090_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_07707_ ), .Q(\ID_EX_imm [13] ), .QN(_08091_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_07707_ ), .Q(\ID_EX_imm [12] ), .QN(_08092_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_07707_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_07707_ ), .Q(\ID_EX_imm [11] ), .QN(_08093_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_07707_ ), .Q(\ID_EX_imm [10] ), .QN(_08094_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_07707_ ), .Q(\ID_EX_imm [9] ), .QN(_08095_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_07707_ ), .Q(\ID_EX_imm [8] ), .QN(_08096_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_07707_ ), .Q(\ID_EX_imm [7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_07707_ ), .Q(\ID_EX_imm [6] ), .QN(_08097_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_07707_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_07707_ ), .Q(\ID_EX_imm [4] ), .QN(_08098_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_07707_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_07707_ ), .Q(\ID_EX_imm [2] ), .QN(_08099_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_07707_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_07707_ ), .Q(\ID_EX_imm [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_07707_ ), .Q(\ID_EX_imm [0] ), .QN(_08100_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_07707_ ), .Q(\ID_EX_imm [27] ), .QN(_08101_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_07707_ ), .Q(\ID_EX_imm [26] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_07707_ ), .Q(\ID_EX_imm [25] ), .QN(_08102_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_07707_ ), .Q(\ID_EX_imm [24] ), .QN(_08103_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_07707_ ), .Q(\ID_EX_imm [23] ), .QN(_08104_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_07707_ ), .Q(\ID_EX_imm [22] ), .QN(_08105_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07706_ ), .Q(\ID_EX_pc [31] ), .QN(_08106_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07706_ ), .Q(\ID_EX_pc [30] ), .QN(_08107_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07706_ ), .Q(\ID_EX_pc [21] ), .QN(_08108_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07706_ ), .Q(\ID_EX_pc [20] ), .QN(_08109_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07706_ ), .Q(\ID_EX_pc [19] ), .QN(_08110_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07706_ ), .Q(\ID_EX_pc [18] ), .QN(_08111_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07706_ ), .Q(\ID_EX_pc [17] ), .QN(_08112_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07706_ ), .Q(\ID_EX_pc [16] ), .QN(_08113_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07706_ ), .Q(\ID_EX_pc [15] ), .QN(_08114_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07706_ ), .Q(\ID_EX_pc [14] ), .QN(_08115_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07706_ ), .Q(\ID_EX_pc [13] ), .QN(_08116_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07706_ ), .Q(\ID_EX_pc [12] ), .QN(_08117_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07706_ ), .Q(\ID_EX_pc [29] ), .QN(_08118_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07706_ ), .Q(\ID_EX_pc [11] ), .QN(_08119_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07706_ ), .Q(\ID_EX_pc [10] ), .QN(_08120_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07706_ ), .Q(\ID_EX_pc [9] ), .QN(_08121_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07706_ ), .Q(\ID_EX_pc [8] ), .QN(_08122_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07706_ ), .Q(\ID_EX_pc [7] ), .QN(_08123_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07706_ ), .Q(\ID_EX_pc [6] ), .QN(_08124_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07706_ ), .Q(\ID_EX_pc [5] ), .QN(_08125_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07706_ ), .Q(\ID_EX_pc [4] ), .QN(_08126_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_07706_ ), .Q(\ID_EX_pc [3] ), .QN(_08127_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_07706_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07706_ ), .Q(\ID_EX_pc [28] ), .QN(_08128_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_07706_ ), .Q(\ID_EX_pc [1] ), .QN(_08129_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_07706_ ), .Q(\ID_EX_pc [0] ), .QN(_08130_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07706_ ), .Q(\ID_EX_pc [27] ), .QN(_08131_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07706_ ), .Q(\ID_EX_pc [26] ), .QN(_08132_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07706_ ), .Q(\ID_EX_pc [25] ), .QN(_08133_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07706_ ), .Q(\ID_EX_pc [24] ), .QN(_08134_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07706_ ), .Q(\ID_EX_pc [23] ), .QN(_08135_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07706_ ), .Q(\ID_EX_pc [22] ), .QN(_07801_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00206_ ), .CK(_07705_ ), .Q(\ID_EX_rd [4] ), .QN(_07800_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00207_ ), .CK(_07705_ ), .Q(\ID_EX_rd [3] ), .QN(_07799_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00208_ ), .CK(_07705_ ), .Q(\ID_EX_rd [2] ), .QN(_07798_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00209_ ), .CK(_07705_ ), .Q(\ID_EX_rd [1] ), .QN(_07797_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00210_ ), .CK(_07705_ ), .Q(\ID_EX_rd [0] ), .QN(_07796_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00211_ ), .CK(_07704_ ), .Q(\ID_EX_rs1 [4] ), .QN(_07795_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00212_ ), .CK(_07704_ ), .Q(\ID_EX_rs1 [3] ), .QN(_07794_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00214_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_07792_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00213_ ), .CK(_07704_ ), .Q(\ID_EX_rs1 [2] ), .QN(_07793_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00216_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_07790_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00215_ ), .CK(_07704_ ), .Q(\ID_EX_rs1 [1] ), .QN(_07791_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00218_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_07788_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00217_ ), .CK(_07704_ ), .Q(\ID_EX_rs1 [0] ), .QN(_07789_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00220_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_07786_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00219_ ), .CK(_07703_ ), .Q(\ID_EX_rs2 [4] ), .QN(_07787_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00221_ ), .CK(_07703_ ), .Q(\ID_EX_rs2 [3] ), .QN(_07785_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00223_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_07783_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00222_ ), .CK(_07703_ ), .Q(\ID_EX_rs2 [2] ), .QN(_07784_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00225_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_07781_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00224_ ), .CK(_07703_ ), .Q(\ID_EX_rs2 [1] ), .QN(_07782_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00227_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_07779_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00226_ ), .CK(_07703_ ), .Q(\ID_EX_rs2 [0] ), .QN(_07780_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00229_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_07777_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00228_ ), .CK(_07702_ ), .Q(\myidu.stall_quest_fencei ), .QN(_07778_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00230_ ), .CK(_07701_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_07776_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08136_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_ANDNOT__A_Y_$_OR__A_B ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_07700_ ), .Q(\ID_EX_typ [7] ), .QN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00232_ ), .CK(_07700_ ), .Q(\ID_EX_typ [6] ), .QN(_07775_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00233_ ), .CK(_07700_ ), .Q(\ID_EX_typ [5] ), .QN(_07774_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00234_ ), .CK(_07700_ ), .Q(\ID_EX_typ [4] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00235_ ), .CK(_07700_ ), .Q(\ID_EX_typ [3] ), .QN(_07773_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00236_ ), .CK(_07700_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00237_ ), .CK(_07700_ ), .Q(\ID_EX_typ [1] ), .QN(_07772_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00238_ ), .CK(_07700_ ), .Q(\ID_EX_typ [0] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_07699_ ), .Q(check_assert ), .QN(_08137_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.inst_$_DFFE_PP__Q_D ), .CK(_07698_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.inst_$_DFFE_PP__Q_1_D ), .CK(_07698_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.inst_$_DFFE_PP__Q_10_D ), .CK(_07698_ ), .Q(\IF_ID_inst [21] ), .QN(_08138_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.inst_$_DFFE_PP__Q_11_D ), .CK(_07698_ ), .Q(\IF_ID_inst [20] ), .QN(_08139_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.inst_$_DFFE_PP__Q_12_D ), .CK(_07698_ ), .Q(\IF_ID_inst [19] ), .QN(_08140_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.inst_$_DFFE_PP__Q_13_D ), .CK(_07698_ ), .Q(\IF_ID_inst [18] ), .QN(_08141_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.inst_$_DFFE_PP__Q_14_D ), .CK(_07698_ ), .Q(\IF_ID_inst [17] ), .QN(_08142_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.inst_$_DFFE_PP__Q_15_D ), .CK(_07698_ ), .Q(\IF_ID_inst [16] ), .QN(_08143_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.inst_$_DFFE_PP__Q_16_D ), .CK(_07698_ ), .Q(\IF_ID_inst [15] ), .QN(_08144_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.inst_$_DFFE_PP__Q_17_D ), .CK(_07698_ ), .Q(\IF_ID_inst [14] ), .QN(_08145_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.inst_$_DFFE_PP__Q_18_D ), .CK(_07698_ ), .Q(\IF_ID_inst [13] ), .QN(_08146_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.inst_$_DFFE_PP__Q_19_D ), .CK(_07698_ ), .Q(\IF_ID_inst [12] ), .QN(_08147_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.inst_$_DFFE_PP__Q_2_D ), .CK(_07698_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.inst_$_DFFE_PP__Q_20_D ), .CK(_07698_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.inst_$_DFFE_PP__Q_21_D ), .CK(_07698_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.inst_$_DFFE_PP__Q_22_D ), .CK(_07698_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.inst_$_DFFE_PP__Q_23_D ), .CK(_07698_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.inst_$_DFFE_PP__Q_24_D ), .CK(_07698_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.inst_$_DFFE_PP__Q_25_D ), .CK(_07698_ ), .Q(\IF_ID_inst [6] ), .QN(_08148_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.inst_$_DFFE_PP__Q_26_D ), .CK(_07698_ ), .Q(\IF_ID_inst [5] ), .QN(_08149_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.inst_$_DFFE_PP__Q_27_D ), .CK(_07698_ ), .Q(\IF_ID_inst [4] ), .QN(_08150_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.inst_$_DFFE_PP__Q_28_D ), .CK(_07698_ ), .Q(\IF_ID_inst [3] ), .QN(_08151_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.inst_$_DFFE_PP__Q_29_D ), .CK(_07698_ ), .Q(\IF_ID_inst [2] ), .QN(_08152_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.inst_$_DFFE_PP__Q_3_D ), .CK(_07698_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.inst_$_DFFE_PP__Q_30_D ), .CK(_07698_ ), .Q(\IF_ID_inst [1] ), .QN(_08153_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.inst_$_DFFE_PP__Q_31_D ), .CK(_07698_ ), .Q(\IF_ID_inst [0] ), .QN(_08154_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.inst_$_DFFE_PP__Q_4_D ), .CK(_07698_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.inst_$_DFFE_PP__Q_5_D ), .CK(_07698_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.inst_$_DFFE_PP__Q_6_D ), .CK(_07698_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.inst_$_DFFE_PP__Q_7_D ), .CK(_07698_ ), .Q(\IF_ID_inst [24] ), .QN(_08155_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.inst_$_DFFE_PP__Q_8_D ), .CK(_07698_ ), .Q(\IF_ID_inst [23] ), .QN(_08156_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.inst_$_DFFE_PP__Q_9_D ), .CK(_07698_ ), .Q(\IF_ID_inst [22] ), .QN(_08157_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08158_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08159_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08160_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08161_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08162_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08163_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08164_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08165_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08166_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08167_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08168_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08169_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08170_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08171_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08172_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08173_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08174_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08175_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08176_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08177_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08178_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08179_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08180_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08181_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08182_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08183_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08184_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08185_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08186_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08187_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08188_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07697_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08189_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08190_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08191_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08192_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08193_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08194_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08195_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08196_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08197_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08198_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08199_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08200_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08201_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08202_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08203_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08204_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08205_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08206_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08207_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08208_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08209_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08210_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08211_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08212_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08213_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08214_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08215_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08216_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08217_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08218_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08219_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08220_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07696_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08221_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08222_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08223_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08224_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08225_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08226_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08227_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08228_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08229_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08230_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08231_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08232_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08233_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08234_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08235_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08236_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08237_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08238_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08239_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08240_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08241_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08242_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08243_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08244_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08245_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08246_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08247_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08248_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08249_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08250_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08251_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08252_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07695_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08253_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08254_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08255_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08256_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08257_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08258_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08259_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08260_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08261_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08262_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08263_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08264_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08265_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08266_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08267_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08268_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08269_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08270_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08271_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08272_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08273_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08274_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08275_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08276_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08277_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08278_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08279_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08280_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08281_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08282_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08283_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08284_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07694_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08285_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08286_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08287_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08288_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08289_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08290_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08291_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08292_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08293_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08294_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08295_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08296_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08297_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08298_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08299_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08300_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08301_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08302_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08303_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08304_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08305_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08306_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08307_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08308_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08309_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08310_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08311_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08312_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08313_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08314_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08315_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08316_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07693_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08317_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08318_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08319_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08320_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08321_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08322_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08323_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08324_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08325_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08326_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08327_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08328_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08329_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08330_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08331_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08332_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08333_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08334_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08335_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08336_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08337_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08338_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08339_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08340_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08341_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08342_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08343_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08344_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08345_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08346_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08347_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08348_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07692_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08349_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08350_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08351_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08352_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08353_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08354_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08355_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08356_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08357_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08358_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08359_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08360_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08361_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08362_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08363_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08364_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08365_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08366_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08367_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08368_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08369_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08370_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08371_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08372_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08373_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08374_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08375_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08376_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08377_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08378_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08379_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08380_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07691_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08381_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08382_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08383_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08384_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08385_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08386_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08387_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08388_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08389_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08390_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08391_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08392_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08393_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08394_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08395_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08396_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08397_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08398_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08399_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08400_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08401_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08402_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08403_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08404_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08405_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08406_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08407_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08408_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08409_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08410_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08411_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08412_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07690_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08413_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08414_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08415_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08416_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08417_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08418_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08419_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08420_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08421_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08422_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08423_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08424_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08425_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08426_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08427_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08428_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08429_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08430_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08431_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08432_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08433_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08434_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08435_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08436_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08437_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08438_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08439_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07689_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08440_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08441_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08442_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08443_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08444_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08445_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08446_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08447_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08448_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08449_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08450_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08451_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08452_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08453_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08454_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08455_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08456_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08457_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08458_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08459_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08460_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08461_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08462_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08463_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08464_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08465_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08466_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07688_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08467_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08468_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08469_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08470_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08471_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08472_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08473_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08474_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08475_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08476_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08477_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08478_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08479_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08480_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08481_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08482_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08483_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08484_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08485_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08486_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08487_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08488_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08489_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08490_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08491_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08492_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08493_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07687_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08494_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08495_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08496_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08497_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08498_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08499_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08500_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08501_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08502_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08503_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08504_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08505_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08506_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08507_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08508_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08509_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08510_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08511_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08512_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08513_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08514_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08515_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08516_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08517_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08518_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08519_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08520_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07686_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_07771_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00239_ ), .CK(_07685_ ), .Q(\myifu.myicache.valid [0] ), .QN(_07770_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00240_ ), .CK(_07684_ ), .Q(\myifu.myicache.valid [1] ), .QN(_07769_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00241_ ), .CK(_07683_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08521_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_07682_ ), .Q(\myifu.myicache.valid [3] ), .QN(_07768_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00242_ ), .CK(_07681_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00243_ ), .CK(_07680_ ), .Q(\IF_ID_pc [30] ), .QN(_07767_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00244_ ), .CK(_07680_ ), .Q(\IF_ID_pc [21] ), .QN(_07766_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00245_ ), .CK(_07680_ ), .Q(\IF_ID_pc [20] ), .QN(_07765_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00246_ ), .CK(_07680_ ), .Q(\IF_ID_pc [19] ), .QN(_07764_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00247_ ), .CK(_07680_ ), .Q(\IF_ID_pc [18] ), .QN(_07763_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00248_ ), .CK(_07680_ ), .Q(\IF_ID_pc [17] ), .QN(_07762_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00249_ ), .CK(_07680_ ), .Q(\IF_ID_pc [16] ), .QN(_07761_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00250_ ), .CK(_07680_ ), .Q(\IF_ID_pc [15] ), .QN(_07760_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00251_ ), .CK(_07680_ ), .Q(\IF_ID_pc [14] ), .QN(_07759_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00252_ ), .CK(_07680_ ), .Q(\IF_ID_pc [13] ), .QN(_07758_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00253_ ), .CK(_07680_ ), .Q(\IF_ID_pc [12] ), .QN(_07757_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00254_ ), .CK(_07680_ ), .Q(\IF_ID_pc [29] ), .QN(_07756_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00255_ ), .CK(_07680_ ), .Q(\IF_ID_pc [11] ), .QN(_07755_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00256_ ), .CK(_07680_ ), .Q(\IF_ID_pc [10] ), .QN(_07754_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00257_ ), .CK(_07680_ ), .Q(\IF_ID_pc [9] ), .QN(_07753_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00258_ ), .CK(_07680_ ), .Q(\IF_ID_pc [8] ), .QN(_07752_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00259_ ), .CK(_07680_ ), .Q(\IF_ID_pc [7] ), .QN(_07751_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00260_ ), .CK(_07680_ ), .Q(\IF_ID_pc [6] ), .QN(_07750_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00261_ ), .CK(_07680_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00262_ ), .CK(_07680_ ), .Q(\IF_ID_pc [4] ), .QN(_07749_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00264_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_07748_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00263_ ), .CK(_07680_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00266_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_07746_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00265_ ), .CK(_07680_ ), .Q(\IF_ID_pc [2] ), .QN(_07747_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00267_ ), .CK(_07680_ ), .Q(\IF_ID_pc [28] ), .QN(_07745_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00268_ ), .CK(_07680_ ), .Q(\IF_ID_pc [1] ), .QN(_07744_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00269_ ), .CK(_07680_ ), .Q(\IF_ID_pc [27] ), .QN(_07743_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00270_ ), .CK(_07680_ ), .Q(\IF_ID_pc [26] ), .QN(_07742_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00271_ ), .CK(_07680_ ), .Q(\IF_ID_pc [25] ), .QN(_07741_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00272_ ), .CK(_07680_ ), .Q(\IF_ID_pc [24] ), .QN(_07740_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00273_ ), .CK(_07680_ ), .Q(\IF_ID_pc [23] ), .QN(_07739_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00274_ ), .CK(_07680_ ), .Q(\IF_ID_pc [22] ), .QN(_07738_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00275_ ), .CK(_07680_ ), .Q(\IF_ID_pc [31] ), .QN(_07737_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(\myifu.wen_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08523_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_07736_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00276_ ), .CK(_07679_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08522_ ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00277_ ), .CK(_07678_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08524_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08525_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08526_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08527_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08528_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08529_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08530_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08531_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08532_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08533_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08534_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08535_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08536_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08537_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08538_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08539_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08540_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08541_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08542_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08543_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08544_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08545_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08546_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08547_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08548_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08549_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08550_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08551_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08552_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08553_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08554_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08555_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07677_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08556_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08557_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08558_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08559_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08560_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08561_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08562_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08563_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08564_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08565_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08566_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08567_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08568_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08569_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08570_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08571_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08572_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08573_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08574_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08575_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08576_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08577_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08578_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08579_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08580_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08581_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08582_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08583_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08584_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08585_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08586_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08587_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07676_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_07735_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PP0P__Q ( .D(_00278_ ), .CK(_07675_ ), .Q(LS_WB_pc ), .QN(_07734_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PP0P__Q ( .D(_00279_ ), .CK(_07674_ ), .Q(\mylsu.previous_load_done ), .QN(_08588_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08589_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08590_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08591_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(_08592_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_07677_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_07677_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08593_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_07677_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_07733_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00280_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_07732_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00281_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_07731_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00282_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_07730_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00283_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_07729_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00284_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_07728_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00285_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_07727_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00286_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_07726_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00287_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_07725_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00288_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_07724_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00289_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_07723_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00290_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_07722_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00291_ ), .CK(_07673_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08594_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_07677_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08595_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_07677_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08596_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_07677_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08597_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_07677_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08598_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08599_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08600_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08601_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08602_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08603_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08604_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08605_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08606_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08607_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08608_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08609_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08610_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08611_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08612_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08613_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08614_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08615_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08616_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08617_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08618_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08619_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08620_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08621_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08622_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08623_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08624_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08625_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08626_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08627_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08628_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08629_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_07673_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08630_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08631_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_08632_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_08633_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_08634_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_08635_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_08636_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_08637_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_08638_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_08639_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_08640_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_08641_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_08642_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_08643_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_08644_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_08645_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_08646_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_08647_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_08648_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_08649_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_08650_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_08651_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_08652_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_08653_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_08654_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_08655_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_08656_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_08657_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_08658_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_08659_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_08660_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_08661_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_07672_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_07721_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q ( .D(_00292_ ), .CK(_07671_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_07720_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_1 ( .D(_00293_ ), .CK(_07671_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_07719_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_2 ( .D(_00294_ ), .CK(_07671_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_07718_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PP0P__Q ( .D(_00295_ ), .CK(_07671_ ), .Q(LS_WB_wen_reg ), .QN(_08662_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_08663_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_08664_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07670_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07669_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07668_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07667_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07666_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07665_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07664_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07663_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07662_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07661_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07660_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07659_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07658_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07657_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07656_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07655_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00296_ ), .CK(_07654_ ), .Q(loaduse_clear ), .QN(_08665_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_08666_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_08667_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_07717_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(reset ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\ID_EX_typ [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myifu.state [2] ), .Z(fanout_net_39 ) );

endmodule
