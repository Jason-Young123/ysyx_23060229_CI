//Generate the verilog at 2025-09-29T17:45:55 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire _09036_ ;
wire _09037_ ;
wire _09038_ ;
wire _09039_ ;
wire _09040_ ;
wire _09041_ ;
wire _09042_ ;
wire _09043_ ;
wire _09044_ ;
wire _09045_ ;
wire _09046_ ;
wire _09047_ ;
wire _09048_ ;
wire _09049_ ;
wire _09050_ ;
wire _09051_ ;
wire _09052_ ;
wire _09053_ ;
wire _09054_ ;
wire _09055_ ;
wire _09056_ ;
wire _09057_ ;
wire _09058_ ;
wire _09059_ ;
wire _09060_ ;
wire _09061_ ;
wire _09062_ ;
wire _09063_ ;
wire _09064_ ;
wire _09065_ ;
wire _09066_ ;
wire _09067_ ;
wire _09068_ ;
wire _09069_ ;
wire _09070_ ;
wire _09071_ ;
wire _09072_ ;
wire _09073_ ;
wire _09074_ ;
wire _09075_ ;
wire _09076_ ;
wire _09077_ ;
wire _09078_ ;
wire _09079_ ;
wire _09080_ ;
wire _09081_ ;
wire _09082_ ;
wire _09083_ ;
wire _09084_ ;
wire _09085_ ;
wire _09086_ ;
wire _09087_ ;
wire _09088_ ;
wire _09089_ ;
wire _09090_ ;
wire _09091_ ;
wire _09092_ ;
wire _09093_ ;
wire _09094_ ;
wire _09095_ ;
wire _09096_ ;
wire _09097_ ;
wire _09098_ ;
wire _09099_ ;
wire _09100_ ;
wire _09101_ ;
wire _09102_ ;
wire _09103_ ;
wire _09104_ ;
wire _09105_ ;
wire _09106_ ;
wire _09107_ ;
wire _09108_ ;
wire _09109_ ;
wire _09110_ ;
wire _09111_ ;
wire _09112_ ;
wire _09113_ ;
wire _09114_ ;
wire _09115_ ;
wire _09116_ ;
wire _09117_ ;
wire _09118_ ;
wire _09119_ ;
wire _09120_ ;
wire _09121_ ;
wire _09122_ ;
wire _09123_ ;
wire _09124_ ;
wire _09125_ ;
wire _09126_ ;
wire _09127_ ;
wire _09128_ ;
wire _09129_ ;
wire _09130_ ;
wire _09131_ ;
wire _09132_ ;
wire _09133_ ;
wire _09134_ ;
wire _09135_ ;
wire _09136_ ;
wire _09137_ ;
wire _09138_ ;
wire _09139_ ;
wire _09140_ ;
wire _09141_ ;
wire _09142_ ;
wire _09143_ ;
wire _09144_ ;
wire _09145_ ;
wire _09146_ ;
wire _09147_ ;
wire _09148_ ;
wire _09149_ ;
wire _09150_ ;
wire _09151_ ;
wire _09152_ ;
wire _09153_ ;
wire _09154_ ;
wire _09155_ ;
wire _09156_ ;
wire _09157_ ;
wire _09158_ ;
wire _09159_ ;
wire _09160_ ;
wire _09161_ ;
wire _09162_ ;
wire _09163_ ;
wire _09164_ ;
wire _09165_ ;
wire _09166_ ;
wire _09167_ ;
wire _09168_ ;
wire _09169_ ;
wire _09170_ ;
wire _09171_ ;
wire _09172_ ;
wire _09173_ ;
wire _09174_ ;
wire _09175_ ;
wire _09176_ ;
wire _09177_ ;
wire _09178_ ;
wire _09179_ ;
wire _09180_ ;
wire _09181_ ;
wire _09182_ ;
wire _09183_ ;
wire _09184_ ;
wire _09185_ ;
wire _09186_ ;
wire _09187_ ;
wire _09188_ ;
wire _09189_ ;
wire _09190_ ;
wire _09191_ ;
wire _09192_ ;
wire _09193_ ;
wire _09194_ ;
wire _09195_ ;
wire _09196_ ;
wire _09197_ ;
wire _09198_ ;
wire _09199_ ;
wire _09200_ ;
wire _09201_ ;
wire _09202_ ;
wire _09203_ ;
wire _09204_ ;
wire _09205_ ;
wire _09206_ ;
wire _09207_ ;
wire _09208_ ;
wire _09209_ ;
wire _09210_ ;
wire _09211_ ;
wire _09212_ ;
wire _09213_ ;
wire _09214_ ;
wire _09215_ ;
wire _09216_ ;
wire _09217_ ;
wire _09218_ ;
wire _09219_ ;
wire _09220_ ;
wire _09221_ ;
wire _09222_ ;
wire _09223_ ;
wire _09224_ ;
wire _09225_ ;
wire _09226_ ;
wire _09227_ ;
wire _09228_ ;
wire _09229_ ;
wire _09230_ ;
wire _09231_ ;
wire _09232_ ;
wire _09233_ ;
wire _09234_ ;
wire _09235_ ;
wire _09236_ ;
wire _09237_ ;
wire _09238_ ;
wire _09239_ ;
wire _09240_ ;
wire _09241_ ;
wire _09242_ ;
wire _09243_ ;
wire _09244_ ;
wire _09245_ ;
wire _09246_ ;
wire _09247_ ;
wire _09248_ ;
wire _09249_ ;
wire _09250_ ;
wire _09251_ ;
wire _09252_ ;
wire _09253_ ;
wire _09254_ ;
wire _09255_ ;
wire _09256_ ;
wire _09257_ ;
wire _09258_ ;
wire _09259_ ;
wire _09260_ ;
wire _09261_ ;
wire _09262_ ;
wire _09263_ ;
wire _09264_ ;
wire _09265_ ;
wire _09266_ ;
wire _09267_ ;
wire _09268_ ;
wire _09269_ ;
wire _09270_ ;
wire _09271_ ;
wire _09272_ ;
wire _09273_ ;
wire _09274_ ;
wire _09275_ ;
wire _09276_ ;
wire _09277_ ;
wire _09278_ ;
wire _09279_ ;
wire _09280_ ;
wire _09281_ ;
wire _09282_ ;
wire _09283_ ;
wire _09284_ ;
wire _09285_ ;
wire _09286_ ;
wire _09287_ ;
wire _09288_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFF_PP0__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire \myexu.pc_out_$_SDFFE_PP0P__Q_E ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_ANDNOT__A_Y ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

INV_X2 _09289_ ( .A(fanout_net_1 ), .ZN(_01773_ ) );
BUF_X4 _09290_ ( .A(_01773_ ), .Z(_01774_ ) );
AND3_X4 _09291_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01775_ ) );
AND3_X4 _09292_ ( .A1(_01775_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01776_ ) );
AND3_X4 _09293_ ( .A1(_01776_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01777_ ) );
AND2_X4 _09294_ ( .A1(_01777_ ), .A2(\myclint.mtime [7] ), .ZN(_01778_ ) );
AND2_X1 _09295_ ( .A1(\myclint.mtime [8] ), .A2(\myclint.mtime [9] ), .ZN(_01779_ ) );
AND3_X4 _09296_ ( .A1(_01778_ ), .A2(\myclint.mtime [10] ), .A3(_01779_ ), .ZN(_01780_ ) );
AND3_X4 _09297_ ( .A1(_01780_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01781_ ) );
AND3_X4 _09298_ ( .A1(_01781_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01782_ ) );
AND3_X4 _09299_ ( .A1(_01782_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01783_ ) );
AND3_X4 _09300_ ( .A1(_01783_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01784_ ) );
AND3_X4 _09301_ ( .A1(_01784_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01785_ ) );
AND3_X4 _09302_ ( .A1(_01785_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01786_ ) );
AND3_X4 _09303_ ( .A1(_01786_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01787_ ) );
AND3_X4 _09304_ ( .A1(_01787_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01788_ ) );
AND2_X4 _09305_ ( .A1(_01788_ ), .A2(\myclint.mtime [27] ), .ZN(_01789_ ) );
AND2_X1 _09306_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01790_ ) );
AND2_X1 _09307_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01791_ ) );
NAND4_X4 _09308_ ( .A1(_01789_ ), .A2(\myclint.mtime [33] ), .A3(_01790_ ), .A4(_01791_ ), .ZN(_01792_ ) );
INV_X1 _09309_ ( .A(\myclint.mtime [32] ), .ZN(_01793_ ) );
NOR2_X2 _09310_ ( .A1(_01792_ ), .A2(_01793_ ), .ZN(_01794_ ) );
NAND3_X1 _09311_ ( .A1(_01794_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01795_ ) );
INV_X1 _09312_ ( .A(\myclint.mtime [36] ), .ZN(_01796_ ) );
INV_X1 _09313_ ( .A(\myclint.mtime [37] ), .ZN(_01797_ ) );
NOR3_X2 _09314_ ( .A1(_01795_ ), .A2(_01796_ ), .A3(_01797_ ), .ZN(_01798_ ) );
NAND3_X1 _09315_ ( .A1(_01798_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [39] ), .ZN(_01799_ ) );
INV_X1 _09316_ ( .A(\myclint.mtime [40] ), .ZN(_01800_ ) );
NOR2_X1 _09317_ ( .A1(_01799_ ), .A2(_01800_ ), .ZN(_01801_ ) );
AND3_X2 _09318_ ( .A1(_01801_ ), .A2(\myclint.mtime [42] ), .A3(\myclint.mtime [41] ), .ZN(_01802_ ) );
AND2_X1 _09319_ ( .A1(_01802_ ), .A2(\myclint.mtime [43] ), .ZN(_01803_ ) );
AND2_X1 _09320_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01804_ ) );
AND2_X2 _09321_ ( .A1(_01803_ ), .A2(_01804_ ), .ZN(_01805_ ) );
AND2_X1 _09322_ ( .A1(\myclint.mtime [46] ), .A2(\myclint.mtime [47] ), .ZN(_01806_ ) );
NAND2_X1 _09323_ ( .A1(_01805_ ), .A2(_01806_ ), .ZN(_01807_ ) );
AND2_X1 _09324_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01808_ ) );
INV_X1 _09325_ ( .A(_01808_ ), .ZN(_01809_ ) );
NOR2_X1 _09326_ ( .A1(_01807_ ), .A2(_01809_ ), .ZN(_01810_ ) );
AND2_X1 _09327_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01811_ ) );
NAND2_X1 _09328_ ( .A1(_01810_ ), .A2(_01811_ ), .ZN(_01812_ ) );
AND2_X1 _09329_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01813_ ) );
INV_X1 _09330_ ( .A(_01813_ ), .ZN(_01814_ ) );
NOR2_X1 _09331_ ( .A1(_01812_ ), .A2(_01814_ ), .ZN(_01815_ ) );
AND2_X1 _09332_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01816_ ) );
NAND2_X1 _09333_ ( .A1(_01815_ ), .A2(_01816_ ), .ZN(_01817_ ) );
AND2_X1 _09334_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01818_ ) );
INV_X1 _09335_ ( .A(_01818_ ), .ZN(_01819_ ) );
NOR2_X1 _09336_ ( .A1(_01817_ ), .A2(_01819_ ), .ZN(_01820_ ) );
AND2_X1 _09337_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01821_ ) );
AND2_X1 _09338_ ( .A1(_01820_ ), .A2(_01821_ ), .ZN(_01822_ ) );
NAND3_X1 _09339_ ( .A1(_01822_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01823_ ) );
NOR2_X1 _09340_ ( .A1(_01823_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01824_ ) );
OAI21_X1 _09341_ ( .A(_01774_ ), .B1(_01824_ ), .B2(\myclint.mtime [63] ), .ZN(_01825_ ) );
AND2_X4 _09342_ ( .A1(_01789_ ), .A2(_01791_ ), .ZN(_01826_ ) );
AND2_X1 _09343_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01827_ ) );
AND3_X4 _09344_ ( .A1(_01826_ ), .A2(_01827_ ), .A3(_01790_ ), .ZN(_01828_ ) );
NAND2_X2 _09345_ ( .A1(_01828_ ), .A2(\myclint.mtime [34] ), .ZN(_01829_ ) );
INV_X1 _09346_ ( .A(\myclint.mtime [35] ), .ZN(_01830_ ) );
NOR3_X2 _09347_ ( .A1(_01829_ ), .A2(_01796_ ), .A3(_01830_ ), .ZN(_01831_ ) );
AND3_X2 _09348_ ( .A1(_01831_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [37] ), .ZN(_01832_ ) );
AND3_X2 _09349_ ( .A1(_01832_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [39] ), .ZN(_01833_ ) );
AND3_X2 _09350_ ( .A1(_01833_ ), .A2(\myclint.mtime [42] ), .A3(\myclint.mtime [41] ), .ZN(_01834_ ) );
AND2_X2 _09351_ ( .A1(_01834_ ), .A2(\myclint.mtime [43] ), .ZN(_01835_ ) );
AND2_X2 _09352_ ( .A1(_01835_ ), .A2(_01804_ ), .ZN(_01836_ ) );
AND2_X4 _09353_ ( .A1(_01836_ ), .A2(_01806_ ), .ZN(_01837_ ) );
AND2_X2 _09354_ ( .A1(_01837_ ), .A2(_01808_ ), .ZN(_01838_ ) );
AND2_X4 _09355_ ( .A1(_01838_ ), .A2(_01811_ ), .ZN(_01839_ ) );
AND2_X4 _09356_ ( .A1(_01839_ ), .A2(_01813_ ), .ZN(_01840_ ) );
AND2_X4 _09357_ ( .A1(_01840_ ), .A2(_01816_ ), .ZN(_01841_ ) );
AND2_X4 _09358_ ( .A1(_01841_ ), .A2(_01818_ ), .ZN(_01842_ ) );
AND2_X2 _09359_ ( .A1(_01842_ ), .A2(_01821_ ), .ZN(_01843_ ) );
NAND3_X1 _09360_ ( .A1(_01843_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01844_ ) );
NOR2_X1 _09361_ ( .A1(_01844_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01845_ ) );
AOI21_X1 _09362_ ( .A(_01825_ ), .B1(_01845_ ), .B2(\myclint.mtime [63] ), .ZN(_00000_ ) );
AND4_X1 _09363_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01846_ ) );
AND4_X1 _09364_ ( .A1(\myclint.mtime [10] ), .A2(_01846_ ), .A3(\myclint.mtime [11] ), .A4(_01779_ ), .ZN(_01847_ ) );
NAND2_X1 _09365_ ( .A1(_01778_ ), .A2(_01847_ ), .ZN(_01848_ ) );
AND2_X1 _09366_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_01849_ ) );
NAND3_X1 _09367_ ( .A1(_01849_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01850_ ) );
NAND4_X1 _09368_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01851_ ) );
NOR2_X1 _09369_ ( .A1(_01850_ ), .A2(_01851_ ), .ZN(_01852_ ) );
AND2_X1 _09370_ ( .A1(\myclint.mtime [24] ), .A2(\myclint.mtime [25] ), .ZN(_01853_ ) );
AND3_X1 _09371_ ( .A1(_01853_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [27] ), .ZN(_01854_ ) );
NAND4_X1 _09372_ ( .A1(_01852_ ), .A2(_01790_ ), .A3(_01791_ ), .A4(_01854_ ), .ZN(_01855_ ) );
NOR2_X1 _09373_ ( .A1(_01848_ ), .A2(_01855_ ), .ZN(_01856_ ) );
NAND3_X1 _09374_ ( .A1(_01827_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01857_ ) );
NAND4_X1 _09375_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01858_ ) );
NOR2_X1 _09376_ ( .A1(_01857_ ), .A2(_01858_ ), .ZN(_01859_ ) );
AND2_X1 _09377_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01860_ ) );
AND3_X1 _09378_ ( .A1(_01860_ ), .A2(\myclint.mtime [42] ), .A3(\myclint.mtime [43] ), .ZN(_01861_ ) );
AND4_X1 _09379_ ( .A1(_01806_ ), .A2(_01859_ ), .A3(_01804_ ), .A4(_01861_ ), .ZN(_01862_ ) );
NAND2_X1 _09380_ ( .A1(_01856_ ), .A2(_01862_ ), .ZN(_01863_ ) );
INV_X1 _09381_ ( .A(_01863_ ), .ZN(_01864_ ) );
AND4_X1 _09382_ ( .A1(_01816_ ), .A2(_01813_ ), .A3(_01811_ ), .A4(_01808_ ), .ZN(_01865_ ) );
AND2_X1 _09383_ ( .A1(_01864_ ), .A2(_01865_ ), .ZN(_01866_ ) );
AND4_X1 _09384_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01867_ ) );
AND2_X1 _09385_ ( .A1(_01866_ ), .A2(_01867_ ), .ZN(_01868_ ) );
AND3_X1 _09386_ ( .A1(_01868_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01869_ ) );
XNOR2_X1 _09387_ ( .A(_01869_ ), .B(\myclint.mtime [62] ), .ZN(_01870_ ) );
NOR2_X1 _09388_ ( .A1(_01870_ ), .A2(fanout_net_1 ), .ZN(_00001_ ) );
AND2_X1 _09389_ ( .A1(_01811_ ), .A2(_01808_ ), .ZN(_01871_ ) );
INV_X1 _09390_ ( .A(_01871_ ), .ZN(_01872_ ) );
NOR3_X1 _09391_ ( .A1(_01863_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01872_ ), .ZN(_01873_ ) );
XNOR2_X1 _09392_ ( .A(_01873_ ), .B(\myclint.mtime [53] ), .ZN(_01874_ ) );
NOR2_X1 _09393_ ( .A1(_01874_ ), .A2(fanout_net_1 ), .ZN(_00002_ ) );
OR3_X1 _09394_ ( .A1(_01863_ ), .A2(\myclint.mtime [52] ), .A3(_01872_ ), .ZN(_01875_ ) );
OAI21_X1 _09395_ ( .A(\myclint.mtime [52] ), .B1(_01863_ ), .B2(_01872_ ), .ZN(_01876_ ) );
AOI21_X1 _09396_ ( .A(fanout_net_1 ), .B1(_01875_ ), .B2(_01876_ ), .ZN(_00003_ ) );
NOR3_X1 _09397_ ( .A1(_01807_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01809_ ), .ZN(_01877_ ) );
OAI21_X1 _09398_ ( .A(_01774_ ), .B1(_01877_ ), .B2(\myclint.mtime [51] ), .ZN(_01878_ ) );
INV_X1 _09399_ ( .A(_01837_ ), .ZN(_01879_ ) );
NOR3_X1 _09400_ ( .A1(_01879_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01809_ ), .ZN(_01880_ ) );
AOI21_X1 _09401_ ( .A(_01878_ ), .B1(_01880_ ), .B2(\myclint.mtime [51] ), .ZN(_00004_ ) );
NAND3_X1 _09402_ ( .A1(_01856_ ), .A2(_01808_ ), .A3(_01862_ ), .ZN(_01881_ ) );
OR2_X1 _09403_ ( .A1(_01881_ ), .A2(\myclint.mtime [50] ), .ZN(_01882_ ) );
NAND2_X1 _09404_ ( .A1(_01881_ ), .A2(\myclint.mtime [50] ), .ZN(_01883_ ) );
AOI21_X1 _09405_ ( .A(fanout_net_1 ), .B1(_01882_ ), .B2(_01883_ ), .ZN(_00005_ ) );
INV_X1 _09406_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01884_ ) );
AND4_X1 _09407_ ( .A1(\myclint.mtime [49] ), .A2(_01836_ ), .A3(_01884_ ), .A4(_01806_ ), .ZN(_01885_ ) );
BUF_X4 _09408_ ( .A(_01773_ ), .Z(_01886_ ) );
BUF_X4 _09409_ ( .A(_01886_ ), .Z(_01887_ ) );
AND3_X1 _09410_ ( .A1(_01805_ ), .A2(_01884_ ), .A3(_01806_ ), .ZN(_01888_ ) );
OAI21_X1 _09411_ ( .A(_01887_ ), .B1(_01888_ ), .B2(\myclint.mtime [49] ), .ZN(_01889_ ) );
NOR2_X1 _09412_ ( .A1(_01885_ ), .A2(_01889_ ), .ZN(_00006_ ) );
NAND2_X1 _09413_ ( .A1(_01863_ ), .A2(\myclint.mtime [48] ), .ZN(_01890_ ) );
INV_X1 _09414_ ( .A(_01862_ ), .ZN(_01891_ ) );
OR4_X1 _09415_ ( .A1(\myclint.mtime [48] ), .A2(_01848_ ), .A3(_01855_ ), .A4(_01891_ ), .ZN(_01892_ ) );
AOI21_X1 _09416_ ( .A(fanout_net_1 ), .B1(_01890_ ), .B2(_01892_ ), .ZN(_00007_ ) );
AND2_X1 _09417_ ( .A1(_01856_ ), .A2(_01859_ ), .ZN(_01893_ ) );
NAND3_X1 _09418_ ( .A1(_01893_ ), .A2(_01804_ ), .A3(_01861_ ), .ZN(_01894_ ) );
OR3_X1 _09419_ ( .A1(_01894_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [47] ), .ZN(_01895_ ) );
OAI21_X1 _09420_ ( .A(\myclint.mtime [47] ), .B1(_01894_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01896_ ) );
AOI21_X1 _09421_ ( .A(fanout_net_1 ), .B1(_01895_ ), .B2(_01896_ ), .ZN(_00008_ ) );
OR2_X1 _09422_ ( .A1(_01894_ ), .A2(\myclint.mtime [46] ), .ZN(_01897_ ) );
NAND2_X1 _09423_ ( .A1(_01894_ ), .A2(\myclint.mtime [46] ), .ZN(_01898_ ) );
AOI21_X1 _09424_ ( .A(fanout_net_1 ), .B1(_01897_ ), .B2(_01898_ ), .ZN(_00009_ ) );
NAND2_X1 _09425_ ( .A1(_01802_ ), .A2(\myclint.mtime [43] ), .ZN(_01899_ ) );
NOR2_X1 _09426_ ( .A1(_01899_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01900_ ) );
OAI21_X1 _09427_ ( .A(_01774_ ), .B1(_01900_ ), .B2(\myclint.mtime [45] ), .ZN(_01901_ ) );
INV_X1 _09428_ ( .A(_01834_ ), .ZN(_01902_ ) );
INV_X1 _09429_ ( .A(\myclint.mtime [43] ), .ZN(_01903_ ) );
NOR3_X1 _09430_ ( .A1(_01902_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01903_ ), .ZN(_01904_ ) );
AOI21_X1 _09431_ ( .A(_01901_ ), .B1(_01904_ ), .B2(\myclint.mtime [45] ), .ZN(_00010_ ) );
AND2_X1 _09432_ ( .A1(_01893_ ), .A2(_01861_ ), .ZN(_01905_ ) );
XNOR2_X1 _09433_ ( .A(_01905_ ), .B(\myclint.mtime [44] ), .ZN(_01906_ ) );
NOR2_X1 _09434_ ( .A1(_01906_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
INV_X1 _09435_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01907_ ) );
AND3_X1 _09436_ ( .A1(_01820_ ), .A2(_01907_ ), .A3(_01821_ ), .ZN(_01908_ ) );
OAI21_X1 _09437_ ( .A(_01774_ ), .B1(_01908_ ), .B2(\myclint.mtime [61] ), .ZN(_01909_ ) );
AND3_X1 _09438_ ( .A1(_01842_ ), .A2(_01907_ ), .A3(_01821_ ), .ZN(_01910_ ) );
AOI21_X1 _09439_ ( .A(_01909_ ), .B1(_01910_ ), .B2(\myclint.mtime [61] ), .ZN(_00012_ ) );
NAND3_X1 _09440_ ( .A1(_01856_ ), .A2(_01860_ ), .A3(_01859_ ), .ZN(_01911_ ) );
NOR2_X1 _09441_ ( .A1(_01911_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01912_ ) );
XNOR2_X1 _09442_ ( .A(_01912_ ), .B(\myclint.mtime [43] ), .ZN(_01913_ ) );
NOR2_X1 _09443_ ( .A1(_01913_ ), .A2(fanout_net_1 ), .ZN(_00013_ ) );
CLKBUF_X2 _09444_ ( .A(_01886_ ), .Z(_01914_ ) );
INV_X1 _09445_ ( .A(\myclint.mtime [41] ), .ZN(_01915_ ) );
NOR3_X1 _09446_ ( .A1(_01799_ ), .A2(_01800_ ), .A3(_01915_ ), .ZN(_01916_ ) );
OAI21_X1 _09447_ ( .A(_01914_ ), .B1(_01916_ ), .B2(\myclint.mtime [42] ), .ZN(_01917_ ) );
NOR2_X1 _09448_ ( .A1(_01917_ ), .A2(_01802_ ), .ZN(_00014_ ) );
NOR2_X1 _09449_ ( .A1(_01799_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01918_ ) );
OAI21_X1 _09450_ ( .A(_01774_ ), .B1(_01918_ ), .B2(\myclint.mtime [41] ), .ZN(_01919_ ) );
INV_X1 _09451_ ( .A(_01832_ ), .ZN(_01920_ ) );
INV_X1 _09452_ ( .A(\myclint.mtime [39] ), .ZN(_01921_ ) );
NOR3_X1 _09453_ ( .A1(_01920_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01921_ ), .ZN(_01922_ ) );
AOI21_X1 _09454_ ( .A(_01919_ ), .B1(\myclint.mtime [41] ), .B2(_01922_ ), .ZN(_00015_ ) );
INV_X1 _09455_ ( .A(_01801_ ), .ZN(_01923_ ) );
AOI21_X1 _09456_ ( .A(fanout_net_1 ), .B1(_01799_ ), .B2(_01800_ ), .ZN(_01924_ ) );
AND2_X1 _09457_ ( .A1(_01923_ ), .A2(_01924_ ), .ZN(_00016_ ) );
AND4_X1 _09458_ ( .A1(\myclint.mtime [33] ), .A2(_01789_ ), .A3(_01790_ ), .A4(_01791_ ), .ZN(_01925_ ) );
NAND3_X1 _09459_ ( .A1(_01925_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01926_ ) );
NOR3_X1 _09460_ ( .A1(_01926_ ), .A2(_01796_ ), .A3(_01830_ ), .ZN(_01927_ ) );
INV_X1 _09461_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01928_ ) );
NAND3_X1 _09462_ ( .A1(_01927_ ), .A2(_01928_ ), .A3(\myclint.mtime [37] ), .ZN(_01929_ ) );
AOI21_X1 _09463_ ( .A(fanout_net_1 ), .B1(_01929_ ), .B2(_01921_ ), .ZN(_01930_ ) );
NAND4_X1 _09464_ ( .A1(_01831_ ), .A2(_01928_ ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01931_ ) );
AND2_X1 _09465_ ( .A1(_01930_ ), .A2(_01931_ ), .ZN(_00017_ ) );
OAI21_X1 _09466_ ( .A(_01914_ ), .B1(_01798_ ), .B2(\myclint.mtime [38] ), .ZN(_01932_ ) );
AND3_X1 _09467_ ( .A1(_01927_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [37] ), .ZN(_01933_ ) );
NOR2_X1 _09468_ ( .A1(_01932_ ), .A2(_01933_ ), .ZN(_00018_ ) );
BUF_X4 _09469_ ( .A(_01886_ ), .Z(_01934_ ) );
NOR3_X1 _09470_ ( .A1(_01926_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01830_ ), .ZN(_01935_ ) );
OAI21_X1 _09471_ ( .A(_01934_ ), .B1(_01935_ ), .B2(\myclint.mtime [37] ), .ZN(_01936_ ) );
NOR4_X1 _09472_ ( .A1(_01829_ ), .A2(_01797_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A4(_01830_ ), .ZN(_01937_ ) );
NOR2_X1 _09473_ ( .A1(_01936_ ), .A2(_01937_ ), .ZN(_00019_ ) );
AND3_X1 _09474_ ( .A1(_01794_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01938_ ) );
OAI21_X1 _09475_ ( .A(_01934_ ), .B1(_01938_ ), .B2(\myclint.mtime [36] ), .ZN(_01939_ ) );
NOR2_X1 _09476_ ( .A1(_01939_ ), .A2(_01927_ ), .ZN(_00020_ ) );
INV_X1 _09477_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01940_ ) );
AND3_X1 _09478_ ( .A1(_01828_ ), .A2(_01940_ ), .A3(\myclint.mtime [35] ), .ZN(_01941_ ) );
NOR3_X1 _09479_ ( .A1(_01792_ ), .A2(_01793_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01942_ ) );
OAI21_X1 _09480_ ( .A(_01887_ ), .B1(_01942_ ), .B2(\myclint.mtime [35] ), .ZN(_01943_ ) );
NOR2_X1 _09481_ ( .A1(_01941_ ), .A2(_01943_ ), .ZN(_00021_ ) );
OAI21_X1 _09482_ ( .A(_01934_ ), .B1(_01794_ ), .B2(\myclint.mtime [34] ), .ZN(_01944_ ) );
AND3_X1 _09483_ ( .A1(_01925_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01945_ ) );
NOR2_X1 _09484_ ( .A1(_01944_ ), .A2(_01945_ ), .ZN(_00022_ ) );
XNOR2_X1 _09485_ ( .A(_01868_ ), .B(\myclint.mtime [60] ), .ZN(_01946_ ) );
NOR2_X1 _09486_ ( .A1(_01946_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
INV_X1 _09487_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01947_ ) );
AND3_X1 _09488_ ( .A1(_01826_ ), .A2(_01947_ ), .A3(_01790_ ), .ZN(_01948_ ) );
AND2_X1 _09489_ ( .A1(_01948_ ), .A2(\myclint.mtime [33] ), .ZN(_01949_ ) );
OAI21_X1 _09490_ ( .A(_01887_ ), .B1(_01948_ ), .B2(\myclint.mtime [33] ), .ZN(_01950_ ) );
NOR2_X1 _09491_ ( .A1(_01949_ ), .A2(_01950_ ), .ZN(_00024_ ) );
OAI21_X1 _09492_ ( .A(\myclint.mtime [32] ), .B1(_01848_ ), .B2(_01855_ ), .ZN(_01951_ ) );
AND4_X1 _09493_ ( .A1(_01790_ ), .A2(_01852_ ), .A3(_01791_ ), .A4(_01854_ ), .ZN(_01952_ ) );
NAND4_X1 _09494_ ( .A1(_01778_ ), .A2(_01793_ ), .A3(_01847_ ), .A4(_01952_ ), .ZN(_01953_ ) );
AOI21_X1 _09495_ ( .A(fanout_net_1 ), .B1(_01951_ ), .B2(_01953_ ), .ZN(_00025_ ) );
AND2_X1 _09496_ ( .A1(_01778_ ), .A2(_01847_ ), .ZN(_01954_ ) );
AND2_X1 _09497_ ( .A1(_01954_ ), .A2(_01852_ ), .ZN(_01955_ ) );
NAND3_X1 _09498_ ( .A1(_01955_ ), .A2(_01791_ ), .A3(_01854_ ), .ZN(_01956_ ) );
OR3_X1 _09499_ ( .A1(_01956_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [31] ), .ZN(_01957_ ) );
OAI21_X1 _09500_ ( .A(\myclint.mtime [31] ), .B1(_01956_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01958_ ) );
AOI21_X1 _09501_ ( .A(fanout_net_1 ), .B1(_01957_ ), .B2(_01958_ ), .ZN(_00026_ ) );
OR2_X1 _09502_ ( .A1(_01956_ ), .A2(\myclint.mtime [30] ), .ZN(_01959_ ) );
NAND2_X1 _09503_ ( .A1(_01956_ ), .A2(\myclint.mtime [30] ), .ZN(_01960_ ) );
AOI21_X1 _09504_ ( .A(fanout_net_1 ), .B1(_01959_ ), .B2(_01960_ ), .ZN(_00027_ ) );
INV_X1 _09505_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01961_ ) );
AND3_X1 _09506_ ( .A1(_01788_ ), .A2(_01961_ ), .A3(\myclint.mtime [27] ), .ZN(_01962_ ) );
AND2_X1 _09507_ ( .A1(_01962_ ), .A2(\myclint.mtime [29] ), .ZN(_01963_ ) );
OAI21_X1 _09508_ ( .A(_01887_ ), .B1(_01962_ ), .B2(\myclint.mtime [29] ), .ZN(_01964_ ) );
NOR2_X1 _09509_ ( .A1(_01963_ ), .A2(_01964_ ), .ZN(_00028_ ) );
NAND2_X1 _09510_ ( .A1(_01955_ ), .A2(_01854_ ), .ZN(_01965_ ) );
OR2_X1 _09511_ ( .A1(_01965_ ), .A2(\myclint.mtime [28] ), .ZN(_01966_ ) );
NAND2_X1 _09512_ ( .A1(_01965_ ), .A2(\myclint.mtime [28] ), .ZN(_01967_ ) );
AOI21_X1 _09513_ ( .A(fanout_net_1 ), .B1(_01966_ ), .B2(_01967_ ), .ZN(_00029_ ) );
NAND3_X1 _09514_ ( .A1(_01954_ ), .A2(_01853_ ), .A3(_01852_ ), .ZN(_01968_ ) );
OR3_X1 _09515_ ( .A1(_01968_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01969_ ) );
OAI21_X1 _09516_ ( .A(\myclint.mtime [27] ), .B1(_01968_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01970_ ) );
AOI21_X1 _09517_ ( .A(fanout_net_1 ), .B1(_01969_ ), .B2(_01970_ ), .ZN(_00030_ ) );
AND2_X1 _09518_ ( .A1(_01787_ ), .A2(\myclint.mtime [25] ), .ZN(_01971_ ) );
OAI21_X1 _09519_ ( .A(_01934_ ), .B1(_01971_ ), .B2(\myclint.mtime [26] ), .ZN(_01972_ ) );
NOR2_X1 _09520_ ( .A1(_01972_ ), .A2(_01788_ ), .ZN(_00031_ ) );
INV_X1 _09521_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01973_ ) );
AND3_X1 _09522_ ( .A1(_01786_ ), .A2(_01973_ ), .A3(\myclint.mtime [23] ), .ZN(_01974_ ) );
AND2_X1 _09523_ ( .A1(_01974_ ), .A2(\myclint.mtime [25] ), .ZN(_01975_ ) );
OAI21_X1 _09524_ ( .A(_01774_ ), .B1(_01974_ ), .B2(\myclint.mtime [25] ), .ZN(_01976_ ) );
NOR2_X1 _09525_ ( .A1(_01975_ ), .A2(_01976_ ), .ZN(_00032_ ) );
AND2_X1 _09526_ ( .A1(_01786_ ), .A2(\myclint.mtime [23] ), .ZN(_01977_ ) );
OAI21_X1 _09527_ ( .A(_01934_ ), .B1(_01977_ ), .B2(\myclint.mtime [24] ), .ZN(_01978_ ) );
NOR2_X1 _09528_ ( .A1(_01978_ ), .A2(_01787_ ), .ZN(_00033_ ) );
NOR3_X1 _09529_ ( .A1(_01817_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01819_ ), .ZN(_01979_ ) );
OAI21_X1 _09530_ ( .A(_01774_ ), .B1(_01979_ ), .B2(\myclint.mtime [59] ), .ZN(_01980_ ) );
INV_X1 _09531_ ( .A(_01841_ ), .ZN(_01981_ ) );
NOR3_X1 _09532_ ( .A1(_01981_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01819_ ), .ZN(_01982_ ) );
AOI21_X1 _09533_ ( .A(_01980_ ), .B1(_01982_ ), .B2(\myclint.mtime [59] ), .ZN(_00034_ ) );
NOR2_X1 _09534_ ( .A1(_01848_ ), .A2(_01850_ ), .ZN(_01983_ ) );
NAND3_X1 _09535_ ( .A1(_01983_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01984_ ) );
OR3_X1 _09536_ ( .A1(_01984_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01985_ ) );
OAI21_X1 _09537_ ( .A(\myclint.mtime [23] ), .B1(_01984_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01986_ ) );
AOI21_X1 _09538_ ( .A(fanout_net_1 ), .B1(_01985_ ), .B2(_01986_ ), .ZN(_00035_ ) );
AND2_X1 _09539_ ( .A1(_01785_ ), .A2(\myclint.mtime [21] ), .ZN(_01987_ ) );
OAI21_X1 _09540_ ( .A(_01934_ ), .B1(_01987_ ), .B2(\myclint.mtime [22] ), .ZN(_01988_ ) );
NOR2_X1 _09541_ ( .A1(_01988_ ), .A2(_01786_ ), .ZN(_00036_ ) );
OR3_X1 _09542_ ( .A1(_01848_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01850_ ), .ZN(_01989_ ) );
NAND2_X1 _09543_ ( .A1(_01989_ ), .A2(\myclint.mtime [21] ), .ZN(_01990_ ) );
OR4_X1 _09544_ ( .A1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01848_ ), .A3(\myclint.mtime [21] ), .A4(_01850_ ), .ZN(_01991_ ) );
AOI21_X1 _09545_ ( .A(fanout_net_1 ), .B1(_01990_ ), .B2(_01991_ ), .ZN(_00037_ ) );
AND2_X1 _09546_ ( .A1(_01784_ ), .A2(\myclint.mtime [19] ), .ZN(_01992_ ) );
OAI21_X1 _09547_ ( .A(_01934_ ), .B1(_01992_ ), .B2(\myclint.mtime [20] ), .ZN(_01993_ ) );
NOR2_X1 _09548_ ( .A1(_01993_ ), .A2(_01785_ ), .ZN(_00038_ ) );
NAND3_X1 _09549_ ( .A1(_01954_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01994_ ) );
OR3_X1 _09550_ ( .A1(_01994_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01995_ ) );
OAI21_X1 _09551_ ( .A(\myclint.mtime [19] ), .B1(_01994_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01996_ ) );
AOI21_X1 _09552_ ( .A(fanout_net_1 ), .B1(_01995_ ), .B2(_01996_ ), .ZN(_00039_ ) );
AND2_X1 _09553_ ( .A1(_01783_ ), .A2(\myclint.mtime [17] ), .ZN(_01997_ ) );
OAI21_X1 _09554_ ( .A(_01934_ ), .B1(_01997_ ), .B2(\myclint.mtime [18] ), .ZN(_01998_ ) );
NOR2_X1 _09555_ ( .A1(_01998_ ), .A2(_01784_ ), .ZN(_00040_ ) );
INV_X1 _09556_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01999_ ) );
AND3_X1 _09557_ ( .A1(_01782_ ), .A2(_01999_ ), .A3(\myclint.mtime [15] ), .ZN(_02000_ ) );
AND2_X1 _09558_ ( .A1(_02000_ ), .A2(\myclint.mtime [17] ), .ZN(_02001_ ) );
OAI21_X1 _09559_ ( .A(_01774_ ), .B1(_02000_ ), .B2(\myclint.mtime [17] ), .ZN(_02002_ ) );
NOR2_X1 _09560_ ( .A1(_02001_ ), .A2(_02002_ ), .ZN(_00041_ ) );
AND2_X1 _09561_ ( .A1(_01782_ ), .A2(\myclint.mtime [15] ), .ZN(_02003_ ) );
OAI21_X1 _09562_ ( .A(_01934_ ), .B1(_02003_ ), .B2(\myclint.mtime [16] ), .ZN(_02004_ ) );
NOR2_X1 _09563_ ( .A1(_02004_ ), .A2(_01783_ ), .ZN(_00042_ ) );
AND3_X1 _09564_ ( .A1(_01779_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [11] ), .ZN(_02005_ ) );
AND2_X1 _09565_ ( .A1(_01778_ ), .A2(_02005_ ), .ZN(_02006_ ) );
NAND3_X1 _09566_ ( .A1(_02006_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_02007_ ) );
OR3_X1 _09567_ ( .A1(_02007_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_02008_ ) );
OAI21_X1 _09568_ ( .A(\myclint.mtime [15] ), .B1(_02007_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02009_ ) );
AOI21_X1 _09569_ ( .A(fanout_net_1 ), .B1(_02008_ ), .B2(_02009_ ), .ZN(_00043_ ) );
AND2_X1 _09570_ ( .A1(_01781_ ), .A2(\myclint.mtime [13] ), .ZN(_02010_ ) );
OAI21_X1 _09571_ ( .A(_01934_ ), .B1(_02010_ ), .B2(\myclint.mtime [14] ), .ZN(_02011_ ) );
NOR2_X1 _09572_ ( .A1(_02011_ ), .A2(_01782_ ), .ZN(_00044_ ) );
NAND3_X1 _09573_ ( .A1(_01864_ ), .A2(_01818_ ), .A3(_01865_ ), .ZN(_02012_ ) );
OR2_X1 _09574_ ( .A1(_02012_ ), .A2(\myclint.mtime [58] ), .ZN(_02013_ ) );
NAND2_X1 _09575_ ( .A1(_02012_ ), .A2(\myclint.mtime [58] ), .ZN(_02014_ ) );
AOI21_X1 _09576_ ( .A(fanout_net_1 ), .B1(_02013_ ), .B2(_02014_ ), .ZN(_00045_ ) );
INV_X1 _09577_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02015_ ) );
AND3_X1 _09578_ ( .A1(_01780_ ), .A2(_02015_ ), .A3(\myclint.mtime [11] ), .ZN(_02016_ ) );
AND2_X1 _09579_ ( .A1(_02016_ ), .A2(\myclint.mtime [13] ), .ZN(_02017_ ) );
OAI21_X1 _09580_ ( .A(_01774_ ), .B1(_02016_ ), .B2(\myclint.mtime [13] ), .ZN(_02018_ ) );
NOR2_X1 _09581_ ( .A1(_02017_ ), .A2(_02018_ ), .ZN(_00046_ ) );
AND2_X1 _09582_ ( .A1(_01780_ ), .A2(\myclint.mtime [11] ), .ZN(_02019_ ) );
OAI21_X1 _09583_ ( .A(_01887_ ), .B1(_02019_ ), .B2(\myclint.mtime [12] ), .ZN(_02020_ ) );
NOR2_X1 _09584_ ( .A1(_02020_ ), .A2(_01781_ ), .ZN(_00047_ ) );
AND2_X1 _09585_ ( .A1(_01778_ ), .A2(_01779_ ), .ZN(_02021_ ) );
INV_X1 _09586_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02022_ ) );
AND2_X1 _09587_ ( .A1(_02021_ ), .A2(_02022_ ), .ZN(_02023_ ) );
OAI21_X1 _09588_ ( .A(_01887_ ), .B1(_02023_ ), .B2(\myclint.mtime [11] ), .ZN(_02024_ ) );
AND3_X1 _09589_ ( .A1(_02021_ ), .A2(_02022_ ), .A3(\myclint.mtime [11] ), .ZN(_02025_ ) );
NOR2_X1 _09590_ ( .A1(_02024_ ), .A2(_02025_ ), .ZN(_00048_ ) );
OAI21_X1 _09591_ ( .A(_01887_ ), .B1(_02021_ ), .B2(\myclint.mtime [10] ), .ZN(_02026_ ) );
NOR2_X1 _09592_ ( .A1(_02026_ ), .A2(_01780_ ), .ZN(_00049_ ) );
INV_X1 _09593_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02027_ ) );
AND3_X1 _09594_ ( .A1(_01778_ ), .A2(\myclint.mtime [9] ), .A3(_02027_ ), .ZN(_02028_ ) );
AOI21_X1 _09595_ ( .A(\myclint.mtime [9] ), .B1(_01778_ ), .B2(_02027_ ), .ZN(_02029_ ) );
NOR3_X1 _09596_ ( .A1(_02028_ ), .A2(_02029_ ), .A3(fanout_net_1 ), .ZN(_00050_ ) );
OAI21_X1 _09597_ ( .A(_01774_ ), .B1(_01778_ ), .B2(\myclint.mtime [8] ), .ZN(_02030_ ) );
AOI21_X1 _09598_ ( .A(_02030_ ), .B1(\myclint.mtime [8] ), .B2(_01778_ ), .ZN(_00051_ ) );
AND2_X1 _09599_ ( .A1(_01776_ ), .A2(\myclint.mtime [5] ), .ZN(_02031_ ) );
INV_X1 _09600_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02032_ ) );
AND3_X1 _09601_ ( .A1(_02031_ ), .A2(_02032_ ), .A3(\myclint.mtime [7] ), .ZN(_02033_ ) );
AOI21_X1 _09602_ ( .A(\myclint.mtime [7] ), .B1(_02031_ ), .B2(_02032_ ), .ZN(_02034_ ) );
NOR3_X1 _09603_ ( .A1(_02033_ ), .A2(_02034_ ), .A3(fanout_net_1 ), .ZN(_00052_ ) );
OAI21_X1 _09604_ ( .A(_01887_ ), .B1(_02031_ ), .B2(\myclint.mtime [6] ), .ZN(_02035_ ) );
NOR2_X1 _09605_ ( .A1(_02035_ ), .A2(_01777_ ), .ZN(_00053_ ) );
AND2_X1 _09606_ ( .A1(_01775_ ), .A2(\myclint.mtime [3] ), .ZN(_02036_ ) );
INV_X1 _09607_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02037_ ) );
AND3_X1 _09608_ ( .A1(_02036_ ), .A2(\myclint.mtime [5] ), .A3(_02037_ ), .ZN(_02038_ ) );
AOI21_X1 _09609_ ( .A(\myclint.mtime [5] ), .B1(_02036_ ), .B2(_02037_ ), .ZN(_02039_ ) );
NOR3_X1 _09610_ ( .A1(_02038_ ), .A2(_02039_ ), .A3(fanout_net_1 ), .ZN(_00054_ ) );
OAI21_X1 _09611_ ( .A(_01887_ ), .B1(_02036_ ), .B2(\myclint.mtime [4] ), .ZN(_02040_ ) );
NOR2_X1 _09612_ ( .A1(_02040_ ), .A2(_01776_ ), .ZN(_00055_ ) );
BUF_X4 _09613_ ( .A(_01773_ ), .Z(_02041_ ) );
INV_X1 _09614_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02042_ ) );
AND3_X1 _09615_ ( .A1(_01815_ ), .A2(_02042_ ), .A3(_01816_ ), .ZN(_02043_ ) );
OAI21_X1 _09616_ ( .A(_02041_ ), .B1(_02043_ ), .B2(\myclint.mtime [57] ), .ZN(_02044_ ) );
AND3_X1 _09617_ ( .A1(_01840_ ), .A2(_02042_ ), .A3(_01816_ ), .ZN(_02045_ ) );
AOI21_X1 _09618_ ( .A(_02044_ ), .B1(_02045_ ), .B2(\myclint.mtime [57] ), .ZN(_00056_ ) );
AND2_X1 _09619_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_02046_ ) );
INV_X1 _09620_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02047_ ) );
AND3_X1 _09621_ ( .A1(_02046_ ), .A2(_02047_ ), .A3(\myclint.mtime [3] ), .ZN(_02048_ ) );
AOI21_X1 _09622_ ( .A(\myclint.mtime [3] ), .B1(_02046_ ), .B2(_02047_ ), .ZN(_02049_ ) );
NOR3_X1 _09623_ ( .A1(_02048_ ), .A2(_02049_ ), .A3(fanout_net_1 ), .ZN(_00057_ ) );
AOI21_X1 _09624_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_02050_ ) );
NOR3_X1 _09625_ ( .A1(_01775_ ), .A2(_02050_ ), .A3(fanout_net_1 ), .ZN(_00058_ ) );
NOR2_X1 _09626_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_02051_ ) );
NOR3_X1 _09627_ ( .A1(_02046_ ), .A2(_02051_ ), .A3(fanout_net_1 ), .ZN(_00059_ ) );
INV_X1 _09628_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_02052_ ) );
NOR2_X1 _09629_ ( .A1(_02052_ ), .A2(fanout_net_1 ), .ZN(_00060_ ) );
XNOR2_X1 _09630_ ( .A(_01866_ ), .B(\myclint.mtime [56] ), .ZN(_02053_ ) );
NOR2_X1 _09631_ ( .A1(_02053_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
NOR3_X1 _09632_ ( .A1(_01812_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01814_ ), .ZN(_02054_ ) );
OAI21_X1 _09633_ ( .A(_02041_ ), .B1(_02054_ ), .B2(\myclint.mtime [55] ), .ZN(_02055_ ) );
INV_X1 _09634_ ( .A(_01839_ ), .ZN(_02056_ ) );
NOR3_X1 _09635_ ( .A1(_02056_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01814_ ), .ZN(_02057_ ) );
AOI21_X1 _09636_ ( .A(_02055_ ), .B1(_02057_ ), .B2(\myclint.mtime [55] ), .ZN(_00062_ ) );
OR4_X1 _09637_ ( .A1(\myclint.mtime [54] ), .A2(_01863_ ), .A3(_01814_ ), .A4(_01872_ ), .ZN(_02058_ ) );
NAND3_X1 _09638_ ( .A1(_01864_ ), .A2(_01813_ ), .A3(_01871_ ), .ZN(_02059_ ) );
NAND2_X1 _09639_ ( .A1(_02059_ ), .A2(\myclint.mtime [54] ), .ZN(_02060_ ) );
AOI21_X1 _09640_ ( .A(fanout_net_2 ), .B1(_02058_ ), .B2(_02060_ ), .ZN(_00063_ ) );
MUX2_X1 _09641_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(fanout_net_44 ), .Z(_02061_ ) );
MUX2_X1 _09642_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(fanout_net_44 ), .Z(_02062_ ) );
MUX2_X1 _09643_ ( .A(_02061_ ), .B(_02062_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02063_ ) );
INV_X1 _09644_ ( .A(\IF_ID_pc [29] ), .ZN(_02064_ ) );
AND2_X1 _09645_ ( .A1(_02063_ ), .A2(_02064_ ), .ZN(_02065_ ) );
MUX2_X1 _09646_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(fanout_net_44 ), .Z(_02066_ ) );
MUX2_X1 _09647_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(fanout_net_44 ), .Z(_02067_ ) );
MUX2_X2 _09648_ ( .A(_02066_ ), .B(_02067_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02068_ ) );
INV_X1 _09649_ ( .A(\IF_ID_pc [20] ), .ZN(_02069_ ) );
MUX2_X1 _09650_ ( .A(\myifu.myicache.tag[0][2] ), .B(\myifu.myicache.tag[1][2] ), .S(fanout_net_44 ), .Z(_02070_ ) );
INV_X32 _09651_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_02071_ ) );
NAND2_X1 _09652_ ( .A1(_02070_ ), .A2(_02071_ ), .ZN(_02072_ ) );
MUX2_X1 _09653_ ( .A(\myifu.myicache.tag[2][2] ), .B(\myifu.myicache.tag[3][2] ), .S(fanout_net_44 ), .Z(_02073_ ) );
NAND2_X1 _09654_ ( .A1(_02073_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_02074_ ) );
NAND2_X1 _09655_ ( .A1(_02072_ ), .A2(_02074_ ), .ZN(_02075_ ) );
INV_X1 _09656_ ( .A(\IF_ID_pc [7] ), .ZN(_02076_ ) );
AOI22_X1 _09657_ ( .A1(_02068_ ), .A2(_02069_ ), .B1(_02075_ ), .B2(_02076_ ), .ZN(_02077_ ) );
MUX2_X1 _09658_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(fanout_net_44 ), .Z(_02078_ ) );
MUX2_X1 _09659_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(fanout_net_44 ), .Z(_02079_ ) );
MUX2_X1 _09660_ ( .A(_02078_ ), .B(_02079_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02080_ ) );
INV_X1 _09661_ ( .A(\IF_ID_pc [14] ), .ZN(_02081_ ) );
NAND2_X1 _09662_ ( .A1(_02080_ ), .A2(_02081_ ), .ZN(_02082_ ) );
INV_X1 _09663_ ( .A(\IF_ID_pc [18] ), .ZN(_02083_ ) );
MUX2_X1 _09664_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(fanout_net_44 ), .Z(_02084_ ) );
MUX2_X1 _09665_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(fanout_net_44 ), .Z(_02085_ ) );
MUX2_X1 _09666_ ( .A(_02084_ ), .B(_02085_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02086_ ) );
OAI211_X1 _09667_ ( .A(_02077_ ), .B(_02082_ ), .C1(_02083_ ), .C2(_02086_ ), .ZN(_02087_ ) );
MUX2_X1 _09668_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(fanout_net_44 ), .Z(_02088_ ) );
MUX2_X1 _09669_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(fanout_net_44 ), .Z(_02089_ ) );
MUX2_X1 _09670_ ( .A(_02088_ ), .B(_02089_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02090_ ) );
INV_X1 _09671_ ( .A(\IF_ID_pc [21] ), .ZN(_02091_ ) );
AND2_X1 _09672_ ( .A1(_02090_ ), .A2(_02091_ ), .ZN(_02092_ ) );
OAI22_X1 _09673_ ( .A1(_02064_ ), .A2(_02063_ ), .B1(_02090_ ), .B2(_02091_ ), .ZN(_02093_ ) );
OR4_X2 _09674_ ( .A1(_02065_ ), .A2(_02087_ ), .A3(_02092_ ), .A4(_02093_ ), .ZN(_02094_ ) );
MUX2_X1 _09675_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(fanout_net_44 ), .Z(_02095_ ) );
MUX2_X1 _09676_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(fanout_net_44 ), .Z(_02096_ ) );
MUX2_X1 _09677_ ( .A(_02095_ ), .B(_02096_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02097_ ) );
INV_X1 _09678_ ( .A(\IF_ID_pc [12] ), .ZN(_02098_ ) );
NAND2_X1 _09679_ ( .A1(_02097_ ), .A2(_02098_ ), .ZN(_02099_ ) );
INV_X1 _09680_ ( .A(\IF_ID_pc [25] ), .ZN(_02100_ ) );
MUX2_X1 _09681_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(fanout_net_44 ), .Z(_02101_ ) );
MUX2_X1 _09682_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_44 ), .Z(_02102_ ) );
MUX2_X1 _09683_ ( .A(_02101_ ), .B(_02102_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02103_ ) );
OAI221_X1 _09684_ ( .A(_02099_ ), .B1(_02069_ ), .B2(_02068_ ), .C1(_02100_ ), .C2(_02103_ ), .ZN(_02104_ ) );
MUX2_X1 _09685_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_44 ), .Z(_02105_ ) );
MUX2_X1 _09686_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_44 ), .Z(_02106_ ) );
MUX2_X1 _09687_ ( .A(_02105_ ), .B(_02106_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02107_ ) );
INV_X1 _09688_ ( .A(\IF_ID_pc [16] ), .ZN(_02108_ ) );
NAND2_X1 _09689_ ( .A1(_02107_ ), .A2(_02108_ ), .ZN(_02109_ ) );
OAI21_X1 _09690_ ( .A(_02109_ ), .B1(_02098_ ), .B2(_02097_ ), .ZN(_02110_ ) );
OAI22_X1 _09691_ ( .A1(_02081_ ), .A2(_02080_ ), .B1(_02107_ ), .B2(_02108_ ), .ZN(_02111_ ) );
NOR4_X4 _09692_ ( .A1(_02094_ ), .A2(_02104_ ), .A3(_02110_ ), .A4(_02111_ ), .ZN(_02112_ ) );
OR2_X1 _09693_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_02113_ ) );
BUF_X4 _09694_ ( .A(_02071_ ), .Z(_02114_ ) );
INV_X32 _09695_ ( .A(fanout_net_44 ), .ZN(_02115_ ) );
BUF_X4 _09696_ ( .A(_02115_ ), .Z(_02116_ ) );
OAI211_X1 _09697_ ( .A(_02113_ ), .B(_02114_ ), .C1(_02116_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_02117_ ) );
OR2_X1 _09698_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][1] ), .ZN(_02118_ ) );
OAI211_X1 _09699_ ( .A(_02118_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02116_ ), .C2(\myifu.myicache.tag[3][1] ), .ZN(_02119_ ) );
AND3_X1 _09700_ ( .A1(_02117_ ), .A2(_02119_ ), .A3(\IF_ID_pc [6] ), .ZN(_02120_ ) );
OR2_X1 _09701_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][26] ), .ZN(_02121_ ) );
BUF_X4 _09702_ ( .A(_02115_ ), .Z(_02122_ ) );
OAI211_X1 _09703_ ( .A(_02121_ ), .B(_02114_ ), .C1(_02122_ ), .C2(\myifu.myicache.tag[1][26] ), .ZN(_02123_ ) );
OR2_X1 _09704_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][26] ), .ZN(_02124_ ) );
BUF_X32 _09705_ ( .A(_02115_ ), .Z(_02125_ ) );
OAI211_X1 _09706_ ( .A(_02124_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02125_ ), .C2(\myifu.myicache.tag[3][26] ), .ZN(_02126_ ) );
INV_X1 _09707_ ( .A(\IF_ID_pc [31] ), .ZN(_02127_ ) );
AND3_X1 _09708_ ( .A1(_02123_ ), .A2(_02126_ ), .A3(_02127_ ), .ZN(_02128_ ) );
AOI21_X1 _09709_ ( .A(_02127_ ), .B1(_02123_ ), .B2(_02126_ ), .ZN(_02129_ ) );
OR2_X1 _09710_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][0] ), .ZN(_02130_ ) );
OAI211_X1 _09711_ ( .A(_02130_ ), .B(_02071_ ), .C1(_02125_ ), .C2(\myifu.myicache.tag[1][0] ), .ZN(_02131_ ) );
OR2_X1 _09712_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][0] ), .ZN(_02132_ ) );
OAI211_X1 _09713_ ( .A(_02132_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02125_ ), .C2(\myifu.myicache.tag[3][0] ), .ZN(_02133_ ) );
AND3_X1 _09714_ ( .A1(_02131_ ), .A2(_02133_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02134_ ) );
AOI21_X1 _09715_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02131_ ), .B2(_02133_ ), .ZN(_02135_ ) );
OAI22_X1 _09716_ ( .A1(_02128_ ), .A2(_02129_ ), .B1(_02134_ ), .B2(_02135_ ), .ZN(_02136_ ) );
OR2_X1 _09717_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][12] ), .ZN(_02137_ ) );
OAI211_X1 _09718_ ( .A(_02137_ ), .B(_02071_ ), .C1(_02122_ ), .C2(\myifu.myicache.tag[1][12] ), .ZN(_02138_ ) );
OR2_X1 _09719_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][12] ), .ZN(_02139_ ) );
OAI211_X1 _09720_ ( .A(_02139_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02122_ ), .C2(\myifu.myicache.tag[3][12] ), .ZN(_02140_ ) );
NAND2_X1 _09721_ ( .A1(_02138_ ), .A2(_02140_ ), .ZN(_02141_ ) );
INV_X1 _09722_ ( .A(\IF_ID_pc [17] ), .ZN(_02142_ ) );
XNOR2_X1 _09723_ ( .A(_02141_ ), .B(_02142_ ), .ZN(_02143_ ) );
AOI21_X1 _09724_ ( .A(\IF_ID_pc [6] ), .B1(_02117_ ), .B2(_02119_ ), .ZN(_02144_ ) );
OR4_X1 _09725_ ( .A1(_02120_ ), .A2(_02136_ ), .A3(_02143_ ), .A4(_02144_ ), .ZN(_02145_ ) );
OR2_X1 _09726_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][10] ), .ZN(_02146_ ) );
OAI211_X1 _09727_ ( .A(_02146_ ), .B(_02114_ ), .C1(_02122_ ), .C2(\myifu.myicache.tag[1][10] ), .ZN(_02147_ ) );
OR2_X1 _09728_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][10] ), .ZN(_02148_ ) );
OAI211_X1 _09729_ ( .A(_02148_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02125_ ), .C2(\myifu.myicache.tag[3][10] ), .ZN(_02149_ ) );
INV_X1 _09730_ ( .A(\IF_ID_pc [15] ), .ZN(_02150_ ) );
AND3_X1 _09731_ ( .A1(_02147_ ), .A2(_02149_ ), .A3(_02150_ ), .ZN(_02151_ ) );
AOI21_X1 _09732_ ( .A(_02150_ ), .B1(_02147_ ), .B2(_02149_ ), .ZN(_02152_ ) );
OR2_X1 _09733_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][8] ), .ZN(_02153_ ) );
OAI211_X1 _09734_ ( .A(_02153_ ), .B(_02071_ ), .C1(_02125_ ), .C2(\myifu.myicache.tag[1][8] ), .ZN(_02154_ ) );
OR2_X1 _09735_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][8] ), .ZN(_02155_ ) );
OAI211_X1 _09736_ ( .A(_02155_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02125_ ), .C2(\myifu.myicache.tag[3][8] ), .ZN(_02156_ ) );
INV_X1 _09737_ ( .A(\IF_ID_pc [13] ), .ZN(_02157_ ) );
AND3_X1 _09738_ ( .A1(_02154_ ), .A2(_02156_ ), .A3(_02157_ ), .ZN(_02158_ ) );
AOI21_X1 _09739_ ( .A(_02157_ ), .B1(_02154_ ), .B2(_02156_ ), .ZN(_02159_ ) );
OAI22_X1 _09740_ ( .A1(_02151_ ), .A2(_02152_ ), .B1(_02158_ ), .B2(_02159_ ), .ZN(_02160_ ) );
OR2_X1 _09741_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][17] ), .ZN(_02161_ ) );
OAI211_X1 _09742_ ( .A(_02161_ ), .B(_02071_ ), .C1(_02125_ ), .C2(\myifu.myicache.tag[1][17] ), .ZN(_02162_ ) );
OR2_X1 _09743_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][17] ), .ZN(_02163_ ) );
OAI211_X1 _09744_ ( .A(_02163_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02125_ ), .C2(\myifu.myicache.tag[3][17] ), .ZN(_02164_ ) );
NAND2_X1 _09745_ ( .A1(_02162_ ), .A2(_02164_ ), .ZN(_02165_ ) );
INV_X1 _09746_ ( .A(\IF_ID_pc [22] ), .ZN(_02166_ ) );
XNOR2_X1 _09747_ ( .A(_02165_ ), .B(_02166_ ), .ZN(_02167_ ) );
OR2_X1 _09748_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][4] ), .ZN(_02168_ ) );
OAI211_X1 _09749_ ( .A(_02168_ ), .B(_02114_ ), .C1(_02122_ ), .C2(\myifu.myicache.tag[1][4] ), .ZN(_02169_ ) );
OR2_X1 _09750_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][4] ), .ZN(_02170_ ) );
OAI211_X1 _09751_ ( .A(_02170_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02122_ ), .C2(\myifu.myicache.tag[3][4] ), .ZN(_02171_ ) );
AND3_X1 _09752_ ( .A1(_02169_ ), .A2(_02171_ ), .A3(\IF_ID_pc [9] ), .ZN(_02172_ ) );
AOI21_X1 _09753_ ( .A(\IF_ID_pc [9] ), .B1(_02169_ ), .B2(_02171_ ), .ZN(_02173_ ) );
OR4_X1 _09754_ ( .A1(_02160_ ), .A2(_02167_ ), .A3(_02172_ ), .A4(_02173_ ), .ZN(_02174_ ) );
OR2_X1 _09755_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][6] ), .ZN(_02175_ ) );
OAI211_X1 _09756_ ( .A(_02175_ ), .B(_02114_ ), .C1(_02116_ ), .C2(\myifu.myicache.tag[1][6] ), .ZN(_02176_ ) );
OR2_X1 _09757_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][6] ), .ZN(_02177_ ) );
OAI211_X1 _09758_ ( .A(_02177_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02116_ ), .C2(\myifu.myicache.tag[3][6] ), .ZN(_02178_ ) );
AND3_X1 _09759_ ( .A1(_02176_ ), .A2(_02178_ ), .A3(\IF_ID_pc [11] ), .ZN(_02179_ ) );
OR2_X4 _09760_ ( .A1(_02125_ ), .A2(\myifu.myicache.tag[3][14] ), .ZN(_02180_ ) );
OAI211_X1 _09761_ ( .A(_02180_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][14] ), .ZN(_02181_ ) );
OR2_X1 _09762_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][14] ), .ZN(_02182_ ) );
OAI211_X1 _09763_ ( .A(_02182_ ), .B(_02114_ ), .C1(_02116_ ), .C2(\myifu.myicache.tag[1][14] ), .ZN(_02183_ ) );
AOI21_X1 _09764_ ( .A(\IF_ID_pc [19] ), .B1(_02181_ ), .B2(_02183_ ), .ZN(_02184_ ) );
OR2_X1 _09765_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][23] ), .ZN(_02185_ ) );
OAI211_X1 _09766_ ( .A(_02185_ ), .B(_02114_ ), .C1(_02122_ ), .C2(\myifu.myicache.tag[1][23] ), .ZN(_02186_ ) );
OR2_X1 _09767_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][23] ), .ZN(_02187_ ) );
OAI211_X1 _09768_ ( .A(_02187_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02122_ ), .C2(\myifu.myicache.tag[3][23] ), .ZN(_02188_ ) );
AND3_X1 _09769_ ( .A1(_02186_ ), .A2(_02188_ ), .A3(\IF_ID_pc [28] ), .ZN(_02189_ ) );
AOI21_X1 _09770_ ( .A(\IF_ID_pc [11] ), .B1(_02176_ ), .B2(_02178_ ), .ZN(_02190_ ) );
OR4_X1 _09771_ ( .A1(_02179_ ), .A2(_02184_ ), .A3(_02189_ ), .A4(_02190_ ), .ZN(_02191_ ) );
MUX2_X1 _09772_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02192_ ) );
MUX2_X1 _09773_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02193_ ) );
MUX2_X1 _09774_ ( .A(_02192_ ), .B(_02193_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02194_ ) );
NAND3_X1 _09775_ ( .A1(_02181_ ), .A2(\IF_ID_pc [19] ), .A3(_02183_ ), .ZN(_02195_ ) );
OR2_X1 _09776_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][21] ), .ZN(_02196_ ) );
OAI211_X1 _09777_ ( .A(_02196_ ), .B(_02114_ ), .C1(_02116_ ), .C2(\myifu.myicache.tag[1][21] ), .ZN(_02197_ ) );
OR2_X1 _09778_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][21] ), .ZN(_02198_ ) );
OAI211_X1 _09779_ ( .A(_02198_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02116_ ), .C2(\myifu.myicache.tag[3][21] ), .ZN(_02199_ ) );
INV_X1 _09780_ ( .A(\IF_ID_pc [26] ), .ZN(_02200_ ) );
AND3_X1 _09781_ ( .A1(_02197_ ), .A2(_02199_ ), .A3(_02200_ ), .ZN(_02201_ ) );
AOI21_X1 _09782_ ( .A(_02200_ ), .B1(_02197_ ), .B2(_02199_ ), .ZN(_02202_ ) );
OAI211_X1 _09783_ ( .A(_02194_ ), .B(_02195_ ), .C1(_02201_ ), .C2(_02202_ ), .ZN(_02203_ ) );
NOR4_X2 _09784_ ( .A1(_02145_ ), .A2(_02174_ ), .A3(_02191_ ), .A4(_02203_ ), .ZN(_02204_ ) );
MUX2_X1 _09785_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02205_ ) );
MUX2_X1 _09786_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02206_ ) );
MUX2_X1 _09787_ ( .A(_02205_ ), .B(_02206_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02207_ ) );
INV_X1 _09788_ ( .A(\IF_ID_pc [10] ), .ZN(_02208_ ) );
XNOR2_X1 _09789_ ( .A(_02207_ ), .B(_02208_ ), .ZN(_02209_ ) );
AOI21_X1 _09790_ ( .A(\IF_ID_pc [28] ), .B1(_02186_ ), .B2(_02188_ ), .ZN(_02210_ ) );
OR2_X2 _09791_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][19] ), .ZN(_02211_ ) );
OAI211_X1 _09792_ ( .A(_02211_ ), .B(_02114_ ), .C1(_02116_ ), .C2(\myifu.myicache.tag[1][19] ), .ZN(_02212_ ) );
OR2_X2 _09793_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][19] ), .ZN(_02213_ ) );
OAI211_X2 _09794_ ( .A(_02213_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02122_ ), .C2(\myifu.myicache.tag[3][19] ), .ZN(_02214_ ) );
AND3_X1 _09795_ ( .A1(_02212_ ), .A2(_02214_ ), .A3(\IF_ID_pc [24] ), .ZN(_02215_ ) );
OR3_X1 _09796_ ( .A1(_02209_ ), .A2(_02210_ ), .A3(_02215_ ), .ZN(_02216_ ) );
MUX2_X1 _09797_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02217_ ) );
MUX2_X1 _09798_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02218_ ) );
MUX2_X1 _09799_ ( .A(_02217_ ), .B(_02218_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02219_ ) );
XNOR2_X1 _09800_ ( .A(_02219_ ), .B(\IF_ID_pc [27] ), .ZN(_02220_ ) );
NAND2_X1 _09801_ ( .A1(_02086_ ), .A2(_02083_ ), .ZN(_02221_ ) );
INV_X1 _09802_ ( .A(\IF_ID_pc [23] ), .ZN(_02222_ ) );
AND2_X1 _09803_ ( .A1(_02125_ ), .A2(\myifu.myicache.tag[0][18] ), .ZN(_02223_ ) );
AOI211_X1 _09804_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B(_02223_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[1][18] ), .ZN(_02224_ ) );
AND2_X1 _09805_ ( .A1(_02122_ ), .A2(\myifu.myicache.tag[2][18] ), .ZN(_02225_ ) );
AOI21_X1 _09806_ ( .A(_02225_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myifu.myicache.tag[3][18] ), .ZN(_02226_ ) );
AOI21_X1 _09807_ ( .A(_02224_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_02226_ ), .ZN(_02227_ ) );
OAI211_X1 _09808_ ( .A(_02220_ ), .B(_02221_ ), .C1(_02222_ ), .C2(_02227_ ), .ZN(_02228_ ) );
NAND2_X1 _09809_ ( .A1(_02227_ ), .A2(_02222_ ), .ZN(_02229_ ) );
MUX2_X1 _09810_ ( .A(\myifu.myicache.tag[0][3] ), .B(\myifu.myicache.tag[1][3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02230_ ) );
MUX2_X1 _09811_ ( .A(\myifu.myicache.tag[2][3] ), .B(\myifu.myicache.tag[3][3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02231_ ) );
MUX2_X1 _09812_ ( .A(_02230_ ), .B(_02231_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02232_ ) );
INV_X1 _09813_ ( .A(\IF_ID_pc [8] ), .ZN(_02233_ ) );
AOI22_X1 _09814_ ( .A1(_02100_ ), .A2(_02103_ ), .B1(_02232_ ), .B2(_02233_ ), .ZN(_02234_ ) );
OAI211_X1 _09815_ ( .A(_02229_ ), .B(_02234_ ), .C1(_02233_ ), .C2(_02232_ ), .ZN(_02235_ ) );
OR2_X2 _09816_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][25] ), .ZN(_02236_ ) );
OAI211_X1 _09817_ ( .A(_02236_ ), .B(_02114_ ), .C1(_02116_ ), .C2(\myifu.myicache.tag[1][25] ), .ZN(_02237_ ) );
OR2_X4 _09818_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][25] ), .ZN(_02238_ ) );
OAI211_X1 _09819_ ( .A(_02238_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02116_ ), .C2(\myifu.myicache.tag[3][25] ), .ZN(_02239_ ) );
AND3_X1 _09820_ ( .A1(_02237_ ), .A2(_02239_ ), .A3(\IF_ID_pc [30] ), .ZN(_02240_ ) );
AND3_X1 _09821_ ( .A1(_02072_ ), .A2(_02074_ ), .A3(\IF_ID_pc [7] ), .ZN(_02241_ ) );
AOI21_X1 _09822_ ( .A(\IF_ID_pc [30] ), .B1(_02237_ ), .B2(_02239_ ), .ZN(_02242_ ) );
AOI21_X1 _09823_ ( .A(\IF_ID_pc [24] ), .B1(_02212_ ), .B2(_02214_ ), .ZN(_02243_ ) );
OR4_X1 _09824_ ( .A1(_02240_ ), .A2(_02241_ ), .A3(_02242_ ), .A4(_02243_ ), .ZN(_02244_ ) );
NOR4_X2 _09825_ ( .A1(_02216_ ), .A2(_02228_ ), .A3(_02235_ ), .A4(_02244_ ), .ZN(_02245_ ) );
NAND3_X2 _09826_ ( .A1(_02112_ ), .A2(_02204_ ), .A3(_02245_ ), .ZN(_02246_ ) );
AND2_X4 _09827_ ( .A1(_02246_ ), .A2(\myifu.state [0] ), .ZN(_02247_ ) );
INV_X1 _09828_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_02248_ ) );
NOR2_X4 _09829_ ( .A1(_02247_ ), .A2(_02248_ ), .ZN(_02249_ ) );
NOR2_X1 _09830_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_02250_ ) );
NOR2_X4 _09831_ ( .A1(_02249_ ), .A2(_02250_ ), .ZN(_02251_ ) );
INV_X1 _09832_ ( .A(\EX_LS_flag [2] ), .ZN(_02252_ ) );
NAND4_X1 _09833_ ( .A1(_02252_ ), .A2(\mylsu.state [0] ), .A3(\EX_LS_flag [1] ), .A4(\EX_LS_flag [0] ), .ZN(_02253_ ) );
INV_X1 _09834_ ( .A(EXU_valid_LSU ), .ZN(_02254_ ) );
NOR2_X1 _09835_ ( .A1(_02253_ ), .A2(_02254_ ), .ZN(_02255_ ) );
INV_X1 _09836_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_02256_ ) );
NOR2_X2 _09837_ ( .A1(_02255_ ), .A2(_02256_ ), .ZN(_02257_ ) );
NOR2_X4 _09838_ ( .A1(_02251_ ), .A2(_02257_ ), .ZN(_02258_ ) );
BUF_X8 _09839_ ( .A(_02258_ ), .Z(_02259_ ) );
CLKBUF_X2 _09840_ ( .A(_02254_ ), .Z(_02260_ ) );
OR3_X1 _09841_ ( .A1(_02253_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(_02260_ ), .ZN(_02261_ ) );
BUF_X4 _09842_ ( .A(_02255_ ), .Z(_02262_ ) );
OAI211_X1 _09843_ ( .A(_02259_ ), .B(_02261_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_02262_ ), .ZN(_02263_ ) );
INV_X1 _09844_ ( .A(\IF_ID_pc [30] ), .ZN(_02264_ ) );
INV_X4 _09845_ ( .A(_02251_ ), .ZN(_02265_ ) );
BUF_X8 _09846_ ( .A(_02265_ ), .Z(_02266_ ) );
OAI21_X1 _09847_ ( .A(_02263_ ), .B1(_02264_ ), .B2(_02266_ ), .ZN(\io_master_araddr [30] ) );
OR3_X1 _09848_ ( .A1(_02253_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(_02260_ ), .ZN(_02267_ ) );
OAI211_X1 _09849_ ( .A(_02259_ ), .B(_02267_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_02255_ ), .ZN(_02268_ ) );
INV_X1 _09850_ ( .A(\IF_ID_pc [28] ), .ZN(_02269_ ) );
OAI21_X1 _09851_ ( .A(_02268_ ), .B1(_02269_ ), .B2(_02265_ ), .ZN(\io_master_araddr [28] ) );
BUF_X16 _09852_ ( .A(_02259_ ), .Z(_02270_ ) );
CLKBUF_X2 _09853_ ( .A(_02253_ ), .Z(_02271_ ) );
CLKBUF_X2 _09854_ ( .A(_02254_ ), .Z(_02272_ ) );
OR3_X1 _09855_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(_02272_ ), .ZN(_02273_ ) );
BUF_X4 _09856_ ( .A(_02262_ ), .Z(_02274_ ) );
OAI211_X1 _09857_ ( .A(_02270_ ), .B(_02273_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_02274_ ), .ZN(_02275_ ) );
INV_X1 _09858_ ( .A(\IF_ID_pc [24] ), .ZN(_02276_ ) );
OAI21_X1 _09859_ ( .A(_02275_ ), .B1(_02276_ ), .B2(_02266_ ), .ZN(\io_master_araddr [24] ) );
INV_X1 _09860_ ( .A(_02257_ ), .ZN(_02277_ ) );
OR3_X1 _09861_ ( .A1(_02253_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(_02260_ ), .ZN(_02278_ ) );
OAI211_X1 _09862_ ( .A(_02277_ ), .B(_02278_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_02262_ ), .ZN(_02279_ ) );
INV_X1 _09863_ ( .A(\IF_ID_pc [27] ), .ZN(_02280_ ) );
MUX2_X1 _09864_ ( .A(_02279_ ), .B(_02280_ ), .S(_02251_ ), .Z(_02281_ ) );
INV_X1 _09865_ ( .A(_02281_ ), .ZN(\io_master_araddr [27] ) );
OR4_X1 _09866_ ( .A1(\io_master_araddr [30] ), .A2(\io_master_araddr [28] ), .A3(\io_master_araddr [24] ), .A4(\io_master_araddr [27] ), .ZN(_02282_ ) );
OR3_X1 _09867_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(_02272_ ), .ZN(_02283_ ) );
OAI211_X1 _09868_ ( .A(_02270_ ), .B(_02283_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_02274_ ), .ZN(_02284_ ) );
OAI221_X1 _09869_ ( .A(\IF_ID_pc [26] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02247_ ), .C2(_02248_ ), .ZN(_02285_ ) );
AND2_X1 _09870_ ( .A1(_02284_ ), .A2(_02285_ ), .ZN(_02286_ ) );
OR3_X1 _09871_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [25] ), .A3(_02272_ ), .ZN(_02287_ ) );
OAI211_X4 _09872_ ( .A(_02270_ ), .B(_02287_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_02262_ ), .ZN(_02288_ ) );
OAI21_X2 _09873_ ( .A(_02288_ ), .B1(_02100_ ), .B2(_02266_ ), .ZN(\io_master_araddr [25] ) );
NAND2_X1 _09874_ ( .A1(_02286_ ), .A2(\io_master_araddr [25] ), .ZN(_02289_ ) );
BUF_X2 _09875_ ( .A(_02271_ ), .Z(_02290_ ) );
OR3_X1 _09876_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(_02272_ ), .ZN(_02291_ ) );
OAI211_X1 _09877_ ( .A(_02270_ ), .B(_02291_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_02274_ ), .ZN(_02292_ ) );
BUF_X4 _09878_ ( .A(_02266_ ), .Z(_02293_ ) );
OAI21_X1 _09879_ ( .A(_02292_ ), .B1(_02142_ ), .B2(_02293_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09880_ ( .A1(_02253_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(_02260_ ), .ZN(_02294_ ) );
OAI211_X1 _09881_ ( .A(_02258_ ), .B(_02294_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_02255_ ), .ZN(_02295_ ) );
OAI21_X1 _09882_ ( .A(_02295_ ), .B1(_02166_ ), .B2(_02265_ ), .ZN(\io_master_araddr [22] ) );
NOR4_X1 _09883_ ( .A1(_02282_ ), .A2(_02289_ ), .A3(\io_master_araddr [17] ), .A4(\io_master_araddr [22] ), .ZN(_02296_ ) );
OR3_X1 _09884_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(_02260_ ), .ZN(_02297_ ) );
OAI211_X1 _09885_ ( .A(_02259_ ), .B(_02297_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_02262_ ), .ZN(_02298_ ) );
OAI21_X1 _09886_ ( .A(_02298_ ), .B1(_02127_ ), .B2(_02266_ ), .ZN(\io_master_araddr [31] ) );
OR3_X1 _09887_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(_02260_ ), .ZN(_02299_ ) );
OAI211_X1 _09888_ ( .A(_02259_ ), .B(_02299_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_02262_ ), .ZN(_02300_ ) );
OAI21_X1 _09889_ ( .A(_02300_ ), .B1(_02064_ ), .B2(_02266_ ), .ZN(\io_master_araddr [29] ) );
OR3_X1 _09890_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(_02272_ ), .ZN(_02301_ ) );
OAI211_X1 _09891_ ( .A(_02270_ ), .B(_02301_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_02274_ ), .ZN(_02302_ ) );
OAI21_X1 _09892_ ( .A(_02302_ ), .B1(_02108_ ), .B2(_02293_ ), .ZN(\io_master_araddr [16] ) );
OR3_X1 _09893_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(_02260_ ), .ZN(_02303_ ) );
OAI211_X1 _09894_ ( .A(_02259_ ), .B(_02303_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_02262_ ), .ZN(_02304_ ) );
OAI21_X1 _09895_ ( .A(_02304_ ), .B1(_02222_ ), .B2(_02266_ ), .ZN(\io_master_araddr [23] ) );
NOR4_X1 _09896_ ( .A1(\io_master_araddr [31] ), .A2(\io_master_araddr [29] ), .A3(\io_master_araddr [16] ), .A4(\io_master_araddr [23] ), .ZN(_02305_ ) );
OR3_X1 _09897_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(_02272_ ), .ZN(_02306_ ) );
OAI211_X1 _09898_ ( .A(_02259_ ), .B(_02306_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_02262_ ), .ZN(_02307_ ) );
INV_X1 _09899_ ( .A(\IF_ID_pc [19] ), .ZN(_02308_ ) );
OAI21_X1 _09900_ ( .A(_02307_ ), .B1(_02308_ ), .B2(_02266_ ), .ZN(\io_master_araddr [19] ) );
OR3_X1 _09901_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(_02260_ ), .ZN(_02309_ ) );
OAI211_X1 _09902_ ( .A(_02259_ ), .B(_02309_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_02262_ ), .ZN(_02310_ ) );
OAI21_X1 _09903_ ( .A(_02310_ ), .B1(_02069_ ), .B2(_02266_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09904_ ( .A1(_02271_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(_02260_ ), .ZN(_02311_ ) );
OAI211_X1 _09905_ ( .A(_02259_ ), .B(_02311_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_02262_ ), .ZN(_02312_ ) );
OAI21_X1 _09906_ ( .A(_02312_ ), .B1(_02083_ ), .B2(_02266_ ), .ZN(\io_master_araddr [18] ) );
OR3_X1 _09907_ ( .A1(_02253_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(_02260_ ), .ZN(_02313_ ) );
OAI211_X1 _09908_ ( .A(_02259_ ), .B(_02313_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_02255_ ), .ZN(_02314_ ) );
OAI21_X1 _09909_ ( .A(_02314_ ), .B1(_02091_ ), .B2(_02265_ ), .ZN(\io_master_araddr [21] ) );
NOR4_X1 _09910_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [18] ), .A4(\io_master_araddr [21] ), .ZN(_02315_ ) );
AND2_X1 _09911_ ( .A1(_02305_ ), .A2(_02315_ ), .ZN(_02316_ ) );
AND2_X2 _09912_ ( .A1(_02296_ ), .A2(_02316_ ), .ZN(_02317_ ) );
INV_X1 _09913_ ( .A(_02317_ ), .ZN(_02318_ ) );
CLKBUF_X2 _09914_ ( .A(_02251_ ), .Z(_02319_ ) );
CLKBUF_X2 _09915_ ( .A(_02319_ ), .Z(_02320_ ) );
BUF_X2 _09916_ ( .A(_02320_ ), .Z(_02321_ ) );
OR2_X1 _09917_ ( .A1(\EX_LS_dest_csreg_mem [27] ), .A2(\EX_LS_dest_csreg_mem [25] ), .ZN(_02322_ ) );
OR3_X1 _09918_ ( .A1(_02322_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(\EX_LS_dest_csreg_mem [24] ), .ZN(_02323_ ) );
OR4_X1 _09919_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(_02323_ ), .A3(\EX_LS_dest_csreg_mem [30] ), .A4(\EX_LS_dest_csreg_mem [29] ), .ZN(_02324_ ) );
NOR2_X1 _09920_ ( .A1(_02324_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .ZN(_02325_ ) );
AND2_X4 _09921_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02326_ ) );
AND2_X4 _09922_ ( .A1(_02326_ ), .A2(_02252_ ), .ZN(_02327_ ) );
AND2_X1 _09923_ ( .A1(_02325_ ), .A2(_02327_ ), .ZN(_02328_ ) );
NOR2_X1 _09924_ ( .A1(fanout_net_4 ), .A2(\EX_LS_dest_csreg_mem [1] ), .ZN(_02329_ ) );
INV_X1 _09925_ ( .A(_02329_ ), .ZN(_02330_ ) );
INV_X1 _09926_ ( .A(\EX_LS_typ [1] ), .ZN(_02331_ ) );
INV_X1 _09927_ ( .A(\EX_LS_typ [3] ), .ZN(_02332_ ) );
NAND4_X1 _09928_ ( .A1(_02330_ ), .A2(_02331_ ), .A3(_02332_ ), .A4(\EX_LS_typ [2] ), .ZN(_02333_ ) );
AND2_X1 _09929_ ( .A1(fanout_net_4 ), .A2(\EX_LS_typ [1] ), .ZN(_02334_ ) );
NOR2_X1 _09930_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02335_ ) );
NAND2_X1 _09931_ ( .A1(_02334_ ), .A2(_02335_ ), .ZN(_02336_ ) );
AOI21_X1 _09932_ ( .A(\EX_LS_typ [0] ), .B1(_02333_ ), .B2(_02336_ ), .ZN(_02337_ ) );
AND3_X1 _09933_ ( .A1(_02334_ ), .A2(\EX_LS_typ [0] ), .A3(_02335_ ), .ZN(_02338_ ) );
OR2_X1 _09934_ ( .A1(_02337_ ), .A2(_02338_ ), .ZN(_02339_ ) );
INV_X1 _09935_ ( .A(\EX_LS_typ [4] ), .ZN(_02340_ ) );
AND2_X1 _09936_ ( .A1(_02327_ ), .A2(_02340_ ), .ZN(_02341_ ) );
AND2_X1 _09937_ ( .A1(_02339_ ), .A2(_02341_ ), .ZN(_02342_ ) );
NOR2_X1 _09938_ ( .A1(_02328_ ), .A2(_02342_ ), .ZN(_02343_ ) );
INV_X32 _09939_ ( .A(\EX_LS_flag [1] ), .ZN(_02344_ ) );
NOR2_X2 _09940_ ( .A1(_02344_ ), .A2(\EX_LS_flag [0] ), .ZN(_02345_ ) );
AND2_X1 _09941_ ( .A1(_02345_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02346_ ) );
AND2_X1 _09942_ ( .A1(_02325_ ), .A2(_02346_ ), .ZN(_02347_ ) );
NAND2_X1 _09943_ ( .A1(\EX_LS_typ [2] ), .A2(\EX_LS_typ [0] ), .ZN(_02348_ ) );
NOR4_X1 _09944_ ( .A1(_02329_ ), .A2(_02348_ ), .A3(_02331_ ), .A4(_02332_ ), .ZN(_02349_ ) );
OR2_X1 _09945_ ( .A1(_02349_ ), .A2(_02338_ ), .ZN(_02350_ ) );
NOR3_X1 _09946_ ( .A1(_02344_ ), .A2(\EX_LS_typ [4] ), .A3(\EX_LS_flag [0] ), .ZN(_02351_ ) );
AND2_X1 _09947_ ( .A1(_02351_ ), .A2(_02252_ ), .ZN(_02352_ ) );
AND2_X1 _09948_ ( .A1(_02350_ ), .A2(_02352_ ), .ZN(_02353_ ) );
NOR2_X1 _09949_ ( .A1(_02347_ ), .A2(_02353_ ), .ZN(_02354_ ) );
AND2_X1 _09950_ ( .A1(_02343_ ), .A2(_02354_ ), .ZN(_02355_ ) );
AOI21_X1 _09951_ ( .A(_02321_ ), .B1(_02274_ ), .B2(_02355_ ), .ZN(_02356_ ) );
NOR2_X1 _09952_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02357_ ) );
AOI211_X1 _09953_ ( .A(_02250_ ), .B(_02249_ ), .C1(\myifu.state [0] ), .C2(_02357_ ), .ZN(_02358_ ) );
NOR3_X1 _09954_ ( .A1(_02318_ ), .A2(_02356_ ), .A3(_02358_ ), .ZN(_02359_ ) );
OAI21_X1 _09955_ ( .A(_01887_ ), .B1(_02359_ ), .B2(\myclint.rvalid ), .ZN(_02360_ ) );
OR4_X2 _09956_ ( .A1(\io_master_araddr [31] ), .A2(\io_master_araddr [29] ), .A3(\io_master_araddr [30] ), .A4(\io_master_araddr [28] ), .ZN(_02361_ ) );
INV_X1 _09957_ ( .A(_02286_ ), .ZN(\io_master_araddr [26] ) );
OAI211_X2 _09958_ ( .A(\io_master_araddr [25] ), .B(_02275_ ), .C1(_02276_ ), .C2(_02293_ ), .ZN(_02362_ ) );
OR4_X4 _09959_ ( .A1(\io_master_araddr [27] ), .A2(_02361_ ), .A3(\io_master_araddr [26] ), .A4(_02362_ ), .ZN(_02363_ ) );
OR4_X2 _09960_ ( .A1(\io_master_araddr [23] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [21] ), .A4(\io_master_araddr [22] ), .ZN(_02364_ ) );
OR2_X1 _09961_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [18] ), .ZN(_02365_ ) );
OR4_X4 _09962_ ( .A1(\io_master_araddr [16] ), .A2(_02364_ ), .A3(\io_master_araddr [17] ), .A4(_02365_ ), .ZN(_02366_ ) );
NOR2_X4 _09963_ ( .A1(_02363_ ), .A2(_02366_ ), .ZN(_02367_ ) );
BUF_X2 _09964_ ( .A(_02367_ ), .Z(_02368_ ) );
BUF_X2 _09965_ ( .A(_02368_ ), .Z(_02369_ ) );
AOI211_X1 _09966_ ( .A(_02256_ ), .B(_02321_ ), .C1(_02274_ ), .C2(_02355_ ), .ZN(_02370_ ) );
AND3_X1 _09967_ ( .A1(_02246_ ), .A2(\myifu.state [0] ), .A3(_02357_ ), .ZN(_02371_ ) );
NOR4_X1 _09968_ ( .A1(_02249_ ), .A2(_02248_ ), .A3(_02250_ ), .A4(_02371_ ), .ZN(_02372_ ) );
NOR2_X1 _09969_ ( .A1(_02370_ ), .A2(_02372_ ), .ZN(_02373_ ) );
AND3_X1 _09970_ ( .A1(_02369_ ), .A2(\myclint.rvalid ), .A3(_02373_ ), .ZN(_02374_ ) );
NOR2_X1 _09971_ ( .A1(_02360_ ), .A2(_02374_ ), .ZN(_00064_ ) );
INV_X1 _09972_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02375_ ) );
CLKBUF_X2 _09973_ ( .A(_02375_ ), .Z(_02376_ ) );
AND2_X1 _09974_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00065_ ) );
INV_X1 _09975_ ( .A(\LS_WB_wdata_csreg [4] ), .ZN(_02377_ ) );
NOR2_X1 _09976_ ( .A1(_02377_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00066_ ) );
AND2_X1 _09977_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00067_ ) );
AND2_X1 _09978_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00068_ ) );
AND2_X1 _09979_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00069_ ) );
AND2_X1 _09980_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [20] ), .ZN(_00070_ ) );
AND2_X1 _09981_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [19] ), .ZN(_00071_ ) );
AND2_X1 _09982_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [18] ), .ZN(_00072_ ) );
AND2_X1 _09983_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [17] ), .ZN(_00073_ ) );
AND2_X1 _09984_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00074_ ) );
AND2_X1 _09985_ ( .A1(_02376_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00075_ ) );
CLKBUF_X2 _09986_ ( .A(_02375_ ), .Z(_02378_ ) );
AND2_X1 _09987_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00076_ ) );
AND2_X1 _09988_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00077_ ) );
AND2_X1 _09989_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00078_ ) );
AND2_X1 _09990_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00079_ ) );
AND2_X1 _09991_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00080_ ) );
AND2_X1 _09992_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00081_ ) );
AND2_X1 _09993_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00082_ ) );
AND2_X1 _09994_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00083_ ) );
AND2_X1 _09995_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00084_ ) );
AND2_X1 _09996_ ( .A1(_02378_ ), .A2(\LS_WB_wdata_csreg [6] ), .ZN(_00085_ ) );
AND2_X1 _09997_ ( .A1(_02375_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00086_ ) );
AND2_X1 _09998_ ( .A1(_02375_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00087_ ) );
AND2_X1 _09999_ ( .A1(_02375_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00088_ ) );
AND2_X1 _10000_ ( .A1(_02375_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00089_ ) );
AND2_X1 _10001_ ( .A1(_02375_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00090_ ) );
AND2_X1 _10002_ ( .A1(_02375_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00091_ ) );
AND2_X1 _10003_ ( .A1(_02375_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00092_ ) );
INV_X1 _10004_ ( .A(_02347_ ), .ZN(_02379_ ) );
NAND3_X1 _10005_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02380_ ) );
OAI21_X1 _10006_ ( .A(_02336_ ), .B1(_02329_ ), .B2(_02380_ ), .ZN(_02381_ ) );
NAND3_X1 _10007_ ( .A1(_02252_ ), .A2(_02340_ ), .A3(\EX_LS_typ [0] ), .ZN(_02382_ ) );
NOR3_X1 _10008_ ( .A1(_02382_ ), .A2(_02344_ ), .A3(\EX_LS_flag [0] ), .ZN(_02383_ ) );
NAND2_X1 _10009_ ( .A1(_02381_ ), .A2(_02383_ ), .ZN(_02384_ ) );
AND2_X1 _10010_ ( .A1(_02379_ ), .A2(_02384_ ), .ZN(_02385_ ) );
INV_X1 _10011_ ( .A(_02385_ ), .ZN(_02386_ ) );
INV_X1 _10012_ ( .A(_02343_ ), .ZN(_02387_ ) );
NOR2_X1 _10013_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02388_ ) );
NAND2_X1 _10014_ ( .A1(_02388_ ), .A2(_01886_ ), .ZN(_02389_ ) );
NOR2_X1 _10015_ ( .A1(\myexu.pc_jump [27] ), .A2(\myexu.pc_jump [24] ), .ZN(_02390_ ) );
INV_X1 _10016_ ( .A(\myexu.pc_jump [26] ), .ZN(_02391_ ) );
INV_X1 _10017_ ( .A(\myexu.pc_jump [25] ), .ZN(_02392_ ) );
NAND3_X1 _10018_ ( .A1(_02390_ ), .A2(_02391_ ), .A3(_02392_ ), .ZN(_02393_ ) );
INV_X1 _10019_ ( .A(\myexu.pc_jump [31] ), .ZN(_02394_ ) );
INV_X1 _10020_ ( .A(\myexu.pc_jump [30] ), .ZN(_02395_ ) );
INV_X1 _10021_ ( .A(\myexu.pc_jump [29] ), .ZN(_02396_ ) );
INV_X1 _10022_ ( .A(\myexu.pc_jump [28] ), .ZN(_02397_ ) );
NAND4_X1 _10023_ ( .A1(_02394_ ), .A2(_02395_ ), .A3(_02396_ ), .A4(_02397_ ), .ZN(_02398_ ) );
NOR2_X1 _10024_ ( .A1(_02393_ ), .A2(_02398_ ), .ZN(_02399_ ) );
NOR2_X1 _10025_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02400_ ) );
INV_X1 _10026_ ( .A(_02400_ ), .ZN(_02401_ ) );
NOR3_X1 _10027_ ( .A1(_02399_ ), .A2(exception_quest_IDU ), .A3(_02401_ ), .ZN(_02402_ ) );
NOR4_X1 _10028_ ( .A1(_02386_ ), .A2(_02387_ ), .A3(_02389_ ), .A4(_02402_ ), .ZN(_00094_ ) );
AOI21_X1 _10029_ ( .A(_02389_ ), .B1(_02355_ ), .B2(exception_quest_IDU ), .ZN(_00095_ ) );
NOR2_X1 _10030_ ( .A1(fanout_net_2 ), .A2(fanout_net_16 ), .ZN(_02403_ ) );
INV_X1 _10031_ ( .A(_02403_ ), .ZN(_02404_ ) );
INV_X1 _10032_ ( .A(IDU_valid_EXU ), .ZN(_02405_ ) );
NOR2_X1 _10033_ ( .A1(_02405_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.pc_out_$_SDFFE_PP0P__Q_E ) );
INV_X1 _10034_ ( .A(\ID_EX_typ [7] ), .ZN(_02406_ ) );
NOR2_X1 _10035_ ( .A1(_02406_ ), .A2(\ID_EX_typ [5] ), .ZN(_02407_ ) );
BUF_X4 _10036_ ( .A(_02407_ ), .Z(_02408_ ) );
INV_X1 _10037_ ( .A(\ID_EX_typ [6] ), .ZN(_02409_ ) );
AND2_X1 _10038_ ( .A1(_02408_ ), .A2(_02409_ ), .ZN(_02410_ ) );
BUF_X4 _10039_ ( .A(_02410_ ), .Z(_02411_ ) );
INV_X1 _10040_ ( .A(\ID_EX_typ [5] ), .ZN(_02412_ ) );
NOR2_X1 _10041_ ( .A1(_02412_ ), .A2(\ID_EX_typ [6] ), .ZN(_02413_ ) );
AND2_X1 _10042_ ( .A1(_02413_ ), .A2(\ID_EX_typ [7] ), .ZN(_02414_ ) );
BUF_X2 _10043_ ( .A(_02414_ ), .Z(_02415_ ) );
OAI21_X1 _10044_ ( .A(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .B1(_02411_ ), .B2(_02415_ ), .ZN(_02416_ ) );
INV_X1 _10045_ ( .A(check_quest ), .ZN(_02417_ ) );
OR2_X1 _10046_ ( .A1(_02417_ ), .A2(check_assert ), .ZN(_02418_ ) );
INV_X2 _10047_ ( .A(fanout_net_5 ), .ZN(_02419_ ) );
NAND2_X2 _10048_ ( .A1(_02414_ ), .A2(_02419_ ), .ZN(_02420_ ) );
INV_X1 _10049_ ( .A(_02410_ ), .ZN(_02421_ ) );
OAI21_X1 _10050_ ( .A(_02420_ ), .B1(_02421_ ), .B2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_02422_ ) );
AOI221_X4 _10051_ ( .A(_02404_ ), .B1(_02416_ ), .B2(_02418_ ), .C1(_02422_ ), .C2(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_00096_ ) );
AND2_X1 _10052_ ( .A1(_02345_ ), .A2(\EX_LS_flag [2] ), .ZN(_02423_ ) );
NOR2_X2 _10053_ ( .A1(_02423_ ), .A2(_02327_ ), .ZN(_02424_ ) );
OAI211_X1 _10054_ ( .A(_02344_ ), .B(\EX_LS_flag [0] ), .C1(\EX_LS_flag [2] ), .C2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02425_ ) );
NAND2_X4 _10055_ ( .A1(_02424_ ), .A2(_02425_ ), .ZN(_02426_ ) );
OR4_X4 _10056_ ( .A1(\EX_LS_dest_reg [3] ), .A2(\EX_LS_dest_reg [2] ), .A3(\EX_LS_dest_reg [1] ), .A4(\EX_LS_dest_reg [0] ), .ZN(_02427_ ) );
NOR2_X2 _10057_ ( .A1(_02427_ ), .A2(\EX_LS_dest_reg [4] ), .ZN(_02428_ ) );
INV_X2 _10058_ ( .A(_02428_ ), .ZN(_02429_ ) );
INV_X4 _10059_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02430_ ) );
NAND2_X1 _10060_ ( .A1(_02430_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02431_ ) );
XNOR2_X1 _10061_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02432_ ) );
NAND4_X4 _10062_ ( .A1(_02426_ ), .A2(_02429_ ), .A3(_02431_ ), .A4(_02432_ ), .ZN(_02433_ ) );
BUF_X4 _10063_ ( .A(_02433_ ), .Z(_02434_ ) );
XNOR2_X1 _10064_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .ZN(_02435_ ) );
OAI211_X1 _10065_ ( .A(_02435_ ), .B(\myidu.fc_disenable_$_NOT__A_Y ), .C1(\ID_EX_rs1 [1] ), .C2(_02430_ ), .ZN(_02436_ ) );
XOR2_X1 _10066_ ( .A(\ID_EX_rs1 [3] ), .B(\EX_LS_dest_reg [3] ), .Z(_02437_ ) );
XOR2_X1 _10067_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .Z(_02438_ ) );
OR3_X4 _10068_ ( .A1(_02436_ ), .A2(_02437_ ), .A3(_02438_ ), .ZN(_02439_ ) );
BUF_X4 _10069_ ( .A(_02439_ ), .Z(_02440_ ) );
NOR2_X1 _10070_ ( .A1(_02434_ ), .A2(_02440_ ), .ZN(_02441_ ) );
INV_X2 _10071_ ( .A(_02441_ ), .ZN(_02442_ ) );
OR2_X1 _10072_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02443_ ) );
INV_X1 _10073_ ( .A(fanout_net_25 ), .ZN(_02444_ ) );
BUF_X4 _10074_ ( .A(_02444_ ), .Z(_02445_ ) );
BUF_X4 _10075_ ( .A(_02445_ ), .Z(_02446_ ) );
BUF_X4 _10076_ ( .A(_02446_ ), .Z(_02447_ ) );
BUF_X4 _10077_ ( .A(_02447_ ), .Z(_02448_ ) );
BUF_X4 _10078_ ( .A(_02448_ ), .Z(_02449_ ) );
BUF_X2 _10079_ ( .A(_02449_ ), .Z(_02450_ ) );
INV_X1 _10080_ ( .A(fanout_net_17 ), .ZN(_02451_ ) );
BUF_X4 _10081_ ( .A(_02451_ ), .Z(_02452_ ) );
BUF_X4 _10082_ ( .A(_02452_ ), .Z(_02453_ ) );
BUF_X4 _10083_ ( .A(_02453_ ), .Z(_02454_ ) );
BUF_X4 _10084_ ( .A(_02454_ ), .Z(_02455_ ) );
BUF_X4 _10085_ ( .A(_02455_ ), .Z(_02456_ ) );
OAI211_X1 _10086_ ( .A(_02443_ ), .B(_02450_ ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02457_ ) );
OR2_X1 _10087_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02458_ ) );
OAI211_X1 _10088_ ( .A(_02458_ ), .B(fanout_net_25 ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02459_ ) );
INV_X1 _10089_ ( .A(fanout_net_28 ), .ZN(_02460_ ) );
BUF_X4 _10090_ ( .A(_02460_ ), .Z(_02461_ ) );
BUF_X4 _10091_ ( .A(_02461_ ), .Z(_02462_ ) );
BUF_X4 _10092_ ( .A(_02462_ ), .Z(_02463_ ) );
BUF_X4 _10093_ ( .A(_02463_ ), .Z(_02464_ ) );
BUF_X4 _10094_ ( .A(_02464_ ), .Z(_02465_ ) );
NAND3_X1 _10095_ ( .A1(_02457_ ), .A2(_02459_ ), .A3(_02465_ ), .ZN(_02466_ ) );
MUX2_X1 _10096_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02467_ ) );
MUX2_X1 _10097_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02468_ ) );
BUF_X4 _10098_ ( .A(_02447_ ), .Z(_02469_ ) );
BUF_X4 _10099_ ( .A(_02469_ ), .Z(_02470_ ) );
MUX2_X1 _10100_ ( .A(_02467_ ), .B(_02468_ ), .S(_02470_ ), .Z(_02471_ ) );
OAI211_X1 _10101_ ( .A(fanout_net_30 ), .B(_02466_ ), .C1(_02471_ ), .C2(_02465_ ), .ZN(_02472_ ) );
NOR2_X1 _10102_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02473_ ) );
INV_X1 _10103_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02474_ ) );
AOI211_X1 _10104_ ( .A(_02449_ ), .B(_02473_ ), .C1(fanout_net_17 ), .C2(_02474_ ), .ZN(_02475_ ) );
MUX2_X1 _10105_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02476_ ) );
AOI21_X1 _10106_ ( .A(_02475_ ), .B1(_02470_ ), .B2(_02476_ ), .ZN(_02477_ ) );
MUX2_X1 _10107_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02478_ ) );
AND2_X1 _10108_ ( .A1(_02478_ ), .A2(_02449_ ), .ZN(_02479_ ) );
MUX2_X1 _10109_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02480_ ) );
AOI21_X1 _10110_ ( .A(_02479_ ), .B1(fanout_net_25 ), .B2(_02480_ ), .ZN(_02481_ ) );
MUX2_X1 _10111_ ( .A(_02477_ ), .B(_02481_ ), .S(fanout_net_28 ), .Z(_02482_ ) );
OAI211_X1 _10112_ ( .A(_02442_ ), .B(_02472_ ), .C1(fanout_net_30 ), .C2(_02482_ ), .ZN(_02483_ ) );
INV_X1 _10113_ ( .A(\ID_EX_imm [27] ), .ZN(_02484_ ) );
BUF_X8 _10114_ ( .A(_02434_ ), .Z(_02485_ ) );
BUF_X2 _10115_ ( .A(_02485_ ), .Z(_02486_ ) );
BUF_X2 _10116_ ( .A(_02486_ ), .Z(_02487_ ) );
CLKBUF_X2 _10117_ ( .A(_02487_ ), .Z(_02488_ ) );
BUF_X8 _10118_ ( .A(_02440_ ), .Z(_02489_ ) );
BUF_X2 _10119_ ( .A(_02489_ ), .Z(_02490_ ) );
BUF_X2 _10120_ ( .A(_02490_ ), .Z(_02491_ ) );
CLKBUF_X2 _10121_ ( .A(_02491_ ), .Z(_02492_ ) );
OR3_X1 _10122_ ( .A1(_02488_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02492_ ), .ZN(_02493_ ) );
AND3_X1 _10123_ ( .A1(_02483_ ), .A2(_02484_ ), .A3(_02493_ ), .ZN(_02494_ ) );
AOI21_X1 _10124_ ( .A(_02484_ ), .B1(_02483_ ), .B2(_02493_ ), .ZN(_02495_ ) );
NOR2_X1 _10125_ ( .A1(_02494_ ), .A2(_02495_ ), .ZN(_02496_ ) );
INV_X1 _10126_ ( .A(fanout_net_30 ), .ZN(_02497_ ) );
BUF_X4 _10127_ ( .A(_02497_ ), .Z(_02498_ ) );
BUF_X4 _10128_ ( .A(_02498_ ), .Z(_02499_ ) );
OR2_X1 _10129_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02500_ ) );
BUF_X4 _10130_ ( .A(_02454_ ), .Z(_02501_ ) );
OAI211_X1 _10131_ ( .A(_02500_ ), .B(_02469_ ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02502_ ) );
OR2_X1 _10132_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02503_ ) );
OAI211_X1 _10133_ ( .A(_02503_ ), .B(fanout_net_25 ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02504_ ) );
NAND3_X1 _10134_ ( .A1(_02502_ ), .A2(_02504_ ), .A3(fanout_net_28 ), .ZN(_02505_ ) );
MUX2_X1 _10135_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02506_ ) );
MUX2_X1 _10136_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02507_ ) );
MUX2_X1 _10137_ ( .A(_02506_ ), .B(_02507_ ), .S(_02448_ ), .Z(_02508_ ) );
OAI211_X1 _10138_ ( .A(_02499_ ), .B(_02505_ ), .C1(_02508_ ), .C2(fanout_net_28 ), .ZN(_02509_ ) );
MUX2_X1 _10139_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02510_ ) );
MUX2_X1 _10140_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02511_ ) );
MUX2_X1 _10141_ ( .A(_02510_ ), .B(_02511_ ), .S(fanout_net_28 ), .Z(_02512_ ) );
AND2_X1 _10142_ ( .A1(_02512_ ), .A2(fanout_net_25 ), .ZN(_02513_ ) );
MUX2_X1 _10143_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02514_ ) );
MUX2_X1 _10144_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02515_ ) );
MUX2_X1 _10145_ ( .A(_02514_ ), .B(_02515_ ), .S(fanout_net_28 ), .Z(_02516_ ) );
AND2_X1 _10146_ ( .A1(_02516_ ), .A2(_02449_ ), .ZN(_02517_ ) );
OAI21_X1 _10147_ ( .A(fanout_net_30 ), .B1(_02513_ ), .B2(_02517_ ), .ZN(_02518_ ) );
NAND3_X1 _10148_ ( .A1(_02442_ ), .A2(_02509_ ), .A3(_02518_ ), .ZN(_02519_ ) );
OR3_X1 _10149_ ( .A1(_02486_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02490_ ), .ZN(_02520_ ) );
NAND2_X1 _10150_ ( .A1(_02519_ ), .A2(_02520_ ), .ZN(_02521_ ) );
BUF_X2 _10151_ ( .A(_02521_ ), .Z(_02522_ ) );
INV_X1 _10152_ ( .A(\ID_EX_imm [22] ), .ZN(_02523_ ) );
XNOR2_X1 _10153_ ( .A(_02522_ ), .B(_02523_ ), .ZN(_02524_ ) );
OR2_X1 _10154_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02525_ ) );
OAI211_X1 _10155_ ( .A(_02525_ ), .B(_02448_ ), .C1(_02454_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02526_ ) );
OR2_X1 _10156_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02527_ ) );
OAI211_X1 _10157_ ( .A(_02527_ ), .B(fanout_net_25 ), .C1(_02454_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02528_ ) );
NAND3_X1 _10158_ ( .A1(_02526_ ), .A2(_02528_ ), .A3(fanout_net_28 ), .ZN(_02529_ ) );
MUX2_X1 _10159_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02530_ ) );
MUX2_X1 _10160_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02531_ ) );
MUX2_X1 _10161_ ( .A(_02530_ ), .B(_02531_ ), .S(_02447_ ), .Z(_02532_ ) );
OAI211_X1 _10162_ ( .A(_02499_ ), .B(_02529_ ), .C1(_02532_ ), .C2(fanout_net_28 ), .ZN(_02533_ ) );
MUX2_X1 _10163_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02534_ ) );
MUX2_X1 _10164_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02535_ ) );
MUX2_X1 _10165_ ( .A(_02534_ ), .B(_02535_ ), .S(fanout_net_28 ), .Z(_02536_ ) );
AND2_X1 _10166_ ( .A1(_02536_ ), .A2(fanout_net_25 ), .ZN(_02537_ ) );
MUX2_X1 _10167_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02538_ ) );
MUX2_X1 _10168_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02539_ ) );
MUX2_X1 _10169_ ( .A(_02538_ ), .B(_02539_ ), .S(fanout_net_28 ), .Z(_02540_ ) );
AND2_X1 _10170_ ( .A1(_02540_ ), .A2(_02469_ ), .ZN(_02541_ ) );
OAI21_X1 _10171_ ( .A(fanout_net_30 ), .B1(_02537_ ), .B2(_02541_ ), .ZN(_02542_ ) );
NAND3_X1 _10172_ ( .A1(_02442_ ), .A2(_02533_ ), .A3(_02542_ ), .ZN(_02543_ ) );
INV_X1 _10173_ ( .A(\ID_EX_imm [23] ), .ZN(_02544_ ) );
OR3_X1 _10174_ ( .A1(_02486_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02490_ ), .ZN(_02545_ ) );
NAND3_X1 _10175_ ( .A1(_02543_ ), .A2(_02544_ ), .A3(_02545_ ), .ZN(_02546_ ) );
NAND2_X1 _10176_ ( .A1(_02543_ ), .A2(_02545_ ), .ZN(_02547_ ) );
BUF_X4 _10177_ ( .A(_02547_ ), .Z(_02548_ ) );
NAND2_X1 _10178_ ( .A1(_02548_ ), .A2(\ID_EX_imm [23] ), .ZN(_02549_ ) );
AND3_X1 _10179_ ( .A1(_02524_ ), .A2(_02546_ ), .A3(_02549_ ), .ZN(_02550_ ) );
OR3_X1 _10180_ ( .A1(_02486_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02490_ ), .ZN(_02551_ ) );
OR2_X1 _10181_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02552_ ) );
BUF_X4 _10182_ ( .A(_02454_ ), .Z(_02553_ ) );
OAI211_X1 _10183_ ( .A(_02552_ ), .B(_02448_ ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02554_ ) );
OR2_X1 _10184_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02555_ ) );
OAI211_X1 _10185_ ( .A(_02555_ ), .B(fanout_net_25 ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02556_ ) );
NAND3_X1 _10186_ ( .A1(_02554_ ), .A2(_02556_ ), .A3(_02463_ ), .ZN(_02557_ ) );
MUX2_X1 _10187_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02558_ ) );
MUX2_X1 _10188_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02559_ ) );
MUX2_X1 _10189_ ( .A(_02558_ ), .B(_02559_ ), .S(_02448_ ), .Z(_02560_ ) );
OAI211_X1 _10190_ ( .A(fanout_net_30 ), .B(_02557_ ), .C1(_02560_ ), .C2(_02464_ ), .ZN(_02561_ ) );
OR2_X1 _10191_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02562_ ) );
OAI211_X1 _10192_ ( .A(_02562_ ), .B(_02469_ ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02563_ ) );
OR2_X1 _10193_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02564_ ) );
OAI211_X1 _10194_ ( .A(_02564_ ), .B(fanout_net_25 ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02565_ ) );
NAND3_X1 _10195_ ( .A1(_02563_ ), .A2(_02565_ ), .A3(_02464_ ), .ZN(_02566_ ) );
OR2_X1 _10196_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02567_ ) );
OAI211_X1 _10197_ ( .A(_02567_ ), .B(_02448_ ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02568_ ) );
OR2_X1 _10198_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02569_ ) );
OAI211_X1 _10199_ ( .A(_02569_ ), .B(fanout_net_25 ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02570_ ) );
NAND3_X1 _10200_ ( .A1(_02568_ ), .A2(_02570_ ), .A3(fanout_net_28 ), .ZN(_02571_ ) );
NAND3_X1 _10201_ ( .A1(_02566_ ), .A2(_02571_ ), .A3(_02499_ ), .ZN(_02572_ ) );
OAI211_X1 _10202_ ( .A(_02561_ ), .B(_02572_ ), .C1(_02487_ ), .C2(_02491_ ), .ZN(_02573_ ) );
NAND2_X1 _10203_ ( .A1(_02551_ ), .A2(_02573_ ), .ZN(_02574_ ) );
BUF_X4 _10204_ ( .A(_02574_ ), .Z(_02575_ ) );
INV_X1 _10205_ ( .A(\ID_EX_imm [21] ), .ZN(_02576_ ) );
XNOR2_X1 _10206_ ( .A(_02575_ ), .B(_02576_ ), .ZN(_02577_ ) );
OR3_X1 _10207_ ( .A1(_02487_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02491_ ), .ZN(_02578_ ) );
OR2_X1 _10208_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02579_ ) );
OAI211_X1 _10209_ ( .A(_02579_ ), .B(_02469_ ), .C1(_02455_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02580_ ) );
OR2_X1 _10210_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02581_ ) );
OAI211_X1 _10211_ ( .A(_02581_ ), .B(fanout_net_25 ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02582_ ) );
NAND3_X1 _10212_ ( .A1(_02580_ ), .A2(_02582_ ), .A3(_02464_ ), .ZN(_02583_ ) );
MUX2_X1 _10213_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02584_ ) );
MUX2_X1 _10214_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02585_ ) );
MUX2_X1 _10215_ ( .A(_02584_ ), .B(_02585_ ), .S(_02469_ ), .Z(_02586_ ) );
OAI211_X1 _10216_ ( .A(_02499_ ), .B(_02583_ ), .C1(_02586_ ), .C2(_02464_ ), .ZN(_02587_ ) );
OR2_X1 _10217_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02588_ ) );
OAI211_X1 _10218_ ( .A(_02588_ ), .B(fanout_net_25 ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02589_ ) );
OR2_X1 _10219_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02590_ ) );
OAI211_X1 _10220_ ( .A(_02590_ ), .B(_02469_ ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02591_ ) );
NAND3_X1 _10221_ ( .A1(_02589_ ), .A2(_02591_ ), .A3(fanout_net_28 ), .ZN(_02592_ ) );
MUX2_X1 _10222_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02593_ ) );
MUX2_X1 _10223_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02594_ ) );
MUX2_X1 _10224_ ( .A(_02593_ ), .B(_02594_ ), .S(fanout_net_25 ), .Z(_02595_ ) );
OAI211_X1 _10225_ ( .A(fanout_net_30 ), .B(_02592_ ), .C1(_02595_ ), .C2(fanout_net_28 ), .ZN(_02596_ ) );
OAI211_X1 _10226_ ( .A(_02587_ ), .B(_02596_ ), .C1(_02487_ ), .C2(_02491_ ), .ZN(_02597_ ) );
NAND2_X1 _10227_ ( .A1(_02578_ ), .A2(_02597_ ), .ZN(_02598_ ) );
INV_X1 _10228_ ( .A(\ID_EX_imm [20] ), .ZN(_02599_ ) );
XNOR2_X1 _10229_ ( .A(_02598_ ), .B(_02599_ ), .ZN(_02600_ ) );
AND2_X1 _10230_ ( .A1(_02577_ ), .A2(_02600_ ), .ZN(_02601_ ) );
AND2_X1 _10231_ ( .A1(_02550_ ), .A2(_02601_ ), .ZN(_02602_ ) );
INV_X1 _10232_ ( .A(_02602_ ), .ZN(_02603_ ) );
OR3_X1 _10233_ ( .A1(_02486_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02490_ ), .ZN(_02604_ ) );
OR2_X1 _10234_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02605_ ) );
OAI211_X1 _10235_ ( .A(_02605_ ), .B(_02448_ ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02606_ ) );
OR2_X1 _10236_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02607_ ) );
OAI211_X1 _10237_ ( .A(_02607_ ), .B(fanout_net_25 ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02608_ ) );
NAND3_X1 _10238_ ( .A1(_02606_ ), .A2(_02608_ ), .A3(_02463_ ), .ZN(_02609_ ) );
MUX2_X1 _10239_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02610_ ) );
MUX2_X1 _10240_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02611_ ) );
MUX2_X1 _10241_ ( .A(_02610_ ), .B(_02611_ ), .S(_02448_ ), .Z(_02612_ ) );
OAI211_X1 _10242_ ( .A(fanout_net_30 ), .B(_02609_ ), .C1(_02612_ ), .C2(_02464_ ), .ZN(_02613_ ) );
OR2_X1 _10243_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02614_ ) );
OAI211_X1 _10244_ ( .A(_02614_ ), .B(_02448_ ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02615_ ) );
OR2_X1 _10245_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02616_ ) );
OAI211_X1 _10246_ ( .A(_02616_ ), .B(fanout_net_25 ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02617_ ) );
AOI21_X1 _10247_ ( .A(_02463_ ), .B1(_02615_ ), .B2(_02617_ ), .ZN(_02618_ ) );
OR2_X1 _10248_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02619_ ) );
OAI211_X1 _10249_ ( .A(_02619_ ), .B(_02448_ ), .C1(_02553_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02620_ ) );
OR2_X1 _10250_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02621_ ) );
OAI211_X1 _10251_ ( .A(_02621_ ), .B(fanout_net_25 ), .C1(_02454_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02622_ ) );
AOI21_X1 _10252_ ( .A(fanout_net_28 ), .B1(_02620_ ), .B2(_02622_ ), .ZN(_02623_ ) );
OAI21_X1 _10253_ ( .A(_02499_ ), .B1(_02618_ ), .B2(_02623_ ), .ZN(_02624_ ) );
OAI211_X1 _10254_ ( .A(_02613_ ), .B(_02624_ ), .C1(_02487_ ), .C2(_02491_ ), .ZN(_02625_ ) );
NAND2_X2 _10255_ ( .A1(_02604_ ), .A2(_02625_ ), .ZN(_02626_ ) );
INV_X1 _10256_ ( .A(\ID_EX_imm [18] ), .ZN(_02627_ ) );
XNOR2_X1 _10257_ ( .A(_02626_ ), .B(_02627_ ), .ZN(_02628_ ) );
CLKBUF_X3 _10258_ ( .A(_02434_ ), .Z(_02629_ ) );
CLKBUF_X2 _10259_ ( .A(_02440_ ), .Z(_02630_ ) );
OR3_X1 _10260_ ( .A1(_02629_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02630_ ), .ZN(_02631_ ) );
OR2_X1 _10261_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02632_ ) );
BUF_X4 _10262_ ( .A(_02452_ ), .Z(_02633_ ) );
BUF_X4 _10263_ ( .A(_02633_ ), .Z(_02634_ ) );
OAI211_X1 _10264_ ( .A(_02632_ ), .B(_02447_ ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02635_ ) );
OR2_X1 _10265_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02636_ ) );
OAI211_X1 _10266_ ( .A(_02636_ ), .B(fanout_net_25 ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02637_ ) );
NAND3_X1 _10267_ ( .A1(_02635_ ), .A2(_02637_ ), .A3(_02462_ ), .ZN(_02638_ ) );
MUX2_X1 _10268_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02639_ ) );
MUX2_X1 _10269_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02640_ ) );
BUF_X4 _10270_ ( .A(_02445_ ), .Z(_02641_ ) );
BUF_X4 _10271_ ( .A(_02641_ ), .Z(_02642_ ) );
MUX2_X1 _10272_ ( .A(_02639_ ), .B(_02640_ ), .S(_02642_ ), .Z(_02643_ ) );
OAI211_X1 _10273_ ( .A(_02499_ ), .B(_02638_ ), .C1(_02643_ ), .C2(_02463_ ), .ZN(_02644_ ) );
OR2_X1 _10274_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02645_ ) );
OAI211_X1 _10275_ ( .A(_02645_ ), .B(fanout_net_25 ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02646_ ) );
OR2_X1 _10276_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02647_ ) );
OAI211_X1 _10277_ ( .A(_02647_ ), .B(_02447_ ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02648_ ) );
NAND3_X1 _10278_ ( .A1(_02646_ ), .A2(_02648_ ), .A3(fanout_net_28 ), .ZN(_02649_ ) );
MUX2_X1 _10279_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02650_ ) );
MUX2_X1 _10280_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02651_ ) );
MUX2_X1 _10281_ ( .A(_02650_ ), .B(_02651_ ), .S(fanout_net_25 ), .Z(_02652_ ) );
OAI211_X1 _10282_ ( .A(fanout_net_30 ), .B(_02649_ ), .C1(_02652_ ), .C2(fanout_net_28 ), .ZN(_02653_ ) );
OAI211_X1 _10283_ ( .A(_02644_ ), .B(_02653_ ), .C1(_02486_ ), .C2(_02490_ ), .ZN(_02654_ ) );
NAND2_X2 _10284_ ( .A1(_02631_ ), .A2(_02654_ ), .ZN(_02655_ ) );
INV_X1 _10285_ ( .A(\ID_EX_imm [19] ), .ZN(_02656_ ) );
XNOR2_X1 _10286_ ( .A(_02655_ ), .B(_02656_ ), .ZN(_02657_ ) );
AND2_X1 _10287_ ( .A1(_02628_ ), .A2(_02657_ ), .ZN(_02658_ ) );
OR3_X1 _10288_ ( .A1(_02629_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02630_ ), .ZN(_02659_ ) );
OR2_X1 _10289_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02660_ ) );
BUF_X4 _10290_ ( .A(_02451_ ), .Z(_02661_ ) );
BUF_X4 _10291_ ( .A(_02661_ ), .Z(_02662_ ) );
BUF_X4 _10292_ ( .A(_02662_ ), .Z(_02663_ ) );
OAI211_X1 _10293_ ( .A(_02660_ ), .B(_02642_ ), .C1(_02663_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02664_ ) );
OR2_X1 _10294_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02665_ ) );
OAI211_X1 _10295_ ( .A(_02665_ ), .B(fanout_net_25 ), .C1(_02663_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02666_ ) );
NAND3_X1 _10296_ ( .A1(_02664_ ), .A2(_02666_ ), .A3(_02462_ ), .ZN(_02667_ ) );
MUX2_X1 _10297_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02668_ ) );
MUX2_X1 _10298_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02669_ ) );
MUX2_X1 _10299_ ( .A(_02668_ ), .B(_02669_ ), .S(_02446_ ), .Z(_02670_ ) );
OAI211_X1 _10300_ ( .A(_02498_ ), .B(_02667_ ), .C1(_02670_ ), .C2(_02463_ ), .ZN(_02671_ ) );
OR2_X1 _10301_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02672_ ) );
OAI211_X1 _10302_ ( .A(_02672_ ), .B(fanout_net_25 ), .C1(_02663_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02673_ ) );
OR2_X1 _10303_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02674_ ) );
OAI211_X1 _10304_ ( .A(_02674_ ), .B(_02446_ ), .C1(_02663_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02675_ ) );
NAND3_X1 _10305_ ( .A1(_02673_ ), .A2(_02675_ ), .A3(fanout_net_28 ), .ZN(_02676_ ) );
MUX2_X1 _10306_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02677_ ) );
MUX2_X1 _10307_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02678_ ) );
MUX2_X1 _10308_ ( .A(_02677_ ), .B(_02678_ ), .S(fanout_net_25 ), .Z(_02679_ ) );
OAI211_X1 _10309_ ( .A(fanout_net_30 ), .B(_02676_ ), .C1(_02679_ ), .C2(fanout_net_28 ), .ZN(_02680_ ) );
OAI211_X1 _10310_ ( .A(_02671_ ), .B(_02680_ ), .C1(_02486_ ), .C2(_02490_ ), .ZN(_02681_ ) );
NAND2_X1 _10311_ ( .A1(_02659_ ), .A2(_02681_ ), .ZN(_02682_ ) );
INV_X1 _10312_ ( .A(\ID_EX_imm [17] ), .ZN(_02683_ ) );
XNOR2_X1 _10313_ ( .A(_02682_ ), .B(_02683_ ), .ZN(_02684_ ) );
OR3_X1 _10314_ ( .A1(_02487_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02491_ ), .ZN(_02685_ ) );
BUF_X2 _10315_ ( .A(_02499_ ), .Z(_02686_ ) );
OR2_X1 _10316_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02687_ ) );
OAI211_X1 _10317_ ( .A(_02687_ ), .B(_02449_ ), .C1(_02455_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02688_ ) );
OR2_X1 _10318_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02689_ ) );
OAI211_X1 _10319_ ( .A(_02689_ ), .B(fanout_net_25 ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02690_ ) );
NAND3_X1 _10320_ ( .A1(_02688_ ), .A2(_02690_ ), .A3(_02464_ ), .ZN(_02691_ ) );
MUX2_X1 _10321_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02692_ ) );
MUX2_X1 _10322_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02693_ ) );
MUX2_X1 _10323_ ( .A(_02692_ ), .B(_02693_ ), .S(_02469_ ), .Z(_02694_ ) );
OAI211_X1 _10324_ ( .A(_02686_ ), .B(_02691_ ), .C1(_02694_ ), .C2(_02464_ ), .ZN(_02695_ ) );
OR2_X1 _10325_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02696_ ) );
OAI211_X1 _10326_ ( .A(_02696_ ), .B(fanout_net_25 ), .C1(_02455_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02697_ ) );
OR2_X1 _10327_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02698_ ) );
OAI211_X1 _10328_ ( .A(_02698_ ), .B(_02469_ ), .C1(_02501_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02699_ ) );
NAND3_X1 _10329_ ( .A1(_02697_ ), .A2(_02699_ ), .A3(fanout_net_28 ), .ZN(_02700_ ) );
MUX2_X1 _10330_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02701_ ) );
MUX2_X1 _10331_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02702_ ) );
MUX2_X1 _10332_ ( .A(_02701_ ), .B(_02702_ ), .S(fanout_net_25 ), .Z(_02703_ ) );
OAI211_X1 _10333_ ( .A(fanout_net_30 ), .B(_02700_ ), .C1(_02703_ ), .C2(fanout_net_28 ), .ZN(_02704_ ) );
OAI211_X1 _10334_ ( .A(_02695_ ), .B(_02704_ ), .C1(_02487_ ), .C2(_02491_ ), .ZN(_02705_ ) );
NAND2_X1 _10335_ ( .A1(_02685_ ), .A2(_02705_ ), .ZN(_02706_ ) );
INV_X1 _10336_ ( .A(\ID_EX_imm [16] ), .ZN(_02707_ ) );
XNOR2_X1 _10337_ ( .A(_02706_ ), .B(_02707_ ), .ZN(_02708_ ) );
NAND3_X1 _10338_ ( .A1(_02658_ ), .A2(_02684_ ), .A3(_02708_ ), .ZN(_02709_ ) );
OR2_X1 _10339_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02710_ ) );
BUF_X4 _10340_ ( .A(_02445_ ), .Z(_02711_ ) );
OAI211_X1 _10341_ ( .A(_02710_ ), .B(_02711_ ), .C1(_02662_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02712_ ) );
OR2_X1 _10342_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02713_ ) );
OAI211_X1 _10343_ ( .A(_02713_ ), .B(fanout_net_25 ), .C1(_02662_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02714_ ) );
BUF_X4 _10344_ ( .A(_02461_ ), .Z(_02715_ ) );
NAND3_X1 _10345_ ( .A1(_02712_ ), .A2(_02714_ ), .A3(_02715_ ), .ZN(_02716_ ) );
MUX2_X1 _10346_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02717_ ) );
MUX2_X1 _10347_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02718_ ) );
MUX2_X1 _10348_ ( .A(_02717_ ), .B(_02718_ ), .S(_02711_ ), .Z(_02719_ ) );
OAI211_X1 _10349_ ( .A(fanout_net_30 ), .B(_02716_ ), .C1(_02719_ ), .C2(_02715_ ), .ZN(_02720_ ) );
MUX2_X1 _10350_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02721_ ) );
AND2_X1 _10351_ ( .A1(_02721_ ), .A2(fanout_net_25 ), .ZN(_02722_ ) );
MUX2_X1 _10352_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02723_ ) );
AOI21_X1 _10353_ ( .A(_02722_ ), .B1(_02711_ ), .B2(_02723_ ), .ZN(_02724_ ) );
NOR2_X1 _10354_ ( .A1(_02724_ ), .A2(_02461_ ), .ZN(_02725_ ) );
MUX2_X1 _10355_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02726_ ) );
MUX2_X1 _10356_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02727_ ) );
MUX2_X1 _10357_ ( .A(_02726_ ), .B(_02727_ ), .S(_02445_ ), .Z(_02728_ ) );
AOI21_X1 _10358_ ( .A(_02725_ ), .B1(_02715_ ), .B2(_02728_ ), .ZN(_02729_ ) );
OAI211_X1 _10359_ ( .A(_02442_ ), .B(_02720_ ), .C1(fanout_net_30 ), .C2(_02729_ ), .ZN(_02730_ ) );
OR3_X1 _10360_ ( .A1(_02434_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02440_ ), .ZN(_02731_ ) );
NAND2_X2 _10361_ ( .A1(_02730_ ), .A2(_02731_ ), .ZN(_02732_ ) );
INV_X1 _10362_ ( .A(\ID_EX_imm [3] ), .ZN(_02733_ ) );
XNOR2_X1 _10363_ ( .A(_02732_ ), .B(_02733_ ), .ZN(_02734_ ) );
OR3_X1 _10364_ ( .A1(_02433_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02439_ ), .ZN(_02735_ ) );
OR2_X1 _10365_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02736_ ) );
OAI211_X1 _10366_ ( .A(_02736_ ), .B(_02444_ ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02737_ ) );
OR2_X1 _10367_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02738_ ) );
OAI211_X1 _10368_ ( .A(_02738_ ), .B(fanout_net_25 ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02739_ ) );
NAND3_X1 _10369_ ( .A1(_02737_ ), .A2(_02739_ ), .A3(_02460_ ), .ZN(_02740_ ) );
MUX2_X1 _10370_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02741_ ) );
MUX2_X1 _10371_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02742_ ) );
MUX2_X1 _10372_ ( .A(_02741_ ), .B(_02742_ ), .S(_02444_ ), .Z(_02743_ ) );
OAI211_X1 _10373_ ( .A(_02497_ ), .B(_02740_ ), .C1(_02743_ ), .C2(_02461_ ), .ZN(_02744_ ) );
OR2_X1 _10374_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02745_ ) );
OAI211_X1 _10375_ ( .A(_02745_ ), .B(fanout_net_25 ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02746_ ) );
OR2_X1 _10376_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02747_ ) );
OAI211_X1 _10377_ ( .A(_02747_ ), .B(_02444_ ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02748_ ) );
NAND3_X1 _10378_ ( .A1(_02746_ ), .A2(_02748_ ), .A3(fanout_net_28 ), .ZN(_02749_ ) );
MUX2_X1 _10379_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02750_ ) );
MUX2_X1 _10380_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02751_ ) );
MUX2_X1 _10381_ ( .A(_02750_ ), .B(_02751_ ), .S(fanout_net_25 ), .Z(_02752_ ) );
OAI211_X1 _10382_ ( .A(fanout_net_30 ), .B(_02749_ ), .C1(_02752_ ), .C2(fanout_net_28 ), .ZN(_02753_ ) );
OAI211_X1 _10383_ ( .A(_02744_ ), .B(_02753_ ), .C1(_02434_ ), .C2(_02440_ ), .ZN(_02754_ ) );
NAND2_X1 _10384_ ( .A1(_02735_ ), .A2(_02754_ ), .ZN(_02755_ ) );
INV_X1 _10385_ ( .A(\ID_EX_imm [2] ), .ZN(_02756_ ) );
XNOR2_X1 _10386_ ( .A(_02755_ ), .B(_02756_ ), .ZN(_02757_ ) );
INV_X1 _10387_ ( .A(_02757_ ), .ZN(_02758_ ) );
OR3_X4 _10388_ ( .A1(_02434_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02440_ ), .ZN(_02759_ ) );
OR2_X1 _10389_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(fanout_net_20 ), .ZN(_02760_ ) );
OAI211_X1 _10390_ ( .A(_02760_ ), .B(_02445_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_02661_ ), .ZN(_02761_ ) );
OR2_X1 _10391_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02762_ ) );
OAI211_X1 _10392_ ( .A(_02762_ ), .B(fanout_net_26 ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02763_ ) );
NAND3_X1 _10393_ ( .A1(_02761_ ), .A2(_02763_ ), .A3(_02461_ ), .ZN(_02764_ ) );
MUX2_X1 _10394_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02765_ ) );
MUX2_X1 _10395_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02766_ ) );
MUX2_X1 _10396_ ( .A(_02765_ ), .B(_02766_ ), .S(_02444_ ), .Z(_02767_ ) );
OAI211_X1 _10397_ ( .A(_02497_ ), .B(_02764_ ), .C1(_02767_ ), .C2(_02461_ ), .ZN(_02768_ ) );
OR2_X1 _10398_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02769_ ) );
OAI211_X1 _10399_ ( .A(_02769_ ), .B(fanout_net_26 ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02770_ ) );
OR2_X1 _10400_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02771_ ) );
OAI211_X1 _10401_ ( .A(_02771_ ), .B(_02444_ ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02772_ ) );
NAND3_X1 _10402_ ( .A1(_02770_ ), .A2(_02772_ ), .A3(fanout_net_28 ), .ZN(_02773_ ) );
MUX2_X1 _10403_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02774_ ) );
MUX2_X1 _10404_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02775_ ) );
MUX2_X1 _10405_ ( .A(_02774_ ), .B(_02775_ ), .S(fanout_net_26 ), .Z(_02776_ ) );
OAI211_X1 _10406_ ( .A(fanout_net_30 ), .B(_02773_ ), .C1(_02776_ ), .C2(fanout_net_28 ), .ZN(_02777_ ) );
OAI211_X1 _10407_ ( .A(_02768_ ), .B(_02777_ ), .C1(_02434_ ), .C2(_02440_ ), .ZN(_02778_ ) );
NAND2_X2 _10408_ ( .A1(_02759_ ), .A2(_02778_ ), .ZN(_02779_ ) );
INV_X1 _10409_ ( .A(\ID_EX_imm [1] ), .ZN(_02780_ ) );
XNOR2_X1 _10410_ ( .A(_02779_ ), .B(_02780_ ), .ZN(_02781_ ) );
INV_X1 _10411_ ( .A(\ID_EX_imm [0] ), .ZN(_02782_ ) );
OR3_X1 _10412_ ( .A1(_02434_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_02440_ ), .ZN(_02783_ ) );
OR2_X1 _10413_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02784_ ) );
OAI211_X1 _10414_ ( .A(_02784_ ), .B(_02711_ ), .C1(_02662_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02785_ ) );
OR2_X1 _10415_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02786_ ) );
OAI211_X1 _10416_ ( .A(_02786_ ), .B(fanout_net_26 ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02787_ ) );
NAND3_X1 _10417_ ( .A1(_02785_ ), .A2(_02787_ ), .A3(_02461_ ), .ZN(_02788_ ) );
MUX2_X1 _10418_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02789_ ) );
MUX2_X1 _10419_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02790_ ) );
MUX2_X1 _10420_ ( .A(_02789_ ), .B(_02790_ ), .S(_02445_ ), .Z(_02791_ ) );
OAI211_X1 _10421_ ( .A(_02497_ ), .B(_02788_ ), .C1(_02791_ ), .C2(_02715_ ), .ZN(_02792_ ) );
OR2_X1 _10422_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02793_ ) );
OAI211_X1 _10423_ ( .A(_02793_ ), .B(fanout_net_26 ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02794_ ) );
OR2_X1 _10424_ ( .A1(fanout_net_20 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02795_ ) );
OAI211_X1 _10425_ ( .A(_02795_ ), .B(_02711_ ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02796_ ) );
NAND3_X1 _10426_ ( .A1(_02794_ ), .A2(_02796_ ), .A3(fanout_net_28 ), .ZN(_02797_ ) );
MUX2_X1 _10427_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02798_ ) );
MUX2_X1 _10428_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02799_ ) );
MUX2_X1 _10429_ ( .A(_02798_ ), .B(_02799_ ), .S(fanout_net_26 ), .Z(_02800_ ) );
OAI211_X1 _10430_ ( .A(fanout_net_30 ), .B(_02797_ ), .C1(_02800_ ), .C2(fanout_net_28 ), .ZN(_02801_ ) );
OAI211_X1 _10431_ ( .A(_02792_ ), .B(_02801_ ), .C1(_02485_ ), .C2(_02489_ ), .ZN(_02802_ ) );
AOI21_X1 _10432_ ( .A(_02782_ ), .B1(_02783_ ), .B2(_02802_ ), .ZN(_02803_ ) );
NAND2_X1 _10433_ ( .A1(_02781_ ), .A2(_02803_ ), .ZN(_02804_ ) );
INV_X1 _10434_ ( .A(_02779_ ), .ZN(_02805_ ) );
OR2_X1 _10435_ ( .A1(_02805_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02806_ ) );
AOI21_X4 _10436_ ( .A(_02758_ ), .B1(_02804_ ), .B2(_02806_ ), .ZN(_02807_ ) );
AOI21_X1 _10437_ ( .A(_02756_ ), .B1(_02735_ ), .B2(_02754_ ), .ZN(_02808_ ) );
OAI21_X2 _10438_ ( .A(_02734_ ), .B1(_02807_ ), .B2(_02808_ ), .ZN(_02809_ ) );
INV_X1 _10439_ ( .A(_02732_ ), .ZN(_02810_ ) );
OR2_X1 _10440_ ( .A1(_02810_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02811_ ) );
AND2_X2 _10441_ ( .A1(_02809_ ), .A2(_02811_ ), .ZN(_02812_ ) );
OR3_X1 _10442_ ( .A1(_02485_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02489_ ), .ZN(_02813_ ) );
OR2_X1 _10443_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02814_ ) );
OAI211_X1 _10444_ ( .A(_02814_ ), .B(_02446_ ), .C1(_02453_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02815_ ) );
OR2_X1 _10445_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02816_ ) );
OAI211_X1 _10446_ ( .A(_02816_ ), .B(fanout_net_26 ), .C1(_02633_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02817_ ) );
NAND3_X1 _10447_ ( .A1(_02815_ ), .A2(_02817_ ), .A3(_02715_ ), .ZN(_02818_ ) );
MUX2_X1 _10448_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02819_ ) );
MUX2_X1 _10449_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02820_ ) );
MUX2_X1 _10450_ ( .A(_02819_ ), .B(_02820_ ), .S(_02641_ ), .Z(_02821_ ) );
OAI211_X1 _10451_ ( .A(_02498_ ), .B(_02818_ ), .C1(_02821_ ), .C2(_02462_ ), .ZN(_02822_ ) );
OR2_X1 _10452_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02823_ ) );
OAI211_X1 _10453_ ( .A(_02823_ ), .B(fanout_net_26 ), .C1(_02453_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02824_ ) );
OR2_X1 _10454_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02825_ ) );
OAI211_X1 _10455_ ( .A(_02825_ ), .B(_02641_ ), .C1(_02633_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02826_ ) );
NAND3_X1 _10456_ ( .A1(_02824_ ), .A2(_02826_ ), .A3(fanout_net_28 ), .ZN(_02827_ ) );
MUX2_X1 _10457_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02828_ ) );
MUX2_X1 _10458_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02829_ ) );
MUX2_X1 _10459_ ( .A(_02828_ ), .B(_02829_ ), .S(fanout_net_26 ), .Z(_02830_ ) );
OAI211_X1 _10460_ ( .A(fanout_net_30 ), .B(_02827_ ), .C1(_02830_ ), .C2(fanout_net_28 ), .ZN(_02831_ ) );
OAI211_X1 _10461_ ( .A(_02822_ ), .B(_02831_ ), .C1(_02629_ ), .C2(_02630_ ), .ZN(_02832_ ) );
NAND2_X4 _10462_ ( .A1(_02813_ ), .A2(_02832_ ), .ZN(_02833_ ) );
XNOR2_X2 _10463_ ( .A(_02833_ ), .B(\ID_EX_imm [5] ), .ZN(_02834_ ) );
OR2_X1 _10464_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02835_ ) );
OAI211_X1 _10465_ ( .A(_02835_ ), .B(_02446_ ), .C1(_02453_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02836_ ) );
OR2_X1 _10466_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02837_ ) );
OAI211_X1 _10467_ ( .A(_02837_ ), .B(fanout_net_26 ), .C1(_02453_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02838_ ) );
NAND3_X1 _10468_ ( .A1(_02836_ ), .A2(_02838_ ), .A3(fanout_net_28 ), .ZN(_02839_ ) );
MUX2_X1 _10469_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02840_ ) );
MUX2_X1 _10470_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02841_ ) );
MUX2_X1 _10471_ ( .A(_02840_ ), .B(_02841_ ), .S(_02641_ ), .Z(_02842_ ) );
OAI211_X1 _10472_ ( .A(_02498_ ), .B(_02839_ ), .C1(_02842_ ), .C2(fanout_net_28 ), .ZN(_02843_ ) );
MUX2_X1 _10473_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02844_ ) );
MUX2_X1 _10474_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02845_ ) );
MUX2_X1 _10475_ ( .A(_02844_ ), .B(_02845_ ), .S(fanout_net_29 ), .Z(_02846_ ) );
AND2_X1 _10476_ ( .A1(_02846_ ), .A2(fanout_net_26 ), .ZN(_02847_ ) );
MUX2_X1 _10477_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02848_ ) );
MUX2_X1 _10478_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02849_ ) );
MUX2_X1 _10479_ ( .A(_02848_ ), .B(_02849_ ), .S(fanout_net_29 ), .Z(_02850_ ) );
AND2_X1 _10480_ ( .A1(_02850_ ), .A2(_02446_ ), .ZN(_02851_ ) );
OAI21_X1 _10481_ ( .A(fanout_net_30 ), .B1(_02847_ ), .B2(_02851_ ), .ZN(_02852_ ) );
NAND3_X1 _10482_ ( .A1(_02442_ ), .A2(_02843_ ), .A3(_02852_ ), .ZN(_02853_ ) );
OR3_X1 _10483_ ( .A1(_02485_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02489_ ), .ZN(_02854_ ) );
NAND2_X1 _10484_ ( .A1(_02853_ ), .A2(_02854_ ), .ZN(_02855_ ) );
INV_X1 _10485_ ( .A(\ID_EX_imm [4] ), .ZN(_02856_ ) );
XNOR2_X1 _10486_ ( .A(_02855_ ), .B(_02856_ ), .ZN(_02857_ ) );
INV_X1 _10487_ ( .A(_02857_ ), .ZN(_02858_ ) );
NOR3_X4 _10488_ ( .A1(_02812_ ), .A2(_02834_ ), .A3(_02858_ ), .ZN(_02859_ ) );
INV_X1 _10489_ ( .A(_02855_ ), .ZN(_02860_ ) );
NOR3_X1 _10490_ ( .A1(_02834_ ), .A2(_02856_ ), .A3(_02860_ ), .ZN(_02861_ ) );
INV_X1 _10491_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02862_ ) );
AOI21_X1 _10492_ ( .A(_02861_ ), .B1(_02862_ ), .B2(_02833_ ), .ZN(_02863_ ) );
INV_X1 _10493_ ( .A(_02863_ ), .ZN(_02864_ ) );
NOR2_X1 _10494_ ( .A1(_02859_ ), .A2(_02864_ ), .ZN(_02865_ ) );
OR2_X1 _10495_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02866_ ) );
OAI211_X1 _10496_ ( .A(_02866_ ), .B(_02446_ ), .C1(_02453_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02867_ ) );
OR2_X1 _10497_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02868_ ) );
OAI211_X1 _10498_ ( .A(_02868_ ), .B(fanout_net_26 ), .C1(_02453_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02869_ ) );
NAND3_X1 _10499_ ( .A1(_02867_ ), .A2(_02869_ ), .A3(fanout_net_29 ), .ZN(_02870_ ) );
MUX2_X1 _10500_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02871_ ) );
MUX2_X1 _10501_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02872_ ) );
MUX2_X1 _10502_ ( .A(_02871_ ), .B(_02872_ ), .S(_02446_ ), .Z(_02873_ ) );
OAI211_X1 _10503_ ( .A(_02498_ ), .B(_02870_ ), .C1(_02873_ ), .C2(fanout_net_29 ), .ZN(_02874_ ) );
MUX2_X1 _10504_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02875_ ) );
MUX2_X1 _10505_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02876_ ) );
MUX2_X1 _10506_ ( .A(_02875_ ), .B(_02876_ ), .S(fanout_net_29 ), .Z(_02877_ ) );
AND2_X1 _10507_ ( .A1(_02877_ ), .A2(fanout_net_26 ), .ZN(_02878_ ) );
MUX2_X1 _10508_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02879_ ) );
MUX2_X1 _10509_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02880_ ) );
MUX2_X1 _10510_ ( .A(_02879_ ), .B(_02880_ ), .S(fanout_net_29 ), .Z(_02881_ ) );
AND2_X1 _10511_ ( .A1(_02881_ ), .A2(_02642_ ), .ZN(_02882_ ) );
OAI21_X1 _10512_ ( .A(fanout_net_30 ), .B1(_02878_ ), .B2(_02882_ ), .ZN(_02883_ ) );
NAND3_X1 _10513_ ( .A1(_02442_ ), .A2(_02874_ ), .A3(_02883_ ), .ZN(_02884_ ) );
OR3_X1 _10514_ ( .A1(_02485_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02489_ ), .ZN(_02885_ ) );
NAND2_X2 _10515_ ( .A1(_02884_ ), .A2(_02885_ ), .ZN(_02886_ ) );
XNOR2_X1 _10516_ ( .A(_02886_ ), .B(\ID_EX_imm [7] ), .ZN(_02887_ ) );
OR3_X1 _10517_ ( .A1(_02485_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02489_ ), .ZN(_02888_ ) );
OR2_X1 _10518_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02889_ ) );
OAI211_X1 _10519_ ( .A(_02889_ ), .B(_02446_ ), .C1(_02453_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02890_ ) );
OR2_X1 _10520_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02891_ ) );
OAI211_X1 _10521_ ( .A(_02891_ ), .B(fanout_net_26 ), .C1(_02453_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02892_ ) );
NAND3_X1 _10522_ ( .A1(_02890_ ), .A2(_02892_ ), .A3(_02715_ ), .ZN(_02893_ ) );
MUX2_X1 _10523_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02894_ ) );
MUX2_X1 _10524_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02895_ ) );
MUX2_X1 _10525_ ( .A(_02894_ ), .B(_02895_ ), .S(_02641_ ), .Z(_02896_ ) );
OAI211_X1 _10526_ ( .A(_02498_ ), .B(_02893_ ), .C1(_02896_ ), .C2(_02462_ ), .ZN(_02897_ ) );
OR2_X1 _10527_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02898_ ) );
OAI211_X1 _10528_ ( .A(_02898_ ), .B(fanout_net_26 ), .C1(_02453_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02899_ ) );
OR2_X1 _10529_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02900_ ) );
OAI211_X1 _10530_ ( .A(_02900_ ), .B(_02641_ ), .C1(_02633_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02901_ ) );
NAND3_X1 _10531_ ( .A1(_02899_ ), .A2(_02901_ ), .A3(fanout_net_29 ), .ZN(_02902_ ) );
MUX2_X1 _10532_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02903_ ) );
MUX2_X1 _10533_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02904_ ) );
MUX2_X1 _10534_ ( .A(_02903_ ), .B(_02904_ ), .S(fanout_net_26 ), .Z(_02905_ ) );
OAI211_X1 _10535_ ( .A(fanout_net_30 ), .B(_02902_ ), .C1(_02905_ ), .C2(fanout_net_29 ), .ZN(_02906_ ) );
OAI211_X1 _10536_ ( .A(_02897_ ), .B(_02906_ ), .C1(_02629_ ), .C2(_02630_ ), .ZN(_02907_ ) );
NAND2_X1 _10537_ ( .A1(_02888_ ), .A2(_02907_ ), .ZN(_02908_ ) );
XOR2_X1 _10538_ ( .A(_02908_ ), .B(\ID_EX_imm [6] ), .Z(_02909_ ) );
INV_X1 _10539_ ( .A(_02909_ ), .ZN(_02910_ ) );
NOR3_X2 _10540_ ( .A1(_02865_ ), .A2(_02887_ ), .A3(_02910_ ), .ZN(_02911_ ) );
INV_X1 _10541_ ( .A(_02886_ ), .ZN(_02912_ ) );
OR2_X1 _10542_ ( .A1(_02912_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02913_ ) );
AND2_X1 _10543_ ( .A1(_02908_ ), .A2(\ID_EX_imm [6] ), .ZN(_02914_ ) );
INV_X1 _10544_ ( .A(_02914_ ), .ZN(_02915_ ) );
OAI21_X1 _10545_ ( .A(_02913_ ), .B1(_02887_ ), .B2(_02915_ ), .ZN(_02916_ ) );
NOR2_X2 _10546_ ( .A1(_02911_ ), .A2(_02916_ ), .ZN(_02917_ ) );
OR3_X1 _10547_ ( .A1(_02485_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02489_ ), .ZN(_02918_ ) );
OR2_X1 _10548_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02919_ ) );
OAI211_X1 _10549_ ( .A(_02919_ ), .B(_02641_ ), .C1(_02633_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02920_ ) );
OR2_X1 _10550_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02921_ ) );
OAI211_X1 _10551_ ( .A(_02921_ ), .B(fanout_net_26 ), .C1(_02633_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02922_ ) );
NAND3_X1 _10552_ ( .A1(_02920_ ), .A2(_02922_ ), .A3(_02715_ ), .ZN(_02923_ ) );
MUX2_X1 _10553_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02924_ ) );
MUX2_X1 _10554_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02925_ ) );
MUX2_X1 _10555_ ( .A(_02924_ ), .B(_02925_ ), .S(_02711_ ), .Z(_02926_ ) );
OAI211_X1 _10556_ ( .A(_02498_ ), .B(_02923_ ), .C1(_02926_ ), .C2(_02462_ ), .ZN(_02927_ ) );
OR2_X1 _10557_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02928_ ) );
OAI211_X1 _10558_ ( .A(_02928_ ), .B(fanout_net_26 ), .C1(_02633_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02929_ ) );
OR2_X1 _10559_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02930_ ) );
OAI211_X1 _10560_ ( .A(_02930_ ), .B(_02641_ ), .C1(_02633_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02931_ ) );
NAND3_X1 _10561_ ( .A1(_02929_ ), .A2(_02931_ ), .A3(fanout_net_29 ), .ZN(_02932_ ) );
MUX2_X1 _10562_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02933_ ) );
MUX2_X1 _10563_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02934_ ) );
MUX2_X1 _10564_ ( .A(_02933_ ), .B(_02934_ ), .S(fanout_net_26 ), .Z(_02935_ ) );
OAI211_X1 _10565_ ( .A(fanout_net_30 ), .B(_02932_ ), .C1(_02935_ ), .C2(fanout_net_29 ), .ZN(_02936_ ) );
OAI211_X1 _10566_ ( .A(_02927_ ), .B(_02936_ ), .C1(_02629_ ), .C2(_02630_ ), .ZN(_02937_ ) );
NAND2_X1 _10567_ ( .A1(_02918_ ), .A2(_02937_ ), .ZN(_02938_ ) );
INV_X1 _10568_ ( .A(\ID_EX_imm [8] ), .ZN(_02939_ ) );
XNOR2_X1 _10569_ ( .A(_02938_ ), .B(_02939_ ), .ZN(_02940_ ) );
OR3_X1 _10570_ ( .A1(_02434_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02440_ ), .ZN(_02941_ ) );
OR2_X1 _10571_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02942_ ) );
OAI211_X1 _10572_ ( .A(_02942_ ), .B(_02445_ ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02943_ ) );
OR2_X1 _10573_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02944_ ) );
OAI211_X1 _10574_ ( .A(_02944_ ), .B(fanout_net_26 ), .C1(_02661_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02945_ ) );
NAND3_X1 _10575_ ( .A1(_02943_ ), .A2(_02945_ ), .A3(_02461_ ), .ZN(_02946_ ) );
MUX2_X1 _10576_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02947_ ) );
MUX2_X1 _10577_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02948_ ) );
MUX2_X1 _10578_ ( .A(_02947_ ), .B(_02948_ ), .S(_02445_ ), .Z(_02949_ ) );
OAI211_X1 _10579_ ( .A(fanout_net_30 ), .B(_02946_ ), .C1(_02949_ ), .C2(_02461_ ), .ZN(_02950_ ) );
OR2_X1 _10580_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02951_ ) );
OAI211_X1 _10581_ ( .A(_02951_ ), .B(_02445_ ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02952_ ) );
OR2_X1 _10582_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02953_ ) );
OAI211_X1 _10583_ ( .A(_02953_ ), .B(fanout_net_26 ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02954_ ) );
NAND3_X1 _10584_ ( .A1(_02952_ ), .A2(_02954_ ), .A3(_02461_ ), .ZN(_02955_ ) );
OR2_X1 _10585_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02956_ ) );
OAI211_X1 _10586_ ( .A(_02956_ ), .B(_02445_ ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02957_ ) );
OR2_X1 _10587_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02958_ ) );
OAI211_X1 _10588_ ( .A(_02958_ ), .B(fanout_net_26 ), .C1(_02452_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02959_ ) );
NAND3_X1 _10589_ ( .A1(_02957_ ), .A2(_02959_ ), .A3(fanout_net_29 ), .ZN(_02960_ ) );
NAND3_X1 _10590_ ( .A1(_02955_ ), .A2(_02960_ ), .A3(_02497_ ), .ZN(_02961_ ) );
OAI211_X1 _10591_ ( .A(_02950_ ), .B(_02961_ ), .C1(_02434_ ), .C2(_02440_ ), .ZN(_02962_ ) );
NAND2_X4 _10592_ ( .A1(_02941_ ), .A2(_02962_ ), .ZN(_02963_ ) );
INV_X1 _10593_ ( .A(\ID_EX_imm [9] ), .ZN(_02964_ ) );
XNOR2_X1 _10594_ ( .A(_02963_ ), .B(_02964_ ), .ZN(_02965_ ) );
NAND2_X1 _10595_ ( .A1(_02940_ ), .A2(_02965_ ), .ZN(_02966_ ) );
OR3_X1 _10596_ ( .A1(_02485_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_02489_ ), .ZN(_02967_ ) );
INV_X1 _10597_ ( .A(\ID_EX_imm [11] ), .ZN(_02968_ ) );
OR2_X1 _10598_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02969_ ) );
OAI211_X1 _10599_ ( .A(_02969_ ), .B(_02641_ ), .C1(_02633_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02970_ ) );
OR2_X1 _10600_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02971_ ) );
OAI211_X1 _10601_ ( .A(_02971_ ), .B(fanout_net_26 ), .C1(_02662_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02972_ ) );
NAND3_X1 _10602_ ( .A1(_02970_ ), .A2(_02972_ ), .A3(_02715_ ), .ZN(_02973_ ) );
MUX2_X1 _10603_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02974_ ) );
MUX2_X1 _10604_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02975_ ) );
MUX2_X1 _10605_ ( .A(_02974_ ), .B(_02975_ ), .S(_02711_ ), .Z(_02976_ ) );
OAI211_X1 _10606_ ( .A(_02498_ ), .B(_02973_ ), .C1(_02976_ ), .C2(_02462_ ), .ZN(_02977_ ) );
OR2_X1 _10607_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02978_ ) );
OAI211_X1 _10608_ ( .A(_02978_ ), .B(fanout_net_26 ), .C1(_02633_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02979_ ) );
OR2_X1 _10609_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02980_ ) );
OAI211_X1 _10610_ ( .A(_02980_ ), .B(_02641_ ), .C1(_02662_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02981_ ) );
NAND3_X1 _10611_ ( .A1(_02979_ ), .A2(_02981_ ), .A3(fanout_net_29 ), .ZN(_02982_ ) );
MUX2_X1 _10612_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02983_ ) );
MUX2_X1 _10613_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02984_ ) );
MUX2_X1 _10614_ ( .A(_02983_ ), .B(_02984_ ), .S(fanout_net_26 ), .Z(_02985_ ) );
OAI211_X1 _10615_ ( .A(fanout_net_30 ), .B(_02982_ ), .C1(_02985_ ), .C2(fanout_net_29 ), .ZN(_02986_ ) );
OAI211_X1 _10616_ ( .A(_02977_ ), .B(_02986_ ), .C1(_02629_ ), .C2(_02630_ ), .ZN(_02987_ ) );
AND3_X1 _10617_ ( .A1(_02967_ ), .A2(_02968_ ), .A3(_02987_ ), .ZN(_02988_ ) );
AOI21_X1 _10618_ ( .A(_02968_ ), .B1(_02967_ ), .B2(_02987_ ), .ZN(_02989_ ) );
NOR2_X1 _10619_ ( .A1(_02988_ ), .A2(_02989_ ), .ZN(_02990_ ) );
INV_X1 _10620_ ( .A(_02990_ ), .ZN(_02991_ ) );
OR3_X1 _10621_ ( .A1(_02629_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02630_ ), .ZN(_02992_ ) );
OR2_X1 _10622_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02993_ ) );
OAI211_X1 _10623_ ( .A(_02993_ ), .B(_02642_ ), .C1(_02663_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02994_ ) );
OR2_X1 _10624_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02995_ ) );
OAI211_X1 _10625_ ( .A(_02995_ ), .B(fanout_net_26 ), .C1(_02663_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02996_ ) );
NAND3_X1 _10626_ ( .A1(_02994_ ), .A2(_02996_ ), .A3(_02462_ ), .ZN(_02997_ ) );
MUX2_X1 _10627_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02998_ ) );
MUX2_X1 _10628_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02999_ ) );
MUX2_X1 _10629_ ( .A(_02998_ ), .B(_02999_ ), .S(_02446_ ), .Z(_03000_ ) );
OAI211_X1 _10630_ ( .A(_02498_ ), .B(_02997_ ), .C1(_03000_ ), .C2(_02463_ ), .ZN(_03001_ ) );
OR2_X1 _10631_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03002_ ) );
OAI211_X1 _10632_ ( .A(_03002_ ), .B(fanout_net_26 ), .C1(_02663_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03003_ ) );
OR2_X1 _10633_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03004_ ) );
OAI211_X1 _10634_ ( .A(_03004_ ), .B(_02642_ ), .C1(_02663_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03005_ ) );
NAND3_X1 _10635_ ( .A1(_03003_ ), .A2(_03005_ ), .A3(fanout_net_29 ), .ZN(_03006_ ) );
MUX2_X1 _10636_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03007_ ) );
MUX2_X1 _10637_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03008_ ) );
MUX2_X1 _10638_ ( .A(_03007_ ), .B(_03008_ ), .S(fanout_net_26 ), .Z(_03009_ ) );
OAI211_X1 _10639_ ( .A(fanout_net_30 ), .B(_03006_ ), .C1(_03009_ ), .C2(fanout_net_29 ), .ZN(_03010_ ) );
OAI211_X1 _10640_ ( .A(_03001_ ), .B(_03010_ ), .C1(_02629_ ), .C2(_02490_ ), .ZN(_03011_ ) );
NAND2_X2 _10641_ ( .A1(_02992_ ), .A2(_03011_ ), .ZN(_03012_ ) );
XNOR2_X1 _10642_ ( .A(_03012_ ), .B(\ID_EX_imm [10] ), .ZN(_03013_ ) );
NOR3_X1 _10643_ ( .A1(_02966_ ), .A2(_02991_ ), .A3(_03013_ ), .ZN(_03014_ ) );
INV_X1 _10644_ ( .A(_03014_ ), .ZN(_03015_ ) );
NOR2_X2 _10645_ ( .A1(_02917_ ), .A2(_03015_ ), .ZN(_03016_ ) );
AND2_X1 _10646_ ( .A1(_02938_ ), .A2(\ID_EX_imm [8] ), .ZN(_03017_ ) );
AND2_X1 _10647_ ( .A1(_02965_ ), .A2(_03017_ ), .ZN(_03018_ ) );
AOI21_X1 _10648_ ( .A(_03018_ ), .B1(\ID_EX_imm [9] ), .B2(_02963_ ), .ZN(_03019_ ) );
OR3_X1 _10649_ ( .A1(_03019_ ), .A2(_02991_ ), .A3(_03013_ ), .ZN(_03020_ ) );
AND2_X1 _10650_ ( .A1(_03012_ ), .A2(\ID_EX_imm [10] ), .ZN(_03021_ ) );
AOI21_X1 _10651_ ( .A(_02989_ ), .B1(_02990_ ), .B2(_03021_ ), .ZN(_03022_ ) );
AND2_X1 _10652_ ( .A1(_03020_ ), .A2(_03022_ ), .ZN(_03023_ ) );
INV_X1 _10653_ ( .A(_03023_ ), .ZN(_03024_ ) );
NOR2_X2 _10654_ ( .A1(_03016_ ), .A2(_03024_ ), .ZN(_03025_ ) );
OR2_X1 _10655_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03026_ ) );
OAI211_X1 _10656_ ( .A(_03026_ ), .B(_02642_ ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03027_ ) );
OR2_X1 _10657_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03028_ ) );
OAI211_X1 _10658_ ( .A(_03028_ ), .B(fanout_net_26 ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03029_ ) );
NAND3_X1 _10659_ ( .A1(_03027_ ), .A2(_03029_ ), .A3(fanout_net_29 ), .ZN(_03030_ ) );
MUX2_X1 _10660_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03031_ ) );
MUX2_X1 _10661_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03032_ ) );
MUX2_X1 _10662_ ( .A(_03031_ ), .B(_03032_ ), .S(_02642_ ), .Z(_03033_ ) );
OAI211_X1 _10663_ ( .A(_02499_ ), .B(_03030_ ), .C1(_03033_ ), .C2(fanout_net_29 ), .ZN(_03034_ ) );
MUX2_X1 _10664_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03035_ ) );
MUX2_X1 _10665_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03036_ ) );
MUX2_X1 _10666_ ( .A(_03035_ ), .B(_03036_ ), .S(fanout_net_29 ), .Z(_03037_ ) );
AND2_X1 _10667_ ( .A1(_03037_ ), .A2(fanout_net_26 ), .ZN(_03038_ ) );
MUX2_X1 _10668_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03039_ ) );
MUX2_X1 _10669_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_03040_ ) );
MUX2_X1 _10670_ ( .A(_03039_ ), .B(_03040_ ), .S(fanout_net_29 ), .Z(_03041_ ) );
AND2_X1 _10671_ ( .A1(_03041_ ), .A2(_02447_ ), .ZN(_03042_ ) );
OAI21_X1 _10672_ ( .A(fanout_net_30 ), .B1(_03038_ ), .B2(_03042_ ), .ZN(_03043_ ) );
NAND3_X1 _10673_ ( .A1(_02442_ ), .A2(_03034_ ), .A3(_03043_ ), .ZN(_03044_ ) );
INV_X1 _10674_ ( .A(\ID_EX_imm [13] ), .ZN(_03045_ ) );
OR3_X2 _10675_ ( .A1(_02629_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02630_ ), .ZN(_03046_ ) );
AND3_X1 _10676_ ( .A1(_03044_ ), .A2(_03045_ ), .A3(_03046_ ), .ZN(_03047_ ) );
AOI21_X1 _10677_ ( .A(_03045_ ), .B1(_03044_ ), .B2(_03046_ ), .ZN(_03048_ ) );
NOR2_X1 _10678_ ( .A1(_03047_ ), .A2(_03048_ ), .ZN(_03049_ ) );
OR3_X1 _10679_ ( .A1(_02629_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02630_ ), .ZN(_03050_ ) );
OR2_X1 _10680_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03051_ ) );
OAI211_X1 _10681_ ( .A(_03051_ ), .B(_02642_ ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03052_ ) );
OR2_X1 _10682_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03053_ ) );
OAI211_X1 _10683_ ( .A(_03053_ ), .B(fanout_net_27 ), .C1(_02663_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03054_ ) );
NAND3_X1 _10684_ ( .A1(_03052_ ), .A2(_03054_ ), .A3(_02462_ ), .ZN(_03055_ ) );
MUX2_X1 _10685_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03056_ ) );
MUX2_X1 _10686_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03057_ ) );
MUX2_X1 _10687_ ( .A(_03056_ ), .B(_03057_ ), .S(_02642_ ), .Z(_03058_ ) );
OAI211_X1 _10688_ ( .A(_02499_ ), .B(_03055_ ), .C1(_03058_ ), .C2(_02463_ ), .ZN(_03059_ ) );
OR2_X1 _10689_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03060_ ) );
OAI211_X1 _10690_ ( .A(_03060_ ), .B(fanout_net_27 ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03061_ ) );
OR2_X1 _10691_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03062_ ) );
OAI211_X1 _10692_ ( .A(_03062_ ), .B(_02642_ ), .C1(_02663_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03063_ ) );
NAND3_X1 _10693_ ( .A1(_03061_ ), .A2(_03063_ ), .A3(fanout_net_29 ), .ZN(_03064_ ) );
MUX2_X1 _10694_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03065_ ) );
MUX2_X1 _10695_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03066_ ) );
MUX2_X1 _10696_ ( .A(_03065_ ), .B(_03066_ ), .S(fanout_net_27 ), .Z(_03067_ ) );
OAI211_X1 _10697_ ( .A(fanout_net_30 ), .B(_03064_ ), .C1(_03067_ ), .C2(fanout_net_29 ), .ZN(_03068_ ) );
OAI211_X1 _10698_ ( .A(_03059_ ), .B(_03068_ ), .C1(_02486_ ), .C2(_02490_ ), .ZN(_03069_ ) );
NAND2_X1 _10699_ ( .A1(_03050_ ), .A2(_03069_ ), .ZN(_03070_ ) );
INV_X1 _10700_ ( .A(\ID_EX_imm [12] ), .ZN(_03071_ ) );
XNOR2_X1 _10701_ ( .A(_03070_ ), .B(_03071_ ), .ZN(_03072_ ) );
AND2_X1 _10702_ ( .A1(_03049_ ), .A2(_03072_ ), .ZN(_03073_ ) );
OR3_X1 _10703_ ( .A1(_02485_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02489_ ), .ZN(_03074_ ) );
OR2_X1 _10704_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03075_ ) );
OAI211_X1 _10705_ ( .A(_03075_ ), .B(_02711_ ), .C1(_02662_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03076_ ) );
OR2_X1 _10706_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03077_ ) );
OAI211_X1 _10707_ ( .A(_03077_ ), .B(fanout_net_27 ), .C1(_02662_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03078_ ) );
NAND3_X1 _10708_ ( .A1(_03076_ ), .A2(_03078_ ), .A3(_02715_ ), .ZN(_03079_ ) );
MUX2_X1 _10709_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03080_ ) );
MUX2_X1 _10710_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03081_ ) );
MUX2_X1 _10711_ ( .A(_03080_ ), .B(_03081_ ), .S(_02711_ ), .Z(_03082_ ) );
OAI211_X1 _10712_ ( .A(_02498_ ), .B(_03079_ ), .C1(_03082_ ), .C2(_02715_ ), .ZN(_03083_ ) );
OR2_X1 _10713_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03084_ ) );
OAI211_X1 _10714_ ( .A(_03084_ ), .B(fanout_net_27 ), .C1(_02662_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03085_ ) );
OR2_X1 _10715_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03086_ ) );
OAI211_X1 _10716_ ( .A(_03086_ ), .B(_02711_ ), .C1(_02662_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03087_ ) );
NAND3_X1 _10717_ ( .A1(_03085_ ), .A2(_03087_ ), .A3(fanout_net_29 ), .ZN(_03088_ ) );
MUX2_X1 _10718_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03089_ ) );
MUX2_X1 _10719_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03090_ ) );
MUX2_X1 _10720_ ( .A(_03089_ ), .B(_03090_ ), .S(fanout_net_27 ), .Z(_03091_ ) );
OAI211_X1 _10721_ ( .A(fanout_net_30 ), .B(_03088_ ), .C1(_03091_ ), .C2(fanout_net_29 ), .ZN(_03092_ ) );
OAI211_X1 _10722_ ( .A(_03083_ ), .B(_03092_ ), .C1(_02485_ ), .C2(_02489_ ), .ZN(_03093_ ) );
NAND2_X2 _10723_ ( .A1(_03074_ ), .A2(_03093_ ), .ZN(_03094_ ) );
XOR2_X1 _10724_ ( .A(_03094_ ), .B(\ID_EX_imm [15] ), .Z(_03095_ ) );
OR3_X1 _10725_ ( .A1(_02486_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02630_ ), .ZN(_03096_ ) );
OR2_X1 _10726_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03097_ ) );
OAI211_X1 _10727_ ( .A(_03097_ ), .B(_02447_ ), .C1(_02454_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03098_ ) );
OR2_X1 _10728_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03099_ ) );
OAI211_X1 _10729_ ( .A(_03099_ ), .B(fanout_net_27 ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03100_ ) );
NAND3_X1 _10730_ ( .A1(_03098_ ), .A2(_03100_ ), .A3(_02463_ ), .ZN(_03101_ ) );
MUX2_X1 _10731_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03102_ ) );
MUX2_X1 _10732_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03103_ ) );
MUX2_X1 _10733_ ( .A(_03102_ ), .B(_03103_ ), .S(_02447_ ), .Z(_03104_ ) );
OAI211_X1 _10734_ ( .A(fanout_net_30 ), .B(_03101_ ), .C1(_03104_ ), .C2(_02463_ ), .ZN(_03105_ ) );
OR2_X1 _10735_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03106_ ) );
OAI211_X1 _10736_ ( .A(_03106_ ), .B(_02447_ ), .C1(_02454_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03107_ ) );
OR2_X1 _10737_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03108_ ) );
OAI211_X1 _10738_ ( .A(_03108_ ), .B(fanout_net_27 ), .C1(_02454_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03109_ ) );
AOI21_X1 _10739_ ( .A(_02462_ ), .B1(_03107_ ), .B2(_03109_ ), .ZN(_03110_ ) );
OR2_X1 _10740_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03111_ ) );
OAI211_X1 _10741_ ( .A(_03111_ ), .B(_02447_ ), .C1(_02454_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03112_ ) );
OR2_X1 _10742_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03113_ ) );
OAI211_X1 _10743_ ( .A(_03113_ ), .B(fanout_net_27 ), .C1(_02634_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03114_ ) );
AOI21_X1 _10744_ ( .A(fanout_net_29 ), .B1(_03112_ ), .B2(_03114_ ), .ZN(_03115_ ) );
OAI21_X1 _10745_ ( .A(_02499_ ), .B1(_03110_ ), .B2(_03115_ ), .ZN(_03116_ ) );
OAI211_X1 _10746_ ( .A(_03105_ ), .B(_03116_ ), .C1(_02486_ ), .C2(_02490_ ), .ZN(_03117_ ) );
NAND2_X2 _10747_ ( .A1(_03096_ ), .A2(_03117_ ), .ZN(_03118_ ) );
INV_X1 _10748_ ( .A(\ID_EX_imm [14] ), .ZN(_03119_ ) );
XNOR2_X1 _10749_ ( .A(_03118_ ), .B(_03119_ ), .ZN(_03120_ ) );
NAND3_X1 _10750_ ( .A1(_03073_ ), .A2(_03095_ ), .A3(_03120_ ), .ZN(_03121_ ) );
OR2_X2 _10751_ ( .A1(_03025_ ), .A2(_03121_ ), .ZN(_03122_ ) );
NAND2_X1 _10752_ ( .A1(_03070_ ), .A2(\ID_EX_imm [12] ), .ZN(_03123_ ) );
NOR3_X1 _10753_ ( .A1(_03047_ ), .A2(_03048_ ), .A3(_03123_ ), .ZN(_03124_ ) );
OAI211_X1 _10754_ ( .A(_03095_ ), .B(_03120_ ), .C1(_03124_ ), .C2(_03048_ ), .ZN(_03125_ ) );
NAND2_X1 _10755_ ( .A1(_03094_ ), .A2(\ID_EX_imm [15] ), .ZN(_03126_ ) );
NAND3_X1 _10756_ ( .A1(_03095_ ), .A2(\ID_EX_imm [14] ), .A3(_03118_ ), .ZN(_03127_ ) );
AND3_X1 _10757_ ( .A1(_03125_ ), .A2(_03126_ ), .A3(_03127_ ), .ZN(_03128_ ) );
AOI211_X1 _10758_ ( .A(_02603_ ), .B(_02709_ ), .C1(_03122_ ), .C2(_03128_ ), .ZN(_03129_ ) );
AND2_X1 _10759_ ( .A1(_02706_ ), .A2(\ID_EX_imm [16] ), .ZN(_03130_ ) );
AND2_X1 _10760_ ( .A1(_02684_ ), .A2(_03130_ ), .ZN(_03131_ ) );
AOI21_X1 _10761_ ( .A(_03131_ ), .B1(\ID_EX_imm [17] ), .B2(_02682_ ), .ZN(_03132_ ) );
INV_X1 _10762_ ( .A(_03132_ ), .ZN(_03133_ ) );
NAND2_X1 _10763_ ( .A1(_03133_ ), .A2(_02658_ ), .ZN(_03134_ ) );
AND2_X1 _10764_ ( .A1(_02626_ ), .A2(\ID_EX_imm [18] ), .ZN(_03135_ ) );
AND2_X1 _10765_ ( .A1(_02657_ ), .A2(_03135_ ), .ZN(_03136_ ) );
AOI21_X1 _10766_ ( .A(_03136_ ), .B1(\ID_EX_imm [19] ), .B2(_02655_ ), .ZN(_03137_ ) );
AND2_X1 _10767_ ( .A1(_03134_ ), .A2(_03137_ ), .ZN(_03138_ ) );
OR2_X1 _10768_ ( .A1(_03138_ ), .A2(_02603_ ), .ZN(_03139_ ) );
AND2_X1 _10769_ ( .A1(_02598_ ), .A2(\ID_EX_imm [20] ), .ZN(_03140_ ) );
AND2_X1 _10770_ ( .A1(_02577_ ), .A2(_03140_ ), .ZN(_03141_ ) );
AOI21_X1 _10771_ ( .A(_03141_ ), .B1(\ID_EX_imm [21] ), .B2(_02575_ ), .ZN(_03142_ ) );
INV_X1 _10772_ ( .A(_03142_ ), .ZN(_03143_ ) );
NAND2_X1 _10773_ ( .A1(_03143_ ), .A2(_02550_ ), .ZN(_03144_ ) );
NAND4_X1 _10774_ ( .A1(_02549_ ), .A2(\ID_EX_imm [22] ), .A3(_02546_ ), .A4(_02522_ ), .ZN(_03145_ ) );
NAND4_X1 _10775_ ( .A1(_03139_ ), .A2(_02549_ ), .A3(_03144_ ), .A4(_03145_ ), .ZN(_03146_ ) );
OR2_X1 _10776_ ( .A1(_03129_ ), .A2(_03146_ ), .ZN(_03147_ ) );
OR3_X1 _10777_ ( .A1(_02488_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02492_ ), .ZN(_03148_ ) );
OR2_X1 _10778_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03149_ ) );
OAI211_X1 _10779_ ( .A(_03149_ ), .B(_02450_ ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03150_ ) );
OR2_X1 _10780_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03151_ ) );
OAI211_X1 _10781_ ( .A(_03151_ ), .B(fanout_net_27 ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03152_ ) );
NAND3_X1 _10782_ ( .A1(_03150_ ), .A2(_03152_ ), .A3(fanout_net_29 ), .ZN(_03153_ ) );
MUX2_X1 _10783_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03154_ ) );
MUX2_X1 _10784_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_03155_ ) );
MUX2_X1 _10785_ ( .A(_03154_ ), .B(_03155_ ), .S(_02470_ ), .Z(_03156_ ) );
OAI211_X1 _10786_ ( .A(_02686_ ), .B(_03153_ ), .C1(_03156_ ), .C2(fanout_net_29 ), .ZN(_03157_ ) );
NOR2_X1 _10787_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03158_ ) );
BUF_X2 _10788_ ( .A(_02501_ ), .Z(_03159_ ) );
OAI21_X1 _10789_ ( .A(_02470_ ), .B1(_03159_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03160_ ) );
INV_X1 _10790_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03161_ ) );
INV_X1 _10791_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03162_ ) );
MUX2_X1 _10792_ ( .A(_03161_ ), .B(_03162_ ), .S(fanout_net_23 ), .Z(_03163_ ) );
OAI221_X1 _10793_ ( .A(_02465_ ), .B1(_03158_ ), .B2(_03160_ ), .C1(_03163_ ), .C2(_02450_ ), .ZN(_03164_ ) );
NOR2_X1 _10794_ ( .A1(_03159_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03165_ ) );
OAI21_X1 _10795_ ( .A(fanout_net_27 ), .B1(fanout_net_23 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03166_ ) );
NOR2_X1 _10796_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03167_ ) );
OAI21_X1 _10797_ ( .A(_02450_ ), .B1(_02456_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03168_ ) );
OAI221_X1 _10798_ ( .A(fanout_net_29 ), .B1(_03165_ ), .B2(_03166_ ), .C1(_03167_ ), .C2(_03168_ ), .ZN(_03169_ ) );
NAND3_X1 _10799_ ( .A1(_03164_ ), .A2(_03169_ ), .A3(fanout_net_30 ), .ZN(_03170_ ) );
OAI211_X1 _10800_ ( .A(_03157_ ), .B(_03170_ ), .C1(_02488_ ), .C2(_02492_ ), .ZN(_03171_ ) );
NAND2_X1 _10801_ ( .A1(_03148_ ), .A2(_03171_ ), .ZN(_03172_ ) );
INV_X1 _10802_ ( .A(\ID_EX_imm [24] ), .ZN(_03173_ ) );
XNOR2_X1 _10803_ ( .A(_03172_ ), .B(_03173_ ), .ZN(_03174_ ) );
AND2_X1 _10804_ ( .A1(_03147_ ), .A2(_03174_ ), .ZN(_03175_ ) );
AOI21_X1 _10805_ ( .A(_03173_ ), .B1(_03148_ ), .B2(_03171_ ), .ZN(_03176_ ) );
NOR2_X2 _10806_ ( .A1(_03175_ ), .A2(_03176_ ), .ZN(_03177_ ) );
OR3_X1 _10807_ ( .A1(_02487_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02491_ ), .ZN(_03178_ ) );
OR2_X1 _10808_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03179_ ) );
OAI211_X1 _10809_ ( .A(_03179_ ), .B(_02470_ ), .C1(_03159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03180_ ) );
OR2_X1 _10810_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03181_ ) );
OAI211_X1 _10811_ ( .A(_03181_ ), .B(fanout_net_27 ), .C1(_02455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03182_ ) );
NAND3_X1 _10812_ ( .A1(_03180_ ), .A2(_03182_ ), .A3(_02465_ ), .ZN(_03183_ ) );
MUX2_X1 _10813_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03184_ ) );
MUX2_X1 _10814_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03185_ ) );
MUX2_X1 _10815_ ( .A(_03184_ ), .B(_03185_ ), .S(_02449_ ), .Z(_03186_ ) );
OAI211_X1 _10816_ ( .A(_02686_ ), .B(_03183_ ), .C1(_03186_ ), .C2(_02465_ ), .ZN(_03187_ ) );
OR2_X1 _10817_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03188_ ) );
OAI211_X1 _10818_ ( .A(_03188_ ), .B(fanout_net_27 ), .C1(_03159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03189_ ) );
OR2_X1 _10819_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03190_ ) );
OAI211_X1 _10820_ ( .A(_03190_ ), .B(_02449_ ), .C1(_02455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03191_ ) );
NAND3_X1 _10821_ ( .A1(_03189_ ), .A2(_03191_ ), .A3(fanout_net_29 ), .ZN(_03192_ ) );
MUX2_X1 _10822_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03193_ ) );
MUX2_X1 _10823_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03194_ ) );
MUX2_X1 _10824_ ( .A(_03193_ ), .B(_03194_ ), .S(fanout_net_27 ), .Z(_03195_ ) );
OAI211_X1 _10825_ ( .A(fanout_net_30 ), .B(_03192_ ), .C1(_03195_ ), .C2(fanout_net_29 ), .ZN(_03196_ ) );
OAI211_X1 _10826_ ( .A(_03187_ ), .B(_03196_ ), .C1(_02488_ ), .C2(_02492_ ), .ZN(_03197_ ) );
NAND2_X1 _10827_ ( .A1(_03178_ ), .A2(_03197_ ), .ZN(_03198_ ) );
NAND2_X1 _10828_ ( .A1(_03198_ ), .A2(\ID_EX_imm [25] ), .ZN(_03199_ ) );
NAND2_X2 _10829_ ( .A1(_03177_ ), .A2(_03199_ ), .ZN(_03200_ ) );
OR3_X1 _10830_ ( .A1(_02488_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02492_ ), .ZN(_03201_ ) );
OR2_X1 _10831_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03202_ ) );
OAI211_X1 _10832_ ( .A(_03202_ ), .B(_02470_ ), .C1(_03159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03203_ ) );
OR2_X1 _10833_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03204_ ) );
OAI211_X1 _10834_ ( .A(_03204_ ), .B(fanout_net_27 ), .C1(_03159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03205_ ) );
NAND3_X1 _10835_ ( .A1(_03203_ ), .A2(_03205_ ), .A3(_02465_ ), .ZN(_03206_ ) );
MUX2_X1 _10836_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03207_ ) );
MUX2_X1 _10837_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03208_ ) );
MUX2_X1 _10838_ ( .A(_03207_ ), .B(_03208_ ), .S(_02470_ ), .Z(_03209_ ) );
OAI211_X1 _10839_ ( .A(_02686_ ), .B(_03206_ ), .C1(_03209_ ), .C2(_02465_ ), .ZN(_03210_ ) );
OR2_X1 _10840_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03211_ ) );
OAI211_X1 _10841_ ( .A(_03211_ ), .B(_02449_ ), .C1(_03159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03212_ ) );
NOR2_X1 _10842_ ( .A1(_03159_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03213_ ) );
OAI21_X1 _10843_ ( .A(fanout_net_27 ), .B1(fanout_net_24 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03214_ ) );
OAI211_X1 _10844_ ( .A(_03212_ ), .B(fanout_net_29 ), .C1(_03213_ ), .C2(_03214_ ), .ZN(_03215_ ) );
MUX2_X1 _10845_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03216_ ) );
MUX2_X1 _10846_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03217_ ) );
MUX2_X1 _10847_ ( .A(_03216_ ), .B(_03217_ ), .S(fanout_net_27 ), .Z(_03218_ ) );
OAI211_X1 _10848_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03215_ ), .C1(_03218_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03219_ ) );
OAI211_X1 _10849_ ( .A(_03210_ ), .B(_03219_ ), .C1(_02488_ ), .C2(_02492_ ), .ZN(_03220_ ) );
NAND2_X1 _10850_ ( .A1(_03201_ ), .A2(_03220_ ), .ZN(_03221_ ) );
XNOR2_X1 _10851_ ( .A(_03221_ ), .B(\ID_EX_imm [26] ), .ZN(_03222_ ) );
INV_X1 _10852_ ( .A(_03222_ ), .ZN(_03223_ ) );
INV_X1 _10853_ ( .A(\ID_EX_imm [25] ), .ZN(_03224_ ) );
NAND3_X1 _10854_ ( .A1(_03178_ ), .A2(_03224_ ), .A3(_03197_ ), .ZN(_03225_ ) );
AND4_X2 _10855_ ( .A1(_02496_ ), .A2(_03200_ ), .A3(_03223_ ), .A4(_03225_ ), .ZN(_03226_ ) );
INV_X1 _10856_ ( .A(_03221_ ), .ZN(_03227_ ) );
OR2_X1 _10857_ ( .A1(_03227_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03228_ ) );
NOR3_X1 _10858_ ( .A1(_03228_ ), .A2(_02494_ ), .A3(_02495_ ), .ZN(_03229_ ) );
OR2_X1 _10859_ ( .A1(_03229_ ), .A2(_02495_ ), .ZN(_03230_ ) );
NOR2_X2 _10860_ ( .A1(_03226_ ), .A2(_03230_ ), .ZN(_03231_ ) );
OR2_X1 _10861_ ( .A1(_02455_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03232_ ) );
OAI211_X1 _10862_ ( .A(_03232_ ), .B(_02450_ ), .C1(fanout_net_24 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03233_ ) );
OR2_X1 _10863_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03234_ ) );
OAI211_X1 _10864_ ( .A(_03234_ ), .B(fanout_net_27 ), .C1(_02456_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03235_ ) );
NAND3_X1 _10865_ ( .A1(_03233_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03235_ ), .ZN(_03236_ ) );
MUX2_X1 _10866_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03237_ ) );
MUX2_X1 _10867_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03238_ ) );
MUX2_X1 _10868_ ( .A(_03237_ ), .B(_03238_ ), .S(_02470_ ), .Z(_03239_ ) );
OAI211_X1 _10869_ ( .A(_02686_ ), .B(_03236_ ), .C1(_03239_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03240_ ) );
MUX2_X1 _10870_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03241_ ) );
AND2_X1 _10871_ ( .A1(_03241_ ), .A2(fanout_net_27 ), .ZN(_03242_ ) );
MUX2_X1 _10872_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03243_ ) );
AOI211_X1 _10873_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_03242_ ), .C1(_02450_ ), .C2(_03243_ ), .ZN(_03244_ ) );
INV_X1 _10874_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03245_ ) );
AOI21_X1 _10875_ ( .A(fanout_net_27 ), .B1(_03245_ ), .B2(fanout_net_24 ), .ZN(_03246_ ) );
OR2_X1 _10876_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03247_ ) );
MUX2_X1 _10877_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03248_ ) );
AOI221_X4 _10878_ ( .A(_02464_ ), .B1(_03246_ ), .B2(_03247_ ), .C1(_03248_ ), .C2(fanout_net_27 ), .ZN(_03249_ ) );
OR3_X1 _10879_ ( .A1(_03244_ ), .A2(_03249_ ), .A3(_02686_ ), .ZN(_03250_ ) );
NAND3_X1 _10880_ ( .A1(_02442_ ), .A2(_03240_ ), .A3(_03250_ ), .ZN(_03251_ ) );
OR3_X1 _10881_ ( .A1(_02488_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02492_ ), .ZN(_03252_ ) );
NAND2_X1 _10882_ ( .A1(_03251_ ), .A2(_03252_ ), .ZN(_03253_ ) );
XNOR2_X1 _10883_ ( .A(_03253_ ), .B(\ID_EX_imm [28] ), .ZN(_03254_ ) );
NOR2_X1 _10884_ ( .A1(_03231_ ), .A2(_03254_ ), .ZN(_03255_ ) );
OR3_X1 _10885_ ( .A1(_02487_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02491_ ), .ZN(_03256_ ) );
OR2_X1 _10886_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03257_ ) );
OAI211_X1 _10887_ ( .A(_03257_ ), .B(_02449_ ), .C1(_02455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03258_ ) );
OR2_X1 _10888_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03259_ ) );
OAI211_X1 _10889_ ( .A(_03259_ ), .B(fanout_net_27 ), .C1(_02455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03260_ ) );
NAND3_X1 _10890_ ( .A1(_03258_ ), .A2(_03260_ ), .A3(_02464_ ), .ZN(_03261_ ) );
MUX2_X1 _10891_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03262_ ) );
MUX2_X1 _10892_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03263_ ) );
MUX2_X1 _10893_ ( .A(_03262_ ), .B(_03263_ ), .S(_02449_ ), .Z(_03264_ ) );
OAI211_X1 _10894_ ( .A(_02686_ ), .B(_03261_ ), .C1(_03264_ ), .C2(_02465_ ), .ZN(_03265_ ) );
OR2_X1 _10895_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03266_ ) );
OAI211_X1 _10896_ ( .A(_03266_ ), .B(_02469_ ), .C1(_02501_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03267_ ) );
NOR2_X1 _10897_ ( .A1(_02455_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03268_ ) );
OAI21_X1 _10898_ ( .A(fanout_net_27 ), .B1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03269_ ) );
OAI211_X1 _10899_ ( .A(_03267_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_03268_ ), .C2(_03269_ ), .ZN(_03270_ ) );
MUX2_X1 _10900_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03271_ ) );
MUX2_X1 _10901_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03272_ ) );
MUX2_X1 _10902_ ( .A(_03271_ ), .B(_03272_ ), .S(fanout_net_27 ), .Z(_03273_ ) );
OAI211_X1 _10903_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03270_ ), .C1(_03273_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03274_ ) );
OAI211_X1 _10904_ ( .A(_03265_ ), .B(_03274_ ), .C1(_02487_ ), .C2(_02491_ ), .ZN(_03275_ ) );
NAND2_X1 _10905_ ( .A1(_03256_ ), .A2(_03275_ ), .ZN(_03276_ ) );
INV_X1 _10906_ ( .A(\ID_EX_imm [29] ), .ZN(_03277_ ) );
XNOR2_X1 _10907_ ( .A(_03276_ ), .B(_03277_ ), .ZN(_03278_ ) );
AND2_X1 _10908_ ( .A1(_03255_ ), .A2(_03278_ ), .ZN(_03279_ ) );
AOI21_X1 _10909_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_03251_ ), .B2(_03252_ ), .ZN(_03280_ ) );
NAND2_X1 _10910_ ( .A1(_03278_ ), .A2(_03280_ ), .ZN(_03281_ ) );
INV_X1 _10911_ ( .A(_03276_ ), .ZN(_03282_ ) );
OAI21_X1 _10912_ ( .A(_03281_ ), .B1(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_03282_ ), .ZN(_03283_ ) );
NOR2_X1 _10913_ ( .A1(_03279_ ), .A2(_03283_ ), .ZN(_03284_ ) );
MUX2_X1 _10914_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03285_ ) );
AND2_X1 _10915_ ( .A1(_03285_ ), .A2(fanout_net_27 ), .ZN(_03286_ ) );
MUX2_X1 _10916_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03287_ ) );
AND2_X1 _10917_ ( .A1(_03287_ ), .A2(_02450_ ), .ZN(_03288_ ) );
NOR3_X1 _10918_ ( .A1(_03286_ ), .A2(_03288_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03289_ ) );
AND2_X1 _10919_ ( .A1(_03159_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03290_ ) );
AOI211_X1 _10920_ ( .A(_02450_ ), .B(_03290_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03291_ ) );
AND2_X1 _10921_ ( .A1(_03159_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03292_ ) );
AOI211_X1 _10922_ ( .A(fanout_net_27 ), .B(_03292_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03293_ ) );
OAI21_X1 _10923_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B1(_03291_ ), .B2(_03293_ ), .ZN(_03294_ ) );
NAND2_X1 _10924_ ( .A1(_03294_ ), .A2(_02686_ ), .ZN(_03295_ ) );
INV_X1 _10925_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03296_ ) );
INV_X1 _10926_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03297_ ) );
MUX2_X1 _10927_ ( .A(_03296_ ), .B(_03297_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03298_ ) );
NOR2_X1 _10928_ ( .A1(_03298_ ), .A2(fanout_net_27 ), .ZN(_03299_ ) );
MUX2_X1 _10929_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03300_ ) );
AOI21_X1 _10930_ ( .A(_03299_ ), .B1(fanout_net_27 ), .B2(_03300_ ), .ZN(_03301_ ) );
MUX2_X1 _10931_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03302_ ) );
AND2_X1 _10932_ ( .A1(_03302_ ), .A2(_02470_ ), .ZN(_03303_ ) );
MUX2_X1 _10933_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03304_ ) );
AOI21_X1 _10934_ ( .A(_03303_ ), .B1(fanout_net_27 ), .B2(_03304_ ), .ZN(_03305_ ) );
MUX2_X1 _10935_ ( .A(_03301_ ), .B(_03305_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(_03306_ ) );
OAI221_X1 _10936_ ( .A(_02442_ ), .B1(_03289_ ), .B2(_03295_ ), .C1(_03306_ ), .C2(_02686_ ), .ZN(_03307_ ) );
OR3_X1 _10937_ ( .A1(_02488_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02492_ ), .ZN(_03308_ ) );
AND2_X1 _10938_ ( .A1(_03307_ ), .A2(_03308_ ), .ZN(_03309_ ) );
BUF_X2 _10939_ ( .A(_03309_ ), .Z(_03310_ ) );
INV_X1 _10940_ ( .A(\ID_EX_imm [30] ), .ZN(_03311_ ) );
XNOR2_X1 _10941_ ( .A(_03310_ ), .B(_03311_ ), .ZN(_03312_ ) );
OR2_X1 _10942_ ( .A1(_03284_ ), .A2(_03312_ ), .ZN(_03313_ ) );
OR2_X1 _10943_ ( .A1(_03310_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03314_ ) );
NAND2_X1 _10944_ ( .A1(_03313_ ), .A2(_03314_ ), .ZN(_03315_ ) );
OR3_X1 _10945_ ( .A1(_02488_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02492_ ), .ZN(_03316_ ) );
OR2_X1 _10946_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03317_ ) );
OAI211_X1 _10947_ ( .A(_03317_ ), .B(_02450_ ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03318_ ) );
OR2_X1 _10948_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03319_ ) );
OAI211_X1 _10949_ ( .A(_03319_ ), .B(fanout_net_27 ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03320_ ) );
NAND3_X1 _10950_ ( .A1(_03318_ ), .A2(_03320_ ), .A3(_02465_ ), .ZN(_03321_ ) );
MUX2_X1 _10951_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03322_ ) );
MUX2_X1 _10952_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03323_ ) );
MUX2_X1 _10953_ ( .A(_03322_ ), .B(_03323_ ), .S(_02470_ ), .Z(_03324_ ) );
OAI211_X1 _10954_ ( .A(_02686_ ), .B(_03321_ ), .C1(_03324_ ), .C2(_02465_ ), .ZN(_03325_ ) );
OR2_X1 _10955_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03326_ ) );
OAI211_X1 _10956_ ( .A(_03326_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03327_ ) );
OR2_X1 _10957_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03328_ ) );
OAI211_X1 _10958_ ( .A(_03328_ ), .B(_02450_ ), .C1(_02456_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03329_ ) );
NAND3_X1 _10959_ ( .A1(_03327_ ), .A2(_03329_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03330_ ) );
MUX2_X1 _10960_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03331_ ) );
MUX2_X1 _10961_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03332_ ) );
MUX2_X1 _10962_ ( .A(_03331_ ), .B(_03332_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03333_ ) );
OAI211_X1 _10963_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03330_ ), .C1(_03333_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03334_ ) );
OAI211_X1 _10964_ ( .A(_03325_ ), .B(_03334_ ), .C1(_02488_ ), .C2(_02492_ ), .ZN(_03335_ ) );
NAND2_X1 _10965_ ( .A1(_03316_ ), .A2(_03335_ ), .ZN(_03336_ ) );
BUF_X2 _10966_ ( .A(_03336_ ), .Z(_03337_ ) );
XOR2_X1 _10967_ ( .A(_03337_ ), .B(\ID_EX_imm [31] ), .Z(_03338_ ) );
XNOR2_X1 _10968_ ( .A(_03315_ ), .B(_03338_ ), .ZN(_03339_ ) );
AND2_X1 _10969_ ( .A1(_02407_ ), .A2(\ID_EX_typ [6] ), .ZN(_03340_ ) );
BUF_X4 _10970_ ( .A(_03340_ ), .Z(_03341_ ) );
AND2_X2 _10971_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03342_ ) );
AND2_X2 _10972_ ( .A1(_03342_ ), .A2(\ID_EX_typ [7] ), .ZN(_03343_ ) );
NOR2_X1 _10973_ ( .A1(_03341_ ), .A2(_03343_ ), .ZN(_03344_ ) );
INV_X1 _10974_ ( .A(_03344_ ), .ZN(_03345_ ) );
BUF_X4 _10975_ ( .A(_03345_ ), .Z(_03346_ ) );
NOR2_X1 _10976_ ( .A1(_03339_ ), .A2(_03346_ ), .ZN(_00097_ ) );
XNOR2_X1 _10977_ ( .A(_03284_ ), .B(_03312_ ), .ZN(_03347_ ) );
NOR2_X1 _10978_ ( .A1(_03347_ ), .A2(_03346_ ), .ZN(_00098_ ) );
AOI21_X1 _10979_ ( .A(_02709_ ), .B1(_03122_ ), .B2(_03128_ ), .ZN(_03348_ ) );
INV_X1 _10980_ ( .A(_03138_ ), .ZN(_03349_ ) );
NOR2_X1 _10981_ ( .A1(_03348_ ), .A2(_03349_ ), .ZN(_03350_ ) );
INV_X1 _10982_ ( .A(_03350_ ), .ZN(_03351_ ) );
AND2_X1 _10983_ ( .A1(_03351_ ), .A2(_02600_ ), .ZN(_03352_ ) );
OR2_X1 _10984_ ( .A1(_03352_ ), .A2(_03140_ ), .ZN(_03353_ ) );
XNOR2_X1 _10985_ ( .A(_03353_ ), .B(_02577_ ), .ZN(_03354_ ) );
NOR2_X1 _10986_ ( .A1(_03354_ ), .A2(_03346_ ), .ZN(_00099_ ) );
XOR2_X1 _10987_ ( .A(_03350_ ), .B(_02600_ ), .Z(_03355_ ) );
NOR2_X1 _10988_ ( .A1(_03355_ ), .A2(_03346_ ), .ZN(_00100_ ) );
INV_X1 _10989_ ( .A(_02708_ ), .ZN(_03356_ ) );
AOI21_X1 _10990_ ( .A(_03356_ ), .B1(_03122_ ), .B2(_03128_ ), .ZN(_03357_ ) );
AND2_X1 _10991_ ( .A1(_03357_ ), .A2(_02684_ ), .ZN(_03358_ ) );
NOR2_X1 _10992_ ( .A1(_03358_ ), .A2(_03133_ ), .ZN(_03359_ ) );
INV_X1 _10993_ ( .A(_02628_ ), .ZN(_03360_ ) );
NOR2_X1 _10994_ ( .A1(_03359_ ), .A2(_03360_ ), .ZN(_03361_ ) );
OR2_X1 _10995_ ( .A1(_03361_ ), .A2(_03135_ ), .ZN(_03362_ ) );
XNOR2_X1 _10996_ ( .A(_03362_ ), .B(_02657_ ), .ZN(_03363_ ) );
NOR2_X1 _10997_ ( .A1(_03363_ ), .A2(_03346_ ), .ZN(_00101_ ) );
XNOR2_X1 _10998_ ( .A(_03359_ ), .B(_03360_ ), .ZN(_03364_ ) );
NOR2_X1 _10999_ ( .A1(_03364_ ), .A2(_03346_ ), .ZN(_00102_ ) );
OR2_X1 _11000_ ( .A1(_03357_ ), .A2(_03130_ ), .ZN(_03365_ ) );
XNOR2_X1 _11001_ ( .A(_03365_ ), .B(_02684_ ), .ZN(_03366_ ) );
NOR2_X1 _11002_ ( .A1(_03366_ ), .A2(_03346_ ), .ZN(_00103_ ) );
AND3_X1 _11003_ ( .A1(_03122_ ), .A2(_03128_ ), .A3(_03356_ ), .ZN(_03367_ ) );
NOR3_X1 _11004_ ( .A1(_03367_ ), .A2(_03357_ ), .A3(_03345_ ), .ZN(_00104_ ) );
INV_X1 _11005_ ( .A(_03072_ ), .ZN(_03368_ ) );
NOR4_X1 _11006_ ( .A1(_03025_ ), .A2(_03047_ ), .A3(_03048_ ), .A4(_03368_ ), .ZN(_03369_ ) );
OR2_X1 _11007_ ( .A1(_03124_ ), .A2(_03048_ ), .ZN(_03370_ ) );
OAI21_X1 _11008_ ( .A(_03120_ ), .B1(_03369_ ), .B2(_03370_ ), .ZN(_03371_ ) );
NAND2_X1 _11009_ ( .A1(_03118_ ), .A2(\ID_EX_imm [14] ), .ZN(_03372_ ) );
NAND2_X1 _11010_ ( .A1(_03371_ ), .A2(_03372_ ), .ZN(_03373_ ) );
XNOR2_X1 _11011_ ( .A(_03373_ ), .B(_03095_ ), .ZN(_03374_ ) );
NOR2_X1 _11012_ ( .A1(_03374_ ), .A2(_03346_ ), .ZN(_00105_ ) );
OR3_X1 _11013_ ( .A1(_03369_ ), .A2(_03120_ ), .A3(_03370_ ), .ZN(_03375_ ) );
AND3_X1 _11014_ ( .A1(_03375_ ), .A2(_03344_ ), .A3(_03371_ ), .ZN(_00106_ ) );
OAI21_X1 _11015_ ( .A(_03072_ ), .B1(_03016_ ), .B2(_03024_ ), .ZN(_03376_ ) );
NAND2_X1 _11016_ ( .A1(_03376_ ), .A2(_03123_ ), .ZN(_03377_ ) );
XNOR2_X1 _11017_ ( .A(_03377_ ), .B(_03049_ ), .ZN(_03378_ ) );
NOR2_X1 _11018_ ( .A1(_03378_ ), .A2(_03346_ ), .ZN(_00107_ ) );
XNOR2_X1 _11019_ ( .A(_03025_ ), .B(_03368_ ), .ZN(_03379_ ) );
NOR2_X1 _11020_ ( .A1(_03379_ ), .A2(_03346_ ), .ZN(_00108_ ) );
NOR2_X1 _11021_ ( .A1(_03255_ ), .A2(_03280_ ), .ZN(_03380_ ) );
XOR2_X1 _11022_ ( .A(_03380_ ), .B(_03278_ ), .Z(_03381_ ) );
BUF_X4 _11023_ ( .A(_03345_ ), .Z(_03382_ ) );
NOR2_X1 _11024_ ( .A1(_03381_ ), .A2(_03382_ ), .ZN(_00109_ ) );
XNOR2_X1 _11025_ ( .A(_03231_ ), .B(_03254_ ), .ZN(_03383_ ) );
NOR2_X1 _11026_ ( .A1(_03383_ ), .A2(_03382_ ), .ZN(_00110_ ) );
NAND3_X1 _11027_ ( .A1(_03200_ ), .A2(_03223_ ), .A3(_03225_ ), .ZN(_03384_ ) );
NAND2_X1 _11028_ ( .A1(_03384_ ), .A2(_03228_ ), .ZN(_03385_ ) );
XNOR2_X1 _11029_ ( .A(_03385_ ), .B(_02496_ ), .ZN(_03386_ ) );
NOR2_X1 _11030_ ( .A1(_03386_ ), .A2(_03382_ ), .ZN(_00111_ ) );
NAND2_X1 _11031_ ( .A1(_03200_ ), .A2(_03225_ ), .ZN(_03387_ ) );
XNOR2_X1 _11032_ ( .A(_03387_ ), .B(_03222_ ), .ZN(_03388_ ) );
NOR2_X1 _11033_ ( .A1(_03388_ ), .A2(_03382_ ), .ZN(_00112_ ) );
NAND2_X1 _11034_ ( .A1(_03199_ ), .A2(_03225_ ), .ZN(_03389_ ) );
XNOR2_X1 _11035_ ( .A(_03177_ ), .B(_03389_ ), .ZN(_03390_ ) );
NOR2_X1 _11036_ ( .A1(_03390_ ), .A2(_03382_ ), .ZN(_00113_ ) );
XNOR2_X1 _11037_ ( .A(_03147_ ), .B(_03174_ ), .ZN(_03391_ ) );
NOR2_X1 _11038_ ( .A1(_03391_ ), .A2(_03382_ ), .ZN(_00114_ ) );
AND2_X1 _11039_ ( .A1(_03351_ ), .A2(_02601_ ), .ZN(_03392_ ) );
OAI21_X1 _11040_ ( .A(_02524_ ), .B1(_03392_ ), .B2(_03143_ ), .ZN(_03393_ ) );
AND2_X1 _11041_ ( .A1(_02522_ ), .A2(\ID_EX_imm [22] ), .ZN(_03394_ ) );
INV_X1 _11042_ ( .A(_03394_ ), .ZN(_03395_ ) );
AND4_X1 _11043_ ( .A1(_02546_ ), .A2(_03393_ ), .A3(_02549_ ), .A4(_03395_ ), .ZN(_03396_ ) );
AOI22_X1 _11044_ ( .A1(_03393_ ), .A2(_03395_ ), .B1(_02546_ ), .B2(_02549_ ), .ZN(_03397_ ) );
NOR2_X1 _11045_ ( .A1(_03396_ ), .A2(_03397_ ), .ZN(_03398_ ) );
NOR2_X1 _11046_ ( .A1(_03398_ ), .A2(_03382_ ), .ZN(_00115_ ) );
OR3_X1 _11047_ ( .A1(_03392_ ), .A2(_02524_ ), .A3(_03143_ ), .ZN(_03399_ ) );
AND3_X1 _11048_ ( .A1(_03399_ ), .A2(_03344_ ), .A3(_03393_ ), .ZN(_00116_ ) );
BUF_X2 _11049_ ( .A(_01886_ ), .Z(_03400_ ) );
INV_X1 _11050_ ( .A(fanout_net_16 ), .ZN(_03401_ ) );
BUF_X4 _11051_ ( .A(_03401_ ), .Z(_03402_ ) );
CLKBUF_X2 _11052_ ( .A(_03402_ ), .Z(_03403_ ) );
AND3_X1 _11053_ ( .A1(_03400_ ), .A2(_03403_ ), .A3(\ID_EX_rd [4] ), .ZN(_00117_ ) );
AND3_X1 _11054_ ( .A1(_03400_ ), .A2(_03403_ ), .A3(\ID_EX_rd [3] ), .ZN(_00118_ ) );
AND3_X1 _11055_ ( .A1(_03400_ ), .A2(_03403_ ), .A3(\ID_EX_rd [2] ), .ZN(_00119_ ) );
AND3_X1 _11056_ ( .A1(_03400_ ), .A2(_03403_ ), .A3(\ID_EX_rd [1] ), .ZN(_00120_ ) );
AND3_X1 _11057_ ( .A1(_01914_ ), .A2(_03403_ ), .A3(\ID_EX_rd [0] ), .ZN(_00121_ ) );
INV_X1 _11058_ ( .A(\ID_EX_pc [31] ), .ZN(_03404_ ) );
NOR3_X1 _11059_ ( .A1(_03404_ ), .A2(fanout_net_2 ), .A3(fanout_net_16 ), .ZN(_00122_ ) );
INV_X1 _11060_ ( .A(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_03405_ ) );
BUF_X4 _11061_ ( .A(_03405_ ), .Z(_03406_ ) );
XOR2_X1 _11062_ ( .A(\ID_EX_pc [25] ), .B(\ID_EX_imm [25] ), .Z(_03407_ ) );
XOR2_X1 _11063_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_03408_ ) );
NOR2_X1 _11064_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03409_ ) );
XOR2_X1 _11065_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_03410_ ) );
NOR2_X1 _11066_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03411_ ) );
XOR2_X1 _11067_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_imm [3] ), .Z(_03412_ ) );
AND2_X1 _11068_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_03413_ ) );
AND2_X1 _11069_ ( .A1(_03412_ ), .A2(_03413_ ), .ZN(_03414_ ) );
AOI21_X1 _11070_ ( .A(_03414_ ), .B1(\ID_EX_pc [3] ), .B2(\ID_EX_imm [3] ), .ZN(_03415_ ) );
XOR2_X1 _11071_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_03416_ ) );
XOR2_X1 _11072_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_03417_ ) );
AND2_X1 _11073_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_03418_ ) );
AND2_X1 _11074_ ( .A1(_03417_ ), .A2(_03418_ ), .ZN(_03419_ ) );
AND2_X1 _11075_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_03420_ ) );
OAI211_X1 _11076_ ( .A(_03416_ ), .B(_03412_ ), .C1(_03419_ ), .C2(_03420_ ), .ZN(_03421_ ) );
NAND2_X1 _11077_ ( .A1(_03415_ ), .A2(_03421_ ), .ZN(_03422_ ) );
XOR2_X1 _11078_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_03423_ ) );
NAND2_X1 _11079_ ( .A1(_03422_ ), .A2(_03423_ ), .ZN(_03424_ ) );
NAND2_X1 _11080_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03425_ ) );
AOI21_X1 _11081_ ( .A(_03411_ ), .B1(_03424_ ), .B2(_03425_ ), .ZN(_03426_ ) );
AND2_X1 _11082_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03427_ ) );
OAI21_X1 _11083_ ( .A(_03410_ ), .B1(_03426_ ), .B2(_03427_ ), .ZN(_03428_ ) );
NAND2_X1 _11084_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03429_ ) );
AOI21_X1 _11085_ ( .A(_03409_ ), .B1(_03428_ ), .B2(_03429_ ), .ZN(_03430_ ) );
AND2_X1 _11086_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03431_ ) );
OR2_X1 _11087_ ( .A1(_03430_ ), .A2(_03431_ ), .ZN(_03432_ ) );
XOR2_X1 _11088_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_03433_ ) );
XOR2_X1 _11089_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_03434_ ) );
AND2_X1 _11090_ ( .A1(_03433_ ), .A2(_03434_ ), .ZN(_03435_ ) );
XOR2_X1 _11091_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_03436_ ) );
XOR2_X1 _11092_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_03437_ ) );
AND2_X1 _11093_ ( .A1(_03436_ ), .A2(_03437_ ), .ZN(_03438_ ) );
AND3_X1 _11094_ ( .A1(_03432_ ), .A2(_03435_ ), .A3(_03438_ ), .ZN(_03439_ ) );
AND2_X1 _11095_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_03440_ ) );
AND2_X1 _11096_ ( .A1(_03433_ ), .A2(_03440_ ), .ZN(_03441_ ) );
AOI21_X1 _11097_ ( .A(_03441_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_03442_ ) );
AND2_X1 _11098_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_03443_ ) );
AND2_X1 _11099_ ( .A1(_03437_ ), .A2(_03443_ ), .ZN(_03444_ ) );
AOI21_X1 _11100_ ( .A(_03444_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_03445_ ) );
INV_X1 _11101_ ( .A(_03435_ ), .ZN(_03446_ ) );
OAI21_X1 _11102_ ( .A(_03442_ ), .B1(_03445_ ), .B2(_03446_ ), .ZN(_03447_ ) );
OR2_X1 _11103_ ( .A1(_03439_ ), .A2(_03447_ ), .ZN(_03448_ ) );
XOR2_X1 _11104_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_03449_ ) );
XOR2_X1 _11105_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_03450_ ) );
AND2_X1 _11106_ ( .A1(_03449_ ), .A2(_03450_ ), .ZN(_03451_ ) );
XOR2_X1 _11107_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_03452_ ) );
INV_X1 _11108_ ( .A(_03452_ ), .ZN(_03453_ ) );
XNOR2_X1 _11109_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .ZN(_03454_ ) );
NOR2_X1 _11110_ ( .A1(_03453_ ), .A2(_03454_ ), .ZN(_03455_ ) );
AND3_X1 _11111_ ( .A1(_03448_ ), .A2(_03451_ ), .A3(_03455_ ), .ZN(_03456_ ) );
AND2_X1 _11112_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_03457_ ) );
AND2_X1 _11113_ ( .A1(_03449_ ), .A2(_03457_ ), .ZN(_03458_ ) );
AOI21_X1 _11114_ ( .A(_03458_ ), .B1(\ID_EX_pc [15] ), .B2(\ID_EX_imm [15] ), .ZN(_03459_ ) );
INV_X1 _11115_ ( .A(_03451_ ), .ZN(_03460_ ) );
NAND2_X1 _11116_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_03461_ ) );
NOR2_X1 _11117_ ( .A1(_03454_ ), .A2(_03461_ ), .ZN(_03462_ ) );
AOI21_X1 _11118_ ( .A(_03462_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_03463_ ) );
OAI21_X1 _11119_ ( .A(_03459_ ), .B1(_03460_ ), .B2(_03463_ ), .ZN(_03464_ ) );
OR2_X1 _11120_ ( .A1(_03456_ ), .A2(_03464_ ), .ZN(_03465_ ) );
XOR2_X1 _11121_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_03466_ ) );
XOR2_X1 _11122_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_03467_ ) );
AND2_X1 _11123_ ( .A1(_03466_ ), .A2(_03467_ ), .ZN(_03468_ ) );
XOR2_X1 _11124_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_03469_ ) );
XOR2_X1 _11125_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_03470_ ) );
AND2_X1 _11126_ ( .A1(_03469_ ), .A2(_03470_ ), .ZN(_03471_ ) );
AND3_X1 _11127_ ( .A1(_03465_ ), .A2(_03468_ ), .A3(_03471_ ), .ZN(_03472_ ) );
AND2_X1 _11128_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_03473_ ) );
AND2_X1 _11129_ ( .A1(_03466_ ), .A2(_03473_ ), .ZN(_03474_ ) );
AOI21_X1 _11130_ ( .A(_03474_ ), .B1(\ID_EX_pc [19] ), .B2(\ID_EX_imm [19] ), .ZN(_03475_ ) );
AND2_X1 _11131_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_03476_ ) );
AND2_X1 _11132_ ( .A1(_03470_ ), .A2(_03476_ ), .ZN(_03477_ ) );
AOI21_X1 _11133_ ( .A(_03477_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_03478_ ) );
INV_X1 _11134_ ( .A(_03468_ ), .ZN(_03479_ ) );
OAI21_X1 _11135_ ( .A(_03475_ ), .B1(_03478_ ), .B2(_03479_ ), .ZN(_03480_ ) );
OR2_X1 _11136_ ( .A1(_03472_ ), .A2(_03480_ ), .ZN(_03481_ ) );
XOR2_X1 _11137_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_03482_ ) );
XOR2_X1 _11138_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_03483_ ) );
AND2_X1 _11139_ ( .A1(_03482_ ), .A2(_03483_ ), .ZN(_03484_ ) );
XOR2_X1 _11140_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_03485_ ) );
XOR2_X1 _11141_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_03486_ ) );
AND2_X1 _11142_ ( .A1(_03485_ ), .A2(_03486_ ), .ZN(_03487_ ) );
AND3_X1 _11143_ ( .A1(_03481_ ), .A2(_03484_ ), .A3(_03487_ ), .ZN(_03488_ ) );
AND2_X1 _11144_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_03489_ ) );
AND2_X1 _11145_ ( .A1(_03482_ ), .A2(_03489_ ), .ZN(_03490_ ) );
AOI21_X1 _11146_ ( .A(_03490_ ), .B1(\ID_EX_pc [23] ), .B2(\ID_EX_imm [23] ), .ZN(_03491_ ) );
AND3_X1 _11147_ ( .A1(_03485_ ), .A2(\ID_EX_pc [20] ), .A3(\ID_EX_imm [20] ), .ZN(_03492_ ) );
AOI21_X1 _11148_ ( .A(_03492_ ), .B1(\ID_EX_pc [21] ), .B2(\ID_EX_imm [21] ), .ZN(_03493_ ) );
INV_X1 _11149_ ( .A(_03484_ ), .ZN(_03494_ ) );
OAI21_X1 _11150_ ( .A(_03491_ ), .B1(_03493_ ), .B2(_03494_ ), .ZN(_03495_ ) );
OAI211_X1 _11151_ ( .A(_03407_ ), .B(_03408_ ), .C1(_03488_ ), .C2(_03495_ ), .ZN(_03496_ ) );
AND2_X1 _11152_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_03497_ ) );
AND2_X1 _11153_ ( .A1(_03407_ ), .A2(_03497_ ), .ZN(_03498_ ) );
AOI21_X1 _11154_ ( .A(_03498_ ), .B1(\ID_EX_pc [25] ), .B2(\ID_EX_imm [25] ), .ZN(_03499_ ) );
NAND2_X1 _11155_ ( .A1(_03496_ ), .A2(_03499_ ), .ZN(_03500_ ) );
XOR2_X1 _11156_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_03501_ ) );
XOR2_X1 _11157_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_03502_ ) );
NAND3_X1 _11158_ ( .A1(_03500_ ), .A2(_03501_ ), .A3(_03502_ ), .ZN(_03503_ ) );
AND3_X1 _11159_ ( .A1(_03501_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_03504_ ) );
AOI21_X1 _11160_ ( .A(_03504_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_03505_ ) );
NAND2_X1 _11161_ ( .A1(_03503_ ), .A2(_03505_ ), .ZN(_03506_ ) );
XOR2_X1 _11162_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_03507_ ) );
NAND2_X1 _11163_ ( .A1(_03506_ ), .A2(_03507_ ), .ZN(_03508_ ) );
NAND2_X1 _11164_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_03509_ ) );
INV_X1 _11165_ ( .A(\ID_EX_pc [29] ), .ZN(_03510_ ) );
AOI22_X1 _11166_ ( .A1(_03508_ ), .A2(_03509_ ), .B1(_03510_ ), .B2(_03277_ ), .ZN(_03511_ ) );
AND2_X1 _11167_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_03512_ ) );
OR2_X1 _11168_ ( .A1(_03511_ ), .A2(_03512_ ), .ZN(_03513_ ) );
XOR2_X1 _11169_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_03514_ ) );
XOR2_X1 _11170_ ( .A(_03513_ ), .B(_03514_ ), .Z(_03515_ ) );
BUF_X2 _11171_ ( .A(_02419_ ), .Z(_03516_ ) );
CLKBUF_X2 _11172_ ( .A(_02415_ ), .Z(_03517_ ) );
AND3_X1 _11173_ ( .A1(_03515_ ), .A2(_03516_ ), .A3(_03517_ ), .ZN(_03518_ ) );
NOR2_X1 _11174_ ( .A1(_02395_ ), .A2(fanout_net_16 ), .ZN(_03519_ ) );
XOR2_X1 _11175_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .Z(_03520_ ) );
INV_X1 _11176_ ( .A(_03520_ ), .ZN(_03521_ ) );
XNOR2_X1 _11177_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_03522_ ) );
XNOR2_X1 _11178_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_03523_ ) );
AND2_X1 _11179_ ( .A1(_03522_ ), .A2(_03523_ ), .ZN(_03524_ ) );
XOR2_X1 _11180_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .Z(_03525_ ) );
XOR2_X1 _11181_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .Z(_03526_ ) );
NOR2_X1 _11182_ ( .A1(_03525_ ), .A2(_03526_ ), .ZN(_03527_ ) );
XNOR2_X1 _11183_ ( .A(\EX_LS_dest_csreg_mem [1] ), .B(\ID_EX_csr [1] ), .ZN(_03528_ ) );
XNOR2_X1 _11184_ ( .A(fanout_net_4 ), .B(\ID_EX_csr [0] ), .ZN(_03529_ ) );
AND2_X1 _11185_ ( .A1(_03528_ ), .A2(_03529_ ), .ZN(_03530_ ) );
XNOR2_X1 _11186_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_03531_ ) );
XNOR2_X1 _11187_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_03532_ ) );
AND2_X1 _11188_ ( .A1(_03531_ ), .A2(_03532_ ), .ZN(_03533_ ) );
AND4_X1 _11189_ ( .A1(_03524_ ), .A2(_03527_ ), .A3(_03530_ ), .A4(_03533_ ), .ZN(_03534_ ) );
XNOR2_X1 _11190_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_03535_ ) );
XNOR2_X1 _11191_ ( .A(\EX_LS_dest_csreg_mem [8] ), .B(\ID_EX_csr [8] ), .ZN(_03536_ ) );
XNOR2_X1 _11192_ ( .A(\EX_LS_dest_csreg_mem [9] ), .B(\ID_EX_csr [9] ), .ZN(_03537_ ) );
AND2_X1 _11193_ ( .A1(_03536_ ), .A2(_03537_ ), .ZN(_03538_ ) );
AND4_X2 _11194_ ( .A1(_03521_ ), .A2(_03534_ ), .A3(_03535_ ), .A4(_03538_ ), .ZN(_03539_ ) );
INV_X1 _11195_ ( .A(_03539_ ), .ZN(_03540_ ) );
INV_X1 _11196_ ( .A(_02423_ ), .ZN(_03541_ ) );
BUF_X4 _11197_ ( .A(_03541_ ), .Z(_03542_ ) );
NOR2_X1 _11198_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_03543_ ) );
INV_X1 _11199_ ( .A(\ID_EX_csr [5] ), .ZN(_03544_ ) );
AND2_X1 _11200_ ( .A1(_03543_ ), .A2(_03544_ ), .ZN(_03545_ ) );
NOR2_X1 _11201_ ( .A1(\ID_EX_csr [3] ), .A2(\ID_EX_csr [2] ), .ZN(_03546_ ) );
INV_X1 _11202_ ( .A(\ID_EX_csr [0] ), .ZN(_03547_ ) );
NOR2_X1 _11203_ ( .A1(_03547_ ), .A2(\ID_EX_csr [1] ), .ZN(_03548_ ) );
AND4_X1 _11204_ ( .A1(\ID_EX_csr [4] ), .A2(_03545_ ), .A3(_03546_ ), .A4(_03548_ ), .ZN(_03549_ ) );
AND2_X1 _11205_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_03550_ ) );
AND3_X1 _11206_ ( .A1(_03550_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_03551_ ) );
NAND2_X1 _11207_ ( .A1(_03549_ ), .A2(_03551_ ), .ZN(_03552_ ) );
INV_X1 _11208_ ( .A(\ID_EX_csr [6] ), .ZN(_03553_ ) );
NOR2_X1 _11209_ ( .A1(_03553_ ), .A2(\ID_EX_csr [7] ), .ZN(_03554_ ) );
NOR2_X1 _11210_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_03555_ ) );
AND4_X1 _11211_ ( .A1(_03546_ ), .A2(_03548_ ), .A3(_03554_ ), .A4(_03555_ ), .ZN(_03556_ ) );
BUF_X4 _11212_ ( .A(_03556_ ), .Z(_03557_ ) );
NOR2_X1 _11213_ ( .A1(\ID_EX_csr [10] ), .A2(\ID_EX_csr [11] ), .ZN(_03558_ ) );
AND2_X1 _11214_ ( .A1(_03550_ ), .A2(_03558_ ), .ZN(_03559_ ) );
BUF_X4 _11215_ ( .A(_03559_ ), .Z(_03560_ ) );
NAND3_X1 _11216_ ( .A1(_03557_ ), .A2(\mepc [30] ), .A3(_03560_ ), .ZN(_03561_ ) );
AND2_X2 _11217_ ( .A1(_03554_ ), .A2(_03555_ ), .ZN(_03562_ ) );
INV_X1 _11218_ ( .A(\ID_EX_csr [1] ), .ZN(_03563_ ) );
NOR2_X1 _11219_ ( .A1(_03563_ ), .A2(\ID_EX_csr [0] ), .ZN(_03564_ ) );
AND2_X1 _11220_ ( .A1(_03564_ ), .A2(_03546_ ), .ZN(_03565_ ) );
NAND4_X1 _11221_ ( .A1(_03562_ ), .A2(_03565_ ), .A3(\mycsreg.CSReg[3][30] ), .A4(_03560_ ), .ZN(_03566_ ) );
INV_X1 _11222_ ( .A(\ID_EX_csr [3] ), .ZN(_03567_ ) );
AND3_X1 _11223_ ( .A1(_03548_ ), .A2(_03567_ ), .A3(\ID_EX_csr [2] ), .ZN(_03568_ ) );
BUF_X4 _11224_ ( .A(_03568_ ), .Z(_03569_ ) );
AND2_X1 _11225_ ( .A1(_03543_ ), .A2(_03555_ ), .ZN(_03570_ ) );
NAND4_X1 _11226_ ( .A1(_03569_ ), .A2(\mtvec [30] ), .A3(_03560_ ), .A4(_03570_ ), .ZN(_03571_ ) );
NAND4_X1 _11227_ ( .A1(_03552_ ), .A2(_03561_ ), .A3(_03566_ ), .A4(_03571_ ), .ZN(_03572_ ) );
AND3_X2 _11228_ ( .A1(_03546_ ), .A2(_03563_ ), .A3(_03547_ ), .ZN(_03573_ ) );
BUF_X4 _11229_ ( .A(_03570_ ), .Z(_03574_ ) );
AND4_X1 _11230_ ( .A1(\mycsreg.CSReg[0][30] ), .A2(_03573_ ), .A3(_03560_ ), .A4(_03574_ ), .ZN(_03575_ ) );
OAI22_X1 _11231_ ( .A1(_03540_ ), .A2(_03542_ ), .B1(_03572_ ), .B2(_03575_ ), .ZN(_03576_ ) );
BUF_X4 _11232_ ( .A(_02423_ ), .Z(_03577_ ) );
NAND3_X1 _11233_ ( .A1(_03539_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_03577_ ), .ZN(_03578_ ) );
AND2_X1 _11234_ ( .A1(_03576_ ), .A2(_03578_ ), .ZN(_03579_ ) );
INV_X2 _11235_ ( .A(fanout_net_6 ), .ZN(_03580_ ) );
OR2_X1 _11236_ ( .A1(_03579_ ), .A2(_03580_ ), .ZN(_03581_ ) );
AND2_X1 _11237_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_03582_ ) );
AND2_X1 _11238_ ( .A1(_03582_ ), .A2(\ID_EX_pc [4] ), .ZN(_03583_ ) );
AND2_X1 _11239_ ( .A1(_03583_ ), .A2(\ID_EX_pc [5] ), .ZN(_03584_ ) );
AND2_X1 _11240_ ( .A1(_03584_ ), .A2(\ID_EX_pc [6] ), .ZN(_03585_ ) );
AND2_X1 _11241_ ( .A1(_03585_ ), .A2(\ID_EX_pc [7] ), .ZN(_03586_ ) );
AND2_X1 _11242_ ( .A1(_03586_ ), .A2(\ID_EX_pc [8] ), .ZN(_03587_ ) );
AND2_X2 _11243_ ( .A1(_03587_ ), .A2(\ID_EX_pc [9] ), .ZN(_03588_ ) );
AND3_X1 _11244_ ( .A1(_03588_ ), .A2(\ID_EX_pc [11] ), .A3(\ID_EX_pc [10] ), .ZN(_03589_ ) );
AND3_X1 _11245_ ( .A1(_03589_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_03590_ ) );
AND3_X1 _11246_ ( .A1(_03590_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_03591_ ) );
AND3_X1 _11247_ ( .A1(_03591_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_03592_ ) );
AND3_X1 _11248_ ( .A1(_03592_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_03593_ ) );
AND3_X1 _11249_ ( .A1(_03593_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_03594_ ) );
AND3_X1 _11250_ ( .A1(_03594_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_03595_ ) );
AND3_X1 _11251_ ( .A1(_03595_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_03596_ ) );
AND3_X1 _11252_ ( .A1(_03596_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_03597_ ) );
NAND3_X1 _11253_ ( .A1(_03597_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_03598_ ) );
INV_X1 _11254_ ( .A(\ID_EX_pc [30] ), .ZN(_03599_ ) );
XNOR2_X1 _11255_ ( .A(_03598_ ), .B(_03599_ ), .ZN(_03600_ ) );
INV_X1 _11256_ ( .A(_03515_ ), .ZN(_03601_ ) );
NOR2_X1 _11257_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_5 ), .ZN(_03602_ ) );
AND2_X1 _11258_ ( .A1(_03602_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_03603_ ) );
INV_X1 _11259_ ( .A(_03603_ ), .ZN(_03604_ ) );
INV_X1 _11260_ ( .A(fanout_net_43 ), .ZN(_03605_ ) );
BUF_X4 _11261_ ( .A(_03605_ ), .Z(_03606_ ) );
OR2_X1 _11262_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][19] ), .ZN(_03607_ ) );
INV_X1 _11263_ ( .A(fanout_net_39 ), .ZN(_03608_ ) );
BUF_X4 _11264_ ( .A(_03608_ ), .Z(_03609_ ) );
BUF_X4 _11265_ ( .A(_03609_ ), .Z(_03610_ ) );
INV_X1 _11266_ ( .A(fanout_net_31 ), .ZN(_03611_ ) );
BUF_X4 _11267_ ( .A(_03611_ ), .Z(_03612_ ) );
BUF_X4 _11268_ ( .A(_03612_ ), .Z(_03613_ ) );
OAI211_X1 _11269_ ( .A(_03607_ ), .B(_03610_ ), .C1(_03613_ ), .C2(\myreg.Reg[1][19] ), .ZN(_03614_ ) );
OR2_X1 _11270_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][19] ), .ZN(_03615_ ) );
OAI211_X1 _11271_ ( .A(_03615_ ), .B(fanout_net_39 ), .C1(_03613_ ), .C2(\myreg.Reg[3][19] ), .ZN(_03616_ ) );
INV_X1 _11272_ ( .A(fanout_net_42 ), .ZN(_03617_ ) );
BUF_X4 _11273_ ( .A(_03617_ ), .Z(_03618_ ) );
BUF_X4 _11274_ ( .A(_03618_ ), .Z(_03619_ ) );
NAND3_X1 _11275_ ( .A1(_03614_ ), .A2(_03616_ ), .A3(_03619_ ), .ZN(_03620_ ) );
MUX2_X1 _11276_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_31 ), .Z(_03621_ ) );
MUX2_X1 _11277_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_31 ), .Z(_03622_ ) );
MUX2_X1 _11278_ ( .A(_03621_ ), .B(_03622_ ), .S(_03610_ ), .Z(_03623_ ) );
BUF_X4 _11279_ ( .A(_03619_ ), .Z(_03624_ ) );
OAI211_X1 _11280_ ( .A(_03606_ ), .B(_03620_ ), .C1(_03623_ ), .C2(_03624_ ), .ZN(_03625_ ) );
OR2_X1 _11281_ ( .A1(_03612_ ), .A2(\myreg.Reg[13][19] ), .ZN(_03626_ ) );
OAI211_X1 _11282_ ( .A(_03626_ ), .B(_03610_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[12][19] ), .ZN(_03627_ ) );
OR2_X1 _11283_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][19] ), .ZN(_03628_ ) );
OAI211_X1 _11284_ ( .A(_03628_ ), .B(fanout_net_39 ), .C1(_03613_ ), .C2(\myreg.Reg[15][19] ), .ZN(_03629_ ) );
NAND3_X1 _11285_ ( .A1(_03627_ ), .A2(fanout_net_42 ), .A3(_03629_ ), .ZN(_03630_ ) );
MUX2_X1 _11286_ ( .A(\myreg.Reg[8][19] ), .B(\myreg.Reg[9][19] ), .S(fanout_net_31 ), .Z(_03631_ ) );
MUX2_X1 _11287_ ( .A(\myreg.Reg[10][19] ), .B(\myreg.Reg[11][19] ), .S(fanout_net_31 ), .Z(_03632_ ) );
MUX2_X1 _11288_ ( .A(_03631_ ), .B(_03632_ ), .S(fanout_net_39 ), .Z(_03633_ ) );
OAI211_X1 _11289_ ( .A(fanout_net_43 ), .B(_03630_ ), .C1(_03633_ ), .C2(fanout_net_42 ), .ZN(_03634_ ) );
NAND2_X1 _11290_ ( .A1(_03625_ ), .A2(_03634_ ), .ZN(_03635_ ) );
XOR2_X2 _11291_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .Z(_03636_ ) );
INV_X1 _11292_ ( .A(\ID_EX_rs2 [3] ), .ZN(_03637_ ) );
OAI22_X1 _11293_ ( .A1(\EX_LS_dest_reg [3] ), .A2(_03637_ ), .B1(_02430_ ), .B2(\ID_EX_rs2 [1] ), .ZN(_03638_ ) );
NOR2_X1 _11294_ ( .A1(_03636_ ), .A2(_03638_ ), .ZN(_03639_ ) );
NAND2_X1 _11295_ ( .A1(_03637_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_03640_ ) );
XNOR2_X1 _11296_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_03641_ ) );
NAND4_X2 _11297_ ( .A1(_03639_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y ), .A3(_03640_ ), .A4(_03641_ ), .ZN(_03642_ ) );
BUF_X4 _11298_ ( .A(_03642_ ), .Z(_03643_ ) );
BUF_X2 _11299_ ( .A(_03643_ ), .Z(_03644_ ) );
XNOR2_X1 _11300_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_03645_ ) );
NAND2_X1 _11301_ ( .A1(_02430_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_03646_ ) );
NAND4_X4 _11302_ ( .A1(_02426_ ), .A2(_02429_ ), .A3(_03645_ ), .A4(_03646_ ), .ZN(_03647_ ) );
BUF_X8 _11303_ ( .A(_03647_ ), .Z(_03648_ ) );
BUF_X2 _11304_ ( .A(_03648_ ), .Z(_03649_ ) );
OAI21_X1 _11305_ ( .A(_03635_ ), .B1(_03644_ ), .B2(_03649_ ), .ZN(_03650_ ) );
BUF_X8 _11306_ ( .A(_03647_ ), .Z(_03651_ ) );
INV_X1 _11307_ ( .A(\EX_LS_result_reg [19] ), .ZN(_03652_ ) );
BUF_X2 _11308_ ( .A(_03642_ ), .Z(_03653_ ) );
OR3_X1 _11309_ ( .A1(_03651_ ), .A2(_03652_ ), .A3(_03653_ ), .ZN(_03654_ ) );
AND2_X1 _11310_ ( .A1(_03650_ ), .A2(_03654_ ), .ZN(_03655_ ) );
INV_X1 _11311_ ( .A(_02655_ ), .ZN(_03656_ ) );
XNOR2_X1 _11312_ ( .A(_03655_ ), .B(_03656_ ), .ZN(_03657_ ) );
BUF_X2 _11313_ ( .A(_03651_ ), .Z(_03658_ ) );
BUF_X2 _11314_ ( .A(_03653_ ), .Z(_03659_ ) );
OR3_X1 _11315_ ( .A1(_03658_ ), .A2(\EX_LS_result_reg [18] ), .A3(_03659_ ), .ZN(_03660_ ) );
BUF_X4 _11316_ ( .A(_03606_ ), .Z(_03661_ ) );
BUF_X4 _11317_ ( .A(_03611_ ), .Z(_03662_ ) );
BUF_X2 _11318_ ( .A(_03662_ ), .Z(_03663_ ) );
BUF_X2 _11319_ ( .A(_03663_ ), .Z(_03664_ ) );
OR2_X1 _11320_ ( .A1(_03664_ ), .A2(\myreg.Reg[3][18] ), .ZN(_03665_ ) );
OAI211_X1 _11321_ ( .A(_03665_ ), .B(fanout_net_39 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[2][18] ), .ZN(_03666_ ) );
BUF_X4 _11322_ ( .A(_03624_ ), .Z(_03667_ ) );
OR2_X1 _11323_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][18] ), .ZN(_03668_ ) );
BUF_X4 _11324_ ( .A(_03610_ ), .Z(_03669_ ) );
BUF_X4 _11325_ ( .A(_03669_ ), .Z(_03670_ ) );
BUF_X4 _11326_ ( .A(_03613_ ), .Z(_03671_ ) );
BUF_X4 _11327_ ( .A(_03671_ ), .Z(_03672_ ) );
OAI211_X1 _11328_ ( .A(_03668_ ), .B(_03670_ ), .C1(_03672_ ), .C2(\myreg.Reg[1][18] ), .ZN(_03673_ ) );
NAND3_X1 _11329_ ( .A1(_03666_ ), .A2(_03667_ ), .A3(_03673_ ), .ZN(_03674_ ) );
MUX2_X1 _11330_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_31 ), .Z(_03675_ ) );
MUX2_X1 _11331_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_31 ), .Z(_03676_ ) );
BUF_X4 _11332_ ( .A(_03610_ ), .Z(_03677_ ) );
MUX2_X1 _11333_ ( .A(_03675_ ), .B(_03676_ ), .S(_03677_ ), .Z(_03678_ ) );
OAI211_X1 _11334_ ( .A(_03661_ ), .B(_03674_ ), .C1(_03678_ ), .C2(_03667_ ), .ZN(_03679_ ) );
OR2_X1 _11335_ ( .A1(_03664_ ), .A2(\myreg.Reg[15][18] ), .ZN(_03680_ ) );
OAI211_X1 _11336_ ( .A(_03680_ ), .B(fanout_net_39 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[14][18] ), .ZN(_03681_ ) );
OR2_X1 _11337_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[12][18] ), .ZN(_03682_ ) );
OAI211_X1 _11338_ ( .A(_03682_ ), .B(_03670_ ), .C1(_03672_ ), .C2(\myreg.Reg[13][18] ), .ZN(_03683_ ) );
NAND3_X1 _11339_ ( .A1(_03681_ ), .A2(fanout_net_42 ), .A3(_03683_ ), .ZN(_03684_ ) );
MUX2_X1 _11340_ ( .A(\myreg.Reg[8][18] ), .B(\myreg.Reg[9][18] ), .S(fanout_net_31 ), .Z(_03685_ ) );
MUX2_X1 _11341_ ( .A(\myreg.Reg[10][18] ), .B(\myreg.Reg[11][18] ), .S(fanout_net_31 ), .Z(_03686_ ) );
MUX2_X1 _11342_ ( .A(_03685_ ), .B(_03686_ ), .S(fanout_net_39 ), .Z(_03687_ ) );
OAI211_X1 _11343_ ( .A(fanout_net_43 ), .B(_03684_ ), .C1(_03687_ ), .C2(fanout_net_42 ), .ZN(_03688_ ) );
BUF_X8 _11344_ ( .A(_03658_ ), .Z(_03689_ ) );
BUF_X2 _11345_ ( .A(_03659_ ), .Z(_03690_ ) );
OAI211_X1 _11346_ ( .A(_03679_ ), .B(_03688_ ), .C1(_03689_ ), .C2(_03690_ ), .ZN(_03691_ ) );
NAND2_X1 _11347_ ( .A1(_03660_ ), .A2(_03691_ ), .ZN(_03692_ ) );
XOR2_X1 _11348_ ( .A(_03692_ ), .B(_02626_ ), .Z(_03693_ ) );
AND2_X1 _11349_ ( .A1(_03657_ ), .A2(_03693_ ), .ZN(_03694_ ) );
INV_X1 _11350_ ( .A(_02682_ ), .ZN(_03695_ ) );
OR2_X1 _11351_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][17] ), .ZN(_03696_ ) );
OAI211_X1 _11352_ ( .A(_03696_ ), .B(_03669_ ), .C1(_03664_ ), .C2(\myreg.Reg[9][17] ), .ZN(_03697_ ) );
OR2_X1 _11353_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[10][17] ), .ZN(_03698_ ) );
BUF_X4 _11354_ ( .A(_03662_ ), .Z(_03699_ ) );
BUF_X4 _11355_ ( .A(_03699_ ), .Z(_03700_ ) );
OAI211_X1 _11356_ ( .A(_03698_ ), .B(fanout_net_39 ), .C1(_03700_ ), .C2(\myreg.Reg[11][17] ), .ZN(_03701_ ) );
NAND3_X1 _11357_ ( .A1(_03697_ ), .A2(_03701_ ), .A3(_03624_ ), .ZN(_03702_ ) );
MUX2_X1 _11358_ ( .A(\myreg.Reg[14][17] ), .B(\myreg.Reg[15][17] ), .S(fanout_net_31 ), .Z(_03703_ ) );
MUX2_X1 _11359_ ( .A(\myreg.Reg[12][17] ), .B(\myreg.Reg[13][17] ), .S(fanout_net_31 ), .Z(_03704_ ) );
BUF_X4 _11360_ ( .A(_03609_ ), .Z(_03705_ ) );
BUF_X4 _11361_ ( .A(_03705_ ), .Z(_03706_ ) );
MUX2_X1 _11362_ ( .A(_03703_ ), .B(_03704_ ), .S(_03706_ ), .Z(_03707_ ) );
BUF_X4 _11363_ ( .A(_03618_ ), .Z(_03708_ ) );
BUF_X4 _11364_ ( .A(_03708_ ), .Z(_03709_ ) );
OAI211_X1 _11365_ ( .A(fanout_net_43 ), .B(_03702_ ), .C1(_03707_ ), .C2(_03709_ ), .ZN(_03710_ ) );
MUX2_X1 _11366_ ( .A(\myreg.Reg[2][17] ), .B(\myreg.Reg[3][17] ), .S(fanout_net_31 ), .Z(_03711_ ) );
AND2_X1 _11367_ ( .A1(_03711_ ), .A2(fanout_net_39 ), .ZN(_03712_ ) );
MUX2_X1 _11368_ ( .A(\myreg.Reg[0][17] ), .B(\myreg.Reg[1][17] ), .S(fanout_net_31 ), .Z(_03713_ ) );
AOI211_X1 _11369_ ( .A(fanout_net_42 ), .B(_03712_ ), .C1(_03670_ ), .C2(_03713_ ), .ZN(_03714_ ) );
MUX2_X1 _11370_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_31 ), .Z(_03715_ ) );
MUX2_X1 _11371_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_31 ), .Z(_03716_ ) );
MUX2_X1 _11372_ ( .A(_03715_ ), .B(_03716_ ), .S(_03706_ ), .Z(_03717_ ) );
OAI21_X1 _11373_ ( .A(_03606_ ), .B1(_03717_ ), .B2(_03624_ ), .ZN(_03718_ ) );
OAI221_X1 _11374_ ( .A(_03710_ ), .B1(_03649_ ), .B2(_03644_ ), .C1(_03714_ ), .C2(_03718_ ), .ZN(_03719_ ) );
OR3_X1 _11375_ ( .A1(_03651_ ), .A2(\EX_LS_result_reg [17] ), .A3(_03653_ ), .ZN(_03720_ ) );
NAND2_X1 _11376_ ( .A1(_03719_ ), .A2(_03720_ ), .ZN(_03721_ ) );
XNOR2_X1 _11377_ ( .A(_03695_ ), .B(_03721_ ), .ZN(_03722_ ) );
OR3_X1 _11378_ ( .A1(_03689_ ), .A2(\EX_LS_result_reg [16] ), .A3(_03690_ ), .ZN(_03723_ ) );
BUF_X4 _11379_ ( .A(_03661_ ), .Z(_03724_ ) );
BUF_X2 _11380_ ( .A(_03613_ ), .Z(_03725_ ) );
OR2_X1 _11381_ ( .A1(_03725_ ), .A2(\myreg.Reg[1][16] ), .ZN(_03726_ ) );
BUF_X4 _11382_ ( .A(_03677_ ), .Z(_03727_ ) );
OAI211_X1 _11383_ ( .A(_03726_ ), .B(_03727_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[0][16] ), .ZN(_03728_ ) );
OR2_X1 _11384_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][16] ), .ZN(_03729_ ) );
OAI211_X1 _11385_ ( .A(_03729_ ), .B(fanout_net_39 ), .C1(_03672_ ), .C2(\myreg.Reg[3][16] ), .ZN(_03730_ ) );
NAND3_X1 _11386_ ( .A1(_03728_ ), .A2(_03667_ ), .A3(_03730_ ), .ZN(_03731_ ) );
MUX2_X1 _11387_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_31 ), .Z(_03732_ ) );
MUX2_X1 _11388_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_31 ), .Z(_03733_ ) );
MUX2_X1 _11389_ ( .A(_03732_ ), .B(_03733_ ), .S(_03670_ ), .Z(_03734_ ) );
OAI211_X1 _11390_ ( .A(_03724_ ), .B(_03731_ ), .C1(_03734_ ), .C2(_03667_ ), .ZN(_03735_ ) );
OR2_X1 _11391_ ( .A1(_03725_ ), .A2(\myreg.Reg[15][16] ), .ZN(_03736_ ) );
OAI211_X1 _11392_ ( .A(_03736_ ), .B(fanout_net_39 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[14][16] ), .ZN(_03737_ ) );
OR2_X1 _11393_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][16] ), .ZN(_03738_ ) );
OAI211_X1 _11394_ ( .A(_03738_ ), .B(_03727_ ), .C1(_03672_ ), .C2(\myreg.Reg[13][16] ), .ZN(_03739_ ) );
NAND3_X1 _11395_ ( .A1(_03737_ ), .A2(fanout_net_42 ), .A3(_03739_ ), .ZN(_03740_ ) );
MUX2_X1 _11396_ ( .A(\myreg.Reg[8][16] ), .B(\myreg.Reg[9][16] ), .S(fanout_net_32 ), .Z(_03741_ ) );
MUX2_X1 _11397_ ( .A(\myreg.Reg[10][16] ), .B(\myreg.Reg[11][16] ), .S(fanout_net_32 ), .Z(_03742_ ) );
MUX2_X1 _11398_ ( .A(_03741_ ), .B(_03742_ ), .S(fanout_net_39 ), .Z(_03743_ ) );
OAI211_X1 _11399_ ( .A(fanout_net_43 ), .B(_03740_ ), .C1(_03743_ ), .C2(fanout_net_42 ), .ZN(_03744_ ) );
OAI211_X1 _11400_ ( .A(_03735_ ), .B(_03744_ ), .C1(_03689_ ), .C2(_03690_ ), .ZN(_03745_ ) );
NAND2_X1 _11401_ ( .A1(_03723_ ), .A2(_03745_ ), .ZN(_03746_ ) );
XOR2_X1 _11402_ ( .A(_03746_ ), .B(_02706_ ), .Z(_03747_ ) );
AND3_X1 _11403_ ( .A1(_03694_ ), .A2(_03722_ ), .A3(_03747_ ), .ZN(_03748_ ) );
OR3_X1 _11404_ ( .A1(_03658_ ), .A2(\EX_LS_result_reg [20] ), .A3(_03659_ ), .ZN(_03749_ ) );
OR2_X1 _11405_ ( .A1(_03725_ ), .A2(\myreg.Reg[1][20] ), .ZN(_03750_ ) );
OAI211_X1 _11406_ ( .A(_03750_ ), .B(_03670_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[0][20] ), .ZN(_03751_ ) );
OR2_X1 _11407_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][20] ), .ZN(_03752_ ) );
OAI211_X1 _11408_ ( .A(_03752_ ), .B(fanout_net_39 ), .C1(_03672_ ), .C2(\myreg.Reg[3][20] ), .ZN(_03753_ ) );
NAND3_X1 _11409_ ( .A1(_03751_ ), .A2(_03667_ ), .A3(_03753_ ), .ZN(_03754_ ) );
MUX2_X1 _11410_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_32 ), .Z(_03755_ ) );
MUX2_X1 _11411_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_32 ), .Z(_03756_ ) );
MUX2_X1 _11412_ ( .A(_03755_ ), .B(_03756_ ), .S(_03670_ ), .Z(_03757_ ) );
OAI211_X1 _11413_ ( .A(_03724_ ), .B(_03754_ ), .C1(_03757_ ), .C2(_03667_ ), .ZN(_03758_ ) );
OR2_X1 _11414_ ( .A1(_03725_ ), .A2(\myreg.Reg[15][20] ), .ZN(_03759_ ) );
OAI211_X1 _11415_ ( .A(_03759_ ), .B(fanout_net_39 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[14][20] ), .ZN(_03760_ ) );
OR2_X1 _11416_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][20] ), .ZN(_03761_ ) );
OAI211_X1 _11417_ ( .A(_03761_ ), .B(_03670_ ), .C1(_03672_ ), .C2(\myreg.Reg[13][20] ), .ZN(_03762_ ) );
NAND3_X1 _11418_ ( .A1(_03760_ ), .A2(fanout_net_42 ), .A3(_03762_ ), .ZN(_03763_ ) );
MUX2_X1 _11419_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_32 ), .Z(_03764_ ) );
MUX2_X1 _11420_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_32 ), .Z(_03765_ ) );
MUX2_X1 _11421_ ( .A(_03764_ ), .B(_03765_ ), .S(fanout_net_39 ), .Z(_03766_ ) );
OAI211_X1 _11422_ ( .A(fanout_net_43 ), .B(_03763_ ), .C1(_03766_ ), .C2(fanout_net_42 ), .ZN(_03767_ ) );
OAI211_X1 _11423_ ( .A(_03758_ ), .B(_03767_ ), .C1(_03689_ ), .C2(_03690_ ), .ZN(_03768_ ) );
NAND2_X1 _11424_ ( .A1(_03749_ ), .A2(_03768_ ), .ZN(_03769_ ) );
XOR2_X1 _11425_ ( .A(_03769_ ), .B(_02598_ ), .Z(_03770_ ) );
OR3_X1 _11426_ ( .A1(_03658_ ), .A2(\EX_LS_result_reg [21] ), .A3(_03659_ ), .ZN(_03771_ ) );
OR2_X1 _11427_ ( .A1(\myreg.Reg[0][21] ), .A2(fanout_net_32 ), .ZN(_03772_ ) );
OAI211_X1 _11428_ ( .A(_03772_ ), .B(_03670_ ), .C1(\myreg.Reg[1][21] ), .C2(_03725_ ), .ZN(_03773_ ) );
OR2_X1 _11429_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][21] ), .ZN(_03774_ ) );
OAI211_X1 _11430_ ( .A(_03774_ ), .B(fanout_net_39 ), .C1(_03672_ ), .C2(\myreg.Reg[3][21] ), .ZN(_03775_ ) );
NAND3_X1 _11431_ ( .A1(_03773_ ), .A2(_03775_ ), .A3(_03709_ ), .ZN(_03776_ ) );
MUX2_X1 _11432_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_32 ), .Z(_03777_ ) );
MUX2_X1 _11433_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_32 ), .Z(_03778_ ) );
MUX2_X1 _11434_ ( .A(_03777_ ), .B(_03778_ ), .S(_03677_ ), .Z(_03779_ ) );
OAI211_X1 _11435_ ( .A(_03661_ ), .B(_03776_ ), .C1(_03779_ ), .C2(_03667_ ), .ZN(_03780_ ) );
OR2_X1 _11436_ ( .A1(_03664_ ), .A2(\myreg.Reg[13][21] ), .ZN(_03781_ ) );
OAI211_X1 _11437_ ( .A(_03781_ ), .B(_03670_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[12][21] ), .ZN(_03782_ ) );
OR2_X1 _11438_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[14][21] ), .ZN(_03783_ ) );
OAI211_X1 _11439_ ( .A(_03783_ ), .B(fanout_net_39 ), .C1(_03725_ ), .C2(\myreg.Reg[15][21] ), .ZN(_03784_ ) );
NAND3_X1 _11440_ ( .A1(_03782_ ), .A2(fanout_net_42 ), .A3(_03784_ ), .ZN(_03785_ ) );
MUX2_X1 _11441_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_32 ), .Z(_03786_ ) );
MUX2_X1 _11442_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_32 ), .Z(_03787_ ) );
MUX2_X1 _11443_ ( .A(_03786_ ), .B(_03787_ ), .S(fanout_net_39 ), .Z(_03788_ ) );
OAI211_X1 _11444_ ( .A(fanout_net_43 ), .B(_03785_ ), .C1(_03788_ ), .C2(fanout_net_42 ), .ZN(_03789_ ) );
OAI211_X1 _11445_ ( .A(_03780_ ), .B(_03789_ ), .C1(_03658_ ), .C2(_03659_ ), .ZN(_03790_ ) );
NAND2_X1 _11446_ ( .A1(_03771_ ), .A2(_03790_ ), .ZN(_03791_ ) );
AND2_X1 _11447_ ( .A1(_03791_ ), .A2(_02574_ ), .ZN(_03792_ ) );
NOR2_X1 _11448_ ( .A1(_03791_ ), .A2(_02575_ ), .ZN(_03793_ ) );
NOR2_X1 _11449_ ( .A1(_03792_ ), .A2(_03793_ ), .ZN(_03794_ ) );
AND2_X1 _11450_ ( .A1(_03770_ ), .A2(_03794_ ), .ZN(_03795_ ) );
OR3_X1 _11451_ ( .A1(_03658_ ), .A2(\EX_LS_result_reg [23] ), .A3(_03644_ ), .ZN(_03796_ ) );
OR2_X1 _11452_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[4][23] ), .ZN(_03797_ ) );
OAI211_X1 _11453_ ( .A(_03797_ ), .B(_03677_ ), .C1(_03725_ ), .C2(\myreg.Reg[5][23] ), .ZN(_03798_ ) );
OR2_X1 _11454_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[6][23] ), .ZN(_03799_ ) );
OAI211_X1 _11455_ ( .A(_03799_ ), .B(fanout_net_39 ), .C1(_03725_ ), .C2(\myreg.Reg[7][23] ), .ZN(_03800_ ) );
NAND3_X1 _11456_ ( .A1(_03798_ ), .A2(_03800_ ), .A3(fanout_net_42 ), .ZN(_03801_ ) );
MUX2_X1 _11457_ ( .A(\myreg.Reg[2][23] ), .B(\myreg.Reg[3][23] ), .S(fanout_net_32 ), .Z(_03802_ ) );
MUX2_X1 _11458_ ( .A(\myreg.Reg[0][23] ), .B(\myreg.Reg[1][23] ), .S(fanout_net_32 ), .Z(_03803_ ) );
MUX2_X1 _11459_ ( .A(_03802_ ), .B(_03803_ ), .S(_03677_ ), .Z(_03804_ ) );
OAI211_X1 _11460_ ( .A(_03661_ ), .B(_03801_ ), .C1(_03804_ ), .C2(fanout_net_42 ), .ZN(_03805_ ) );
NOR2_X1 _11461_ ( .A1(_03671_ ), .A2(\myreg.Reg[11][23] ), .ZN(_03806_ ) );
OAI21_X1 _11462_ ( .A(fanout_net_39 ), .B1(fanout_net_32 ), .B2(\myreg.Reg[10][23] ), .ZN(_03807_ ) );
NOR2_X1 _11463_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][23] ), .ZN(_03808_ ) );
OAI21_X1 _11464_ ( .A(_03677_ ), .B1(_03671_ ), .B2(\myreg.Reg[9][23] ), .ZN(_03809_ ) );
OAI221_X1 _11465_ ( .A(_03709_ ), .B1(_03806_ ), .B2(_03807_ ), .C1(_03808_ ), .C2(_03809_ ), .ZN(_03810_ ) );
MUX2_X1 _11466_ ( .A(\myreg.Reg[12][23] ), .B(\myreg.Reg[13][23] ), .S(fanout_net_32 ), .Z(_03811_ ) );
MUX2_X1 _11467_ ( .A(\myreg.Reg[14][23] ), .B(\myreg.Reg[15][23] ), .S(fanout_net_32 ), .Z(_03812_ ) );
MUX2_X1 _11468_ ( .A(_03811_ ), .B(_03812_ ), .S(fanout_net_39 ), .Z(_03813_ ) );
OAI211_X1 _11469_ ( .A(fanout_net_43 ), .B(_03810_ ), .C1(_03813_ ), .C2(_03709_ ), .ZN(_03814_ ) );
OAI211_X1 _11470_ ( .A(_03805_ ), .B(_03814_ ), .C1(_03658_ ), .C2(_03659_ ), .ZN(_03815_ ) );
NAND2_X1 _11471_ ( .A1(_03796_ ), .A2(_03815_ ), .ZN(_03816_ ) );
XOR2_X1 _11472_ ( .A(_02548_ ), .B(_03816_ ), .Z(_03817_ ) );
OR3_X1 _11473_ ( .A1(_03658_ ), .A2(\EX_LS_result_reg [22] ), .A3(_03659_ ), .ZN(_03818_ ) );
OR2_X1 _11474_ ( .A1(_03671_ ), .A2(\myreg.Reg[7][22] ), .ZN(_03819_ ) );
OAI211_X1 _11475_ ( .A(_03819_ ), .B(fanout_net_39 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[6][22] ), .ZN(_03820_ ) );
OR2_X1 _11476_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[4][22] ), .ZN(_03821_ ) );
OAI211_X1 _11477_ ( .A(_03821_ ), .B(_03670_ ), .C1(_03672_ ), .C2(\myreg.Reg[5][22] ), .ZN(_03822_ ) );
NAND3_X1 _11478_ ( .A1(_03820_ ), .A2(fanout_net_42 ), .A3(_03822_ ), .ZN(_03823_ ) );
MUX2_X1 _11479_ ( .A(\myreg.Reg[2][22] ), .B(\myreg.Reg[3][22] ), .S(fanout_net_32 ), .Z(_03824_ ) );
MUX2_X1 _11480_ ( .A(\myreg.Reg[0][22] ), .B(\myreg.Reg[1][22] ), .S(fanout_net_33 ), .Z(_03825_ ) );
MUX2_X1 _11481_ ( .A(_03824_ ), .B(_03825_ ), .S(_03677_ ), .Z(_03826_ ) );
OAI211_X1 _11482_ ( .A(_03661_ ), .B(_03823_ ), .C1(_03826_ ), .C2(fanout_net_42 ), .ZN(_03827_ ) );
NOR2_X1 _11483_ ( .A1(_03725_ ), .A2(\myreg.Reg[11][22] ), .ZN(_03828_ ) );
OAI21_X1 _11484_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myreg.Reg[10][22] ), .ZN(_03829_ ) );
NOR2_X1 _11485_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[8][22] ), .ZN(_03830_ ) );
OAI21_X1 _11486_ ( .A(_03677_ ), .B1(_03725_ ), .B2(\myreg.Reg[9][22] ), .ZN(_03831_ ) );
OAI221_X1 _11487_ ( .A(_03709_ ), .B1(_03828_ ), .B2(_03829_ ), .C1(_03830_ ), .C2(_03831_ ), .ZN(_03832_ ) );
MUX2_X1 _11488_ ( .A(\myreg.Reg[12][22] ), .B(\myreg.Reg[13][22] ), .S(fanout_net_33 ), .Z(_03833_ ) );
MUX2_X1 _11489_ ( .A(\myreg.Reg[14][22] ), .B(\myreg.Reg[15][22] ), .S(fanout_net_33 ), .Z(_03834_ ) );
MUX2_X1 _11490_ ( .A(_03833_ ), .B(_03834_ ), .S(fanout_net_39 ), .Z(_03835_ ) );
OAI211_X1 _11491_ ( .A(fanout_net_43 ), .B(_03832_ ), .C1(_03835_ ), .C2(_03667_ ), .ZN(_03836_ ) );
OAI211_X1 _11492_ ( .A(_03827_ ), .B(_03836_ ), .C1(_03689_ ), .C2(_03690_ ), .ZN(_03837_ ) );
NAND2_X1 _11493_ ( .A1(_03818_ ), .A2(_03837_ ), .ZN(_03838_ ) );
XOR2_X1 _11494_ ( .A(_02521_ ), .B(_03838_ ), .Z(_03839_ ) );
AND3_X1 _11495_ ( .A1(_03795_ ), .A2(_03817_ ), .A3(_03839_ ), .ZN(_03840_ ) );
AND2_X1 _11496_ ( .A1(_03748_ ), .A2(_03840_ ), .ZN(_03841_ ) );
BUF_X2 _11497_ ( .A(_03689_ ), .Z(_03842_ ) );
BUF_X2 _11498_ ( .A(_03690_ ), .Z(_03843_ ) );
OR3_X1 _11499_ ( .A1(_03842_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_03843_ ), .ZN(_03844_ ) );
OR2_X1 _11500_ ( .A1(fanout_net_33 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03845_ ) );
BUF_X4 _11501_ ( .A(_03727_ ), .Z(_03846_ ) );
BUF_X2 _11502_ ( .A(_03672_ ), .Z(_03847_ ) );
BUF_X4 _11503_ ( .A(_03847_ ), .Z(_03848_ ) );
OAI211_X1 _11504_ ( .A(_03845_ ), .B(_03846_ ), .C1(_03848_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03849_ ) );
OR2_X1 _11505_ ( .A1(fanout_net_33 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03850_ ) );
OAI211_X1 _11506_ ( .A(_03850_ ), .B(fanout_net_39 ), .C1(_03848_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03851_ ) );
BUF_X4 _11507_ ( .A(_03667_ ), .Z(_03852_ ) );
NAND3_X1 _11508_ ( .A1(_03849_ ), .A2(_03851_ ), .A3(_03852_ ), .ZN(_03853_ ) );
MUX2_X1 _11509_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03854_ ) );
MUX2_X1 _11510_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03855_ ) );
MUX2_X1 _11511_ ( .A(_03854_ ), .B(_03855_ ), .S(_03846_ ), .Z(_03856_ ) );
BUF_X4 _11512_ ( .A(_03852_ ), .Z(_03857_ ) );
OAI211_X1 _11513_ ( .A(_03724_ ), .B(_03853_ ), .C1(_03856_ ), .C2(_03857_ ), .ZN(_03858_ ) );
OR2_X1 _11514_ ( .A1(fanout_net_33 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03859_ ) );
OAI211_X1 _11515_ ( .A(_03859_ ), .B(fanout_net_39 ), .C1(_03848_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03860_ ) );
NAND2_X1 _11516_ ( .A1(_03245_ ), .A2(fanout_net_33 ), .ZN(_03861_ ) );
OAI211_X1 _11517_ ( .A(_03861_ ), .B(_03846_ ), .C1(fanout_net_33 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03862_ ) );
NAND3_X1 _11518_ ( .A1(_03860_ ), .A2(_03862_ ), .A3(fanout_net_42 ), .ZN(_03863_ ) );
MUX2_X1 _11519_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03864_ ) );
MUX2_X1 _11520_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03865_ ) );
MUX2_X1 _11521_ ( .A(_03864_ ), .B(_03865_ ), .S(fanout_net_39 ), .Z(_03866_ ) );
OAI211_X1 _11522_ ( .A(fanout_net_43 ), .B(_03863_ ), .C1(_03866_ ), .C2(fanout_net_42 ), .ZN(_03867_ ) );
OAI211_X1 _11523_ ( .A(_03858_ ), .B(_03867_ ), .C1(_03842_ ), .C2(_03843_ ), .ZN(_03868_ ) );
NAND2_X1 _11524_ ( .A1(_03844_ ), .A2(_03868_ ), .ZN(_03869_ ) );
XNOR2_X1 _11525_ ( .A(_03253_ ), .B(_03869_ ), .ZN(_03870_ ) );
OR3_X1 _11526_ ( .A1(_03689_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03690_ ), .ZN(_03871_ ) );
OR2_X1 _11527_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03872_ ) );
OAI211_X1 _11528_ ( .A(_03872_ ), .B(_03727_ ), .C1(_03847_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03873_ ) );
OR2_X1 _11529_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03874_ ) );
OAI211_X1 _11530_ ( .A(_03874_ ), .B(fanout_net_39 ), .C1(_03847_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03875_ ) );
NAND3_X1 _11531_ ( .A1(_03873_ ), .A2(_03875_ ), .A3(fanout_net_42 ), .ZN(_03876_ ) );
MUX2_X1 _11532_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03877_ ) );
MUX2_X1 _11533_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03878_ ) );
MUX2_X1 _11534_ ( .A(_03877_ ), .B(_03878_ ), .S(_03727_ ), .Z(_03879_ ) );
OAI211_X1 _11535_ ( .A(_03724_ ), .B(_03876_ ), .C1(_03879_ ), .C2(fanout_net_42 ), .ZN(_03880_ ) );
NOR2_X1 _11536_ ( .A1(_03847_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03881_ ) );
OAI21_X1 _11537_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03882_ ) );
NOR2_X1 _11538_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03883_ ) );
OAI21_X1 _11539_ ( .A(_03727_ ), .B1(_03847_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03884_ ) );
OAI221_X1 _11540_ ( .A(_03667_ ), .B1(_03881_ ), .B2(_03882_ ), .C1(_03883_ ), .C2(_03884_ ), .ZN(_03885_ ) );
MUX2_X1 _11541_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03886_ ) );
MUX2_X1 _11542_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03887_ ) );
MUX2_X1 _11543_ ( .A(_03886_ ), .B(_03887_ ), .S(fanout_net_39 ), .Z(_03888_ ) );
OAI211_X1 _11544_ ( .A(fanout_net_43 ), .B(_03885_ ), .C1(_03888_ ), .C2(_03852_ ), .ZN(_03889_ ) );
OAI211_X1 _11545_ ( .A(_03880_ ), .B(_03889_ ), .C1(_03689_ ), .C2(_03690_ ), .ZN(_03890_ ) );
NAND2_X1 _11546_ ( .A1(_03871_ ), .A2(_03890_ ), .ZN(_03891_ ) );
XNOR2_X1 _11547_ ( .A(_03276_ ), .B(_03891_ ), .ZN(_03892_ ) );
AND2_X1 _11548_ ( .A1(_03870_ ), .A2(_03892_ ), .ZN(_03893_ ) );
OR3_X1 _11549_ ( .A1(_03689_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03690_ ), .ZN(_03894_ ) );
OR2_X1 _11550_ ( .A1(_03847_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03895_ ) );
OAI211_X1 _11551_ ( .A(_03895_ ), .B(fanout_net_40 ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03896_ ) );
OR2_X1 _11552_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03897_ ) );
BUF_X4 _11553_ ( .A(_03727_ ), .Z(_03898_ ) );
BUF_X4 _11554_ ( .A(_03672_ ), .Z(_03899_ ) );
OAI211_X1 _11555_ ( .A(_03897_ ), .B(_03898_ ), .C1(_03899_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03900_ ) );
NAND3_X1 _11556_ ( .A1(_03896_ ), .A2(_03852_ ), .A3(_03900_ ), .ZN(_03901_ ) );
MUX2_X1 _11557_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03902_ ) );
MUX2_X1 _11558_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03903_ ) );
MUX2_X1 _11559_ ( .A(_03902_ ), .B(_03903_ ), .S(_03727_ ), .Z(_03904_ ) );
OAI211_X1 _11560_ ( .A(_03724_ ), .B(_03901_ ), .C1(_03904_ ), .C2(_03857_ ), .ZN(_03905_ ) );
OR2_X1 _11561_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03906_ ) );
OAI211_X1 _11562_ ( .A(_03906_ ), .B(fanout_net_40 ), .C1(_03899_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03907_ ) );
OR2_X1 _11563_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03908_ ) );
OAI211_X1 _11564_ ( .A(_03908_ ), .B(_03898_ ), .C1(_03899_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03909_ ) );
NAND3_X1 _11565_ ( .A1(_03907_ ), .A2(_03909_ ), .A3(fanout_net_42 ), .ZN(_03910_ ) );
MUX2_X1 _11566_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03911_ ) );
MUX2_X1 _11567_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03912_ ) );
MUX2_X1 _11568_ ( .A(_03911_ ), .B(_03912_ ), .S(fanout_net_40 ), .Z(_03913_ ) );
OAI211_X1 _11569_ ( .A(fanout_net_43 ), .B(_03910_ ), .C1(_03913_ ), .C2(fanout_net_42 ), .ZN(_03914_ ) );
OAI211_X1 _11570_ ( .A(_03905_ ), .B(_03914_ ), .C1(_03842_ ), .C2(_03843_ ), .ZN(_03915_ ) );
NAND2_X1 _11571_ ( .A1(_03894_ ), .A2(_03915_ ), .ZN(_03916_ ) );
XNOR2_X1 _11572_ ( .A(_03916_ ), .B(_03336_ ), .ZN(_03917_ ) );
OR3_X1 _11573_ ( .A1(_03842_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_03843_ ), .ZN(_03918_ ) );
OR2_X1 _11574_ ( .A1(_03847_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03919_ ) );
OAI211_X1 _11575_ ( .A(_03919_ ), .B(fanout_net_40 ), .C1(fanout_net_34 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03920_ ) );
OR2_X1 _11576_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03921_ ) );
OAI211_X1 _11577_ ( .A(_03921_ ), .B(_03846_ ), .C1(_03848_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03922_ ) );
NAND3_X1 _11578_ ( .A1(_03920_ ), .A2(fanout_net_42 ), .A3(_03922_ ), .ZN(_03923_ ) );
MUX2_X1 _11579_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03924_ ) );
MUX2_X1 _11580_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03925_ ) );
MUX2_X1 _11581_ ( .A(_03924_ ), .B(_03925_ ), .S(_03846_ ), .Z(_03926_ ) );
OAI211_X1 _11582_ ( .A(_03724_ ), .B(_03923_ ), .C1(_03926_ ), .C2(fanout_net_42 ), .ZN(_03927_ ) );
NOR2_X1 _11583_ ( .A1(_03899_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03928_ ) );
OAI21_X1 _11584_ ( .A(fanout_net_40 ), .B1(fanout_net_34 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03929_ ) );
MUX2_X1 _11585_ ( .A(_03296_ ), .B(_03297_ ), .S(fanout_net_34 ), .Z(_03930_ ) );
OAI221_X1 _11586_ ( .A(_03852_ ), .B1(_03928_ ), .B2(_03929_ ), .C1(_03930_ ), .C2(fanout_net_40 ), .ZN(_03931_ ) );
MUX2_X1 _11587_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03932_ ) );
MUX2_X1 _11588_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03933_ ) );
MUX2_X1 _11589_ ( .A(_03932_ ), .B(_03933_ ), .S(fanout_net_40 ), .Z(_03934_ ) );
OAI211_X1 _11590_ ( .A(fanout_net_43 ), .B(_03931_ ), .C1(_03934_ ), .C2(_03857_ ), .ZN(_03935_ ) );
OAI211_X1 _11591_ ( .A(_03927_ ), .B(_03935_ ), .C1(_03842_ ), .C2(_03843_ ), .ZN(_03936_ ) );
NAND2_X1 _11592_ ( .A1(_03918_ ), .A2(_03936_ ), .ZN(_03937_ ) );
INV_X1 _11593_ ( .A(_03937_ ), .ZN(_03938_ ) );
XNOR2_X1 _11594_ ( .A(_03309_ ), .B(_03938_ ), .ZN(_03939_ ) );
AND3_X1 _11595_ ( .A1(_03893_ ), .A2(_03917_ ), .A3(_03939_ ), .ZN(_03940_ ) );
NOR2_X2 _11596_ ( .A1(_03647_ ), .A2(_03642_ ), .ZN(_03941_ ) );
NAND2_X1 _11597_ ( .A1(_03941_ ), .A2(\EX_LS_result_reg [24] ), .ZN(_03942_ ) );
OR2_X1 _11598_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03943_ ) );
OAI211_X1 _11599_ ( .A(_03943_ ), .B(_03846_ ), .C1(_03848_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03944_ ) );
OR2_X1 _11600_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03945_ ) );
OAI211_X1 _11601_ ( .A(_03945_ ), .B(fanout_net_40 ), .C1(_03848_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03946_ ) );
NAND3_X1 _11602_ ( .A1(_03944_ ), .A2(_03946_ ), .A3(fanout_net_42 ), .ZN(_03947_ ) );
MUX2_X1 _11603_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03948_ ) );
MUX2_X1 _11604_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03949_ ) );
MUX2_X1 _11605_ ( .A(_03948_ ), .B(_03949_ ), .S(_03846_ ), .Z(_03950_ ) );
OAI211_X1 _11606_ ( .A(_03724_ ), .B(_03947_ ), .C1(_03950_ ), .C2(fanout_net_42 ), .ZN(_03951_ ) );
NOR2_X1 _11607_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03952_ ) );
OAI21_X1 _11608_ ( .A(_03846_ ), .B1(_03848_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03953_ ) );
MUX2_X1 _11609_ ( .A(_03161_ ), .B(_03162_ ), .S(fanout_net_34 ), .Z(_03954_ ) );
OAI221_X1 _11610_ ( .A(_03857_ ), .B1(_03952_ ), .B2(_03953_ ), .C1(_03954_ ), .C2(_03846_ ), .ZN(_03955_ ) );
MUX2_X1 _11611_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03956_ ) );
MUX2_X1 _11612_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03957_ ) );
MUX2_X1 _11613_ ( .A(_03956_ ), .B(_03957_ ), .S(fanout_net_40 ), .Z(_03958_ ) );
OAI211_X1 _11614_ ( .A(fanout_net_43 ), .B(_03955_ ), .C1(_03958_ ), .C2(_03857_ ), .ZN(_03959_ ) );
OAI211_X1 _11615_ ( .A(_03951_ ), .B(_03959_ ), .C1(_03842_ ), .C2(_03843_ ), .ZN(_03960_ ) );
NAND2_X1 _11616_ ( .A1(_03942_ ), .A2(_03960_ ), .ZN(_03961_ ) );
XNOR2_X1 _11617_ ( .A(_03961_ ), .B(_03172_ ), .ZN(_03962_ ) );
INV_X1 _11618_ ( .A(\EX_LS_result_reg [25] ), .ZN(_03963_ ) );
OR3_X1 _11619_ ( .A1(_03689_ ), .A2(_03963_ ), .A3(_03690_ ), .ZN(_03964_ ) );
OR2_X1 _11620_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03965_ ) );
OAI211_X1 _11621_ ( .A(_03965_ ), .B(_03898_ ), .C1(_03899_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03966_ ) );
OR2_X1 _11622_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03967_ ) );
OAI211_X1 _11623_ ( .A(_03967_ ), .B(fanout_net_40 ), .C1(_03899_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03968_ ) );
NAND3_X1 _11624_ ( .A1(_03966_ ), .A2(_03968_ ), .A3(_03852_ ), .ZN(_03969_ ) );
MUX2_X1 _11625_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03970_ ) );
MUX2_X1 _11626_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03971_ ) );
MUX2_X1 _11627_ ( .A(_03970_ ), .B(_03971_ ), .S(_03898_ ), .Z(_03972_ ) );
OAI211_X1 _11628_ ( .A(fanout_net_43 ), .B(_03969_ ), .C1(_03972_ ), .C2(_03857_ ), .ZN(_03973_ ) );
NOR2_X1 _11629_ ( .A1(_03899_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03974_ ) );
OAI21_X1 _11630_ ( .A(fanout_net_40 ), .B1(fanout_net_34 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03975_ ) );
NOR2_X1 _11631_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03976_ ) );
OAI21_X1 _11632_ ( .A(_03898_ ), .B1(_03899_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03977_ ) );
OAI221_X1 _11633_ ( .A(_03852_ ), .B1(_03974_ ), .B2(_03975_ ), .C1(_03976_ ), .C2(_03977_ ), .ZN(_03978_ ) );
MUX2_X1 _11634_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03979_ ) );
MUX2_X1 _11635_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03980_ ) );
MUX2_X1 _11636_ ( .A(_03979_ ), .B(_03980_ ), .S(_03898_ ), .Z(_03981_ ) );
OAI211_X1 _11637_ ( .A(_03724_ ), .B(_03978_ ), .C1(_03981_ ), .C2(_03857_ ), .ZN(_03982_ ) );
OAI211_X1 _11638_ ( .A(_03973_ ), .B(_03982_ ), .C1(_03842_ ), .C2(_03843_ ), .ZN(_03983_ ) );
NAND2_X1 _11639_ ( .A1(_03964_ ), .A2(_03983_ ), .ZN(_03984_ ) );
XNOR2_X1 _11640_ ( .A(_03198_ ), .B(_03984_ ), .ZN(_03985_ ) );
AND2_X1 _11641_ ( .A1(_03962_ ), .A2(_03985_ ), .ZN(_03986_ ) );
NAND2_X1 _11642_ ( .A1(_02483_ ), .A2(_02493_ ), .ZN(_03987_ ) );
INV_X1 _11643_ ( .A(\EX_LS_result_reg [27] ), .ZN(_03988_ ) );
OR3_X1 _11644_ ( .A1(_03842_ ), .A2(_03988_ ), .A3(_03843_ ), .ZN(_03989_ ) );
OR2_X1 _11645_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03990_ ) );
OAI211_X1 _11646_ ( .A(_03990_ ), .B(_03846_ ), .C1(_03848_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03991_ ) );
OR2_X1 _11647_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03992_ ) );
OAI211_X1 _11648_ ( .A(_03992_ ), .B(fanout_net_40 ), .C1(_03848_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03993_ ) );
NAND3_X1 _11649_ ( .A1(_03991_ ), .A2(_03993_ ), .A3(_03852_ ), .ZN(_03994_ ) );
MUX2_X1 _11650_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03995_ ) );
MUX2_X1 _11651_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03996_ ) );
MUX2_X1 _11652_ ( .A(_03995_ ), .B(_03996_ ), .S(_03898_ ), .Z(_03997_ ) );
OAI211_X1 _11653_ ( .A(fanout_net_43 ), .B(_03994_ ), .C1(_03997_ ), .C2(_03857_ ), .ZN(_03998_ ) );
OR2_X1 _11654_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03999_ ) );
OAI211_X1 _11655_ ( .A(_03999_ ), .B(_03898_ ), .C1(_03848_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04000_ ) );
OR2_X1 _11656_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04001_ ) );
OAI211_X1 _11657_ ( .A(_04001_ ), .B(fanout_net_40 ), .C1(_03899_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04002_ ) );
NAND3_X1 _11658_ ( .A1(_04000_ ), .A2(_04002_ ), .A3(_03852_ ), .ZN(_04003_ ) );
MUX2_X1 _11659_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04004_ ) );
MUX2_X1 _11660_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04005_ ) );
MUX2_X1 _11661_ ( .A(_04004_ ), .B(_04005_ ), .S(_03898_ ), .Z(_04006_ ) );
OAI211_X1 _11662_ ( .A(_03724_ ), .B(_04003_ ), .C1(_04006_ ), .C2(_03857_ ), .ZN(_04007_ ) );
OAI211_X1 _11663_ ( .A(_03998_ ), .B(_04007_ ), .C1(_03842_ ), .C2(_03843_ ), .ZN(_04008_ ) );
NAND2_X1 _11664_ ( .A1(_03989_ ), .A2(_04008_ ), .ZN(_04009_ ) );
XNOR2_X1 _11665_ ( .A(_03987_ ), .B(_04009_ ), .ZN(_04010_ ) );
NAND2_X1 _11666_ ( .A1(_03941_ ), .A2(\EX_LS_result_reg [26] ), .ZN(_04011_ ) );
OR2_X1 _11667_ ( .A1(_03847_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04012_ ) );
OAI211_X1 _11668_ ( .A(_04012_ ), .B(_03898_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04013_ ) );
OR2_X1 _11669_ ( .A1(_03847_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04014_ ) );
OAI211_X1 _11670_ ( .A(_04014_ ), .B(fanout_net_40 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04015_ ) );
NAND3_X1 _11671_ ( .A1(_04013_ ), .A2(_04015_ ), .A3(fanout_net_42 ), .ZN(_04016_ ) );
MUX2_X1 _11672_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04017_ ) );
MUX2_X1 _11673_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04018_ ) );
MUX2_X1 _11674_ ( .A(_04017_ ), .B(_04018_ ), .S(_03727_ ), .Z(_04019_ ) );
OAI211_X1 _11675_ ( .A(_03724_ ), .B(_04016_ ), .C1(_04019_ ), .C2(fanout_net_42 ), .ZN(_04020_ ) );
NOR2_X1 _11676_ ( .A1(_03847_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04021_ ) );
OAI21_X1 _11677_ ( .A(fanout_net_40 ), .B1(fanout_net_35 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04022_ ) );
NOR2_X1 _11678_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04023_ ) );
OAI21_X1 _11679_ ( .A(_03727_ ), .B1(_03899_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04024_ ) );
OAI221_X1 _11680_ ( .A(_03852_ ), .B1(_04021_ ), .B2(_04022_ ), .C1(_04023_ ), .C2(_04024_ ), .ZN(_04025_ ) );
MUX2_X1 _11681_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04026_ ) );
MUX2_X1 _11682_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04027_ ) );
MUX2_X1 _11683_ ( .A(_04026_ ), .B(_04027_ ), .S(fanout_net_40 ), .Z(_04028_ ) );
OAI211_X1 _11684_ ( .A(fanout_net_43 ), .B(_04025_ ), .C1(_04028_ ), .C2(_03857_ ), .ZN(_04029_ ) );
OAI211_X1 _11685_ ( .A(_04020_ ), .B(_04029_ ), .C1(_03842_ ), .C2(_03843_ ), .ZN(_04030_ ) );
NAND2_X1 _11686_ ( .A1(_04011_ ), .A2(_04030_ ), .ZN(_04031_ ) );
XNOR2_X1 _11687_ ( .A(_04031_ ), .B(_03221_ ), .ZN(_04032_ ) );
AND3_X1 _11688_ ( .A1(_03986_ ), .A2(_04010_ ), .A3(_04032_ ), .ZN(_04033_ ) );
AND3_X1 _11689_ ( .A1(_03841_ ), .A2(_03940_ ), .A3(_04033_ ), .ZN(_04034_ ) );
OR3_X4 _11690_ ( .A1(_03648_ ), .A2(\EX_LS_result_reg [1] ), .A3(_03643_ ), .ZN(_04035_ ) );
OR2_X1 _11691_ ( .A1(_03662_ ), .A2(\myreg.Reg[7][1] ), .ZN(_04036_ ) );
OAI211_X1 _11692_ ( .A(_04036_ ), .B(fanout_net_40 ), .C1(fanout_net_35 ), .C2(\myreg.Reg[6][1] ), .ZN(_04037_ ) );
OR2_X1 _11693_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[4][1] ), .ZN(_04038_ ) );
OAI211_X1 _11694_ ( .A(_04038_ ), .B(_03705_ ), .C1(_03699_ ), .C2(\myreg.Reg[5][1] ), .ZN(_04039_ ) );
NAND3_X1 _11695_ ( .A1(_04037_ ), .A2(fanout_net_42 ), .A3(_04039_ ), .ZN(_04040_ ) );
MUX2_X1 _11696_ ( .A(\myreg.Reg[2][1] ), .B(\myreg.Reg[3][1] ), .S(fanout_net_35 ), .Z(_04041_ ) );
MUX2_X1 _11697_ ( .A(\myreg.Reg[0][1] ), .B(\myreg.Reg[1][1] ), .S(fanout_net_35 ), .Z(_04042_ ) );
BUF_X4 _11698_ ( .A(_03608_ ), .Z(_04043_ ) );
MUX2_X1 _11699_ ( .A(_04041_ ), .B(_04042_ ), .S(_04043_ ), .Z(_04044_ ) );
OAI211_X1 _11700_ ( .A(_03606_ ), .B(_04040_ ), .C1(_04044_ ), .C2(fanout_net_42 ), .ZN(_04045_ ) );
NOR2_X1 _11701_ ( .A1(_03699_ ), .A2(\myreg.Reg[11][1] ), .ZN(_04046_ ) );
OAI21_X1 _11702_ ( .A(fanout_net_40 ), .B1(fanout_net_35 ), .B2(\myreg.Reg[10][1] ), .ZN(_04047_ ) );
NOR2_X1 _11703_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[8][1] ), .ZN(_04048_ ) );
OAI21_X1 _11704_ ( .A(_04043_ ), .B1(_03699_ ), .B2(\myreg.Reg[9][1] ), .ZN(_04049_ ) );
OAI221_X1 _11705_ ( .A(_03618_ ), .B1(_04046_ ), .B2(_04047_ ), .C1(_04048_ ), .C2(_04049_ ), .ZN(_04050_ ) );
MUX2_X1 _11706_ ( .A(\myreg.Reg[12][1] ), .B(\myreg.Reg[13][1] ), .S(fanout_net_35 ), .Z(_04051_ ) );
MUX2_X1 _11707_ ( .A(\myreg.Reg[14][1] ), .B(\myreg.Reg[15][1] ), .S(fanout_net_35 ), .Z(_04052_ ) );
MUX2_X1 _11708_ ( .A(_04051_ ), .B(_04052_ ), .S(fanout_net_40 ), .Z(_04053_ ) );
OAI211_X1 _11709_ ( .A(fanout_net_43 ), .B(_04050_ ), .C1(_04053_ ), .C2(_03619_ ), .ZN(_04054_ ) );
OAI211_X1 _11710_ ( .A(_04045_ ), .B(_04054_ ), .C1(_03651_ ), .C2(_03653_ ), .ZN(_04055_ ) );
NAND2_X1 _11711_ ( .A1(_04035_ ), .A2(_04055_ ), .ZN(_04056_ ) );
XOR2_X1 _11712_ ( .A(_04056_ ), .B(_02779_ ), .Z(_04057_ ) );
NAND2_X2 _11713_ ( .A1(_02783_ ), .A2(_02802_ ), .ZN(_04058_ ) );
OR2_X1 _11714_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][0] ), .ZN(_04059_ ) );
OAI211_X1 _11715_ ( .A(_04059_ ), .B(_04043_ ), .C1(_03612_ ), .C2(\myreg.Reg[1][0] ), .ZN(_04060_ ) );
OR2_X1 _11716_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][0] ), .ZN(_04061_ ) );
OAI211_X1 _11717_ ( .A(_04061_ ), .B(fanout_net_40 ), .C1(_03612_ ), .C2(\myreg.Reg[3][0] ), .ZN(_04062_ ) );
NAND3_X1 _11718_ ( .A1(_04060_ ), .A2(_04062_ ), .A3(_03618_ ), .ZN(_04063_ ) );
MUX2_X1 _11719_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_35 ), .Z(_04064_ ) );
MUX2_X1 _11720_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_35 ), .Z(_04065_ ) );
MUX2_X1 _11721_ ( .A(_04064_ ), .B(_04065_ ), .S(_04043_ ), .Z(_04066_ ) );
OAI211_X1 _11722_ ( .A(_03605_ ), .B(_04063_ ), .C1(_04066_ ), .C2(_03619_ ), .ZN(_04067_ ) );
OR2_X1 _11723_ ( .A1(_03611_ ), .A2(\myreg.Reg[13][0] ), .ZN(_04068_ ) );
OAI211_X1 _11724_ ( .A(_04068_ ), .B(_04043_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[12][0] ), .ZN(_04069_ ) );
OR2_X1 _11725_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[14][0] ), .ZN(_04070_ ) );
OAI211_X1 _11726_ ( .A(_04070_ ), .B(fanout_net_40 ), .C1(_03612_ ), .C2(\myreg.Reg[15][0] ), .ZN(_04071_ ) );
NAND3_X1 _11727_ ( .A1(_04069_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04071_ ), .ZN(_04072_ ) );
MUX2_X1 _11728_ ( .A(\myreg.Reg[8][0] ), .B(\myreg.Reg[9][0] ), .S(fanout_net_35 ), .Z(_04073_ ) );
MUX2_X1 _11729_ ( .A(\myreg.Reg[10][0] ), .B(\myreg.Reg[11][0] ), .S(fanout_net_35 ), .Z(_04074_ ) );
MUX2_X1 _11730_ ( .A(_04073_ ), .B(_04074_ ), .S(fanout_net_40 ), .Z(_04075_ ) );
OAI211_X1 _11731_ ( .A(fanout_net_43 ), .B(_04072_ ), .C1(_04075_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04076_ ) );
NAND2_X1 _11732_ ( .A1(_04067_ ), .A2(_04076_ ), .ZN(_04077_ ) );
OAI21_X1 _11733_ ( .A(_04077_ ), .B1(_03653_ ), .B2(_03648_ ), .ZN(_04078_ ) );
INV_X1 _11734_ ( .A(\EX_LS_result_reg [0] ), .ZN(_04079_ ) );
OR3_X1 _11735_ ( .A1(_03647_ ), .A2(_04079_ ), .A3(_03642_ ), .ZN(_04080_ ) );
AOI21_X1 _11736_ ( .A(_04058_ ), .B1(_04078_ ), .B2(_04080_ ), .ZN(_04081_ ) );
INV_X1 _11737_ ( .A(_04081_ ), .ZN(_04082_ ) );
NAND3_X1 _11738_ ( .A1(_04058_ ), .A2(_04078_ ), .A3(_04080_ ), .ZN(_04083_ ) );
AND3_X1 _11739_ ( .A1(_04057_ ), .A2(_04082_ ), .A3(_04083_ ), .ZN(_04084_ ) );
OR2_X1 _11740_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04085_ ) );
OAI211_X1 _11741_ ( .A(_04085_ ), .B(_03609_ ), .C1(_03662_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04086_ ) );
OR2_X1 _11742_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04087_ ) );
OAI211_X1 _11743_ ( .A(_04087_ ), .B(fanout_net_40 ), .C1(_03662_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04088_ ) );
NAND3_X1 _11744_ ( .A1(_04086_ ), .A2(_04088_ ), .A3(_03617_ ), .ZN(_04089_ ) );
MUX2_X1 _11745_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04090_ ) );
MUX2_X1 _11746_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04091_ ) );
MUX2_X1 _11747_ ( .A(_04090_ ), .B(_04091_ ), .S(_03608_ ), .Z(_04092_ ) );
OAI211_X1 _11748_ ( .A(_03605_ ), .B(_04089_ ), .C1(_04092_ ), .C2(_03618_ ), .ZN(_04093_ ) );
OR2_X1 _11749_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04094_ ) );
OAI211_X1 _11750_ ( .A(_04094_ ), .B(fanout_net_40 ), .C1(_03662_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04095_ ) );
OR2_X1 _11751_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04096_ ) );
OAI211_X1 _11752_ ( .A(_04096_ ), .B(_03609_ ), .C1(_03611_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04097_ ) );
NAND3_X1 _11753_ ( .A1(_04095_ ), .A2(_04097_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04098_ ) );
MUX2_X1 _11754_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04099_ ) );
MUX2_X1 _11755_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04100_ ) );
MUX2_X1 _11756_ ( .A(_04099_ ), .B(_04100_ ), .S(fanout_net_40 ), .Z(_04101_ ) );
OAI211_X1 _11757_ ( .A(fanout_net_43 ), .B(_04098_ ), .C1(_04101_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04102_ ) );
NAND2_X1 _11758_ ( .A1(_04093_ ), .A2(_04102_ ), .ZN(_04103_ ) );
OAI21_X1 _11759_ ( .A(_04103_ ), .B1(_03643_ ), .B2(_03648_ ), .ZN(_04104_ ) );
NAND2_X1 _11760_ ( .A1(_03941_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04105_ ) );
AND2_X2 _11761_ ( .A1(_04104_ ), .A2(_04105_ ), .ZN(_04106_ ) );
XNOR2_X1 _11762_ ( .A(_02732_ ), .B(_04106_ ), .ZN(_04107_ ) );
INV_X1 _11763_ ( .A(_02755_ ), .ZN(_04108_ ) );
OR2_X1 _11764_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[8][2] ), .ZN(_04109_ ) );
OAI211_X1 _11765_ ( .A(_04109_ ), .B(_03610_ ), .C1(_03663_ ), .C2(\myreg.Reg[9][2] ), .ZN(_04110_ ) );
OR2_X1 _11766_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[10][2] ), .ZN(_04111_ ) );
OAI211_X1 _11767_ ( .A(_04111_ ), .B(fanout_net_40 ), .C1(_03663_ ), .C2(\myreg.Reg[11][2] ), .ZN(_04112_ ) );
NAND3_X1 _11768_ ( .A1(_04110_ ), .A2(_04112_ ), .A3(_03619_ ), .ZN(_04113_ ) );
MUX2_X1 _11769_ ( .A(\myreg.Reg[14][2] ), .B(\myreg.Reg[15][2] ), .S(fanout_net_36 ), .Z(_04114_ ) );
MUX2_X1 _11770_ ( .A(\myreg.Reg[12][2] ), .B(\myreg.Reg[13][2] ), .S(fanout_net_36 ), .Z(_04115_ ) );
MUX2_X1 _11771_ ( .A(_04114_ ), .B(_04115_ ), .S(_03705_ ), .Z(_04116_ ) );
OAI211_X1 _11772_ ( .A(fanout_net_43 ), .B(_04113_ ), .C1(_04116_ ), .C2(_03708_ ), .ZN(_04117_ ) );
MUX2_X1 _11773_ ( .A(\myreg.Reg[0][2] ), .B(\myreg.Reg[1][2] ), .S(fanout_net_36 ), .Z(_04118_ ) );
AND2_X1 _11774_ ( .A1(_04118_ ), .A2(_03705_ ), .ZN(_04119_ ) );
MUX2_X1 _11775_ ( .A(\myreg.Reg[2][2] ), .B(\myreg.Reg[3][2] ), .S(fanout_net_36 ), .Z(_04120_ ) );
AOI211_X1 _11776_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_04119_ ), .C1(fanout_net_40 ), .C2(_04120_ ), .ZN(_04121_ ) );
MUX2_X1 _11777_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_36 ), .Z(_04122_ ) );
MUX2_X1 _11778_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_36 ), .Z(_04123_ ) );
MUX2_X1 _11779_ ( .A(_04122_ ), .B(_04123_ ), .S(_04043_ ), .Z(_04124_ ) );
OAI21_X1 _11780_ ( .A(_03606_ ), .B1(_04124_ ), .B2(_03708_ ), .ZN(_04125_ ) );
OAI221_X1 _11781_ ( .A(_04117_ ), .B1(_03648_ ), .B2(_03643_ ), .C1(_04121_ ), .C2(_04125_ ), .ZN(_04126_ ) );
OR3_X4 _11782_ ( .A1(_03648_ ), .A2(\EX_LS_result_reg [2] ), .A3(_03643_ ), .ZN(_04127_ ) );
NAND2_X1 _11783_ ( .A1(_04126_ ), .A2(_04127_ ), .ZN(_04128_ ) );
XNOR2_X1 _11784_ ( .A(_04108_ ), .B(_04128_ ), .ZN(_04129_ ) );
AND3_X1 _11785_ ( .A1(_04084_ ), .A2(_04107_ ), .A3(_04129_ ), .ZN(_04130_ ) );
OR2_X1 _11786_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[0][15] ), .ZN(_04131_ ) );
OAI211_X1 _11787_ ( .A(_04131_ ), .B(_03609_ ), .C1(_03612_ ), .C2(\myreg.Reg[1][15] ), .ZN(_04132_ ) );
OR2_X1 _11788_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[2][15] ), .ZN(_04133_ ) );
OAI211_X1 _11789_ ( .A(_04133_ ), .B(fanout_net_40 ), .C1(_03662_ ), .C2(\myreg.Reg[3][15] ), .ZN(_04134_ ) );
NAND3_X1 _11790_ ( .A1(_04132_ ), .A2(_04134_ ), .A3(_03618_ ), .ZN(_04135_ ) );
MUX2_X1 _11791_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_36 ), .Z(_04136_ ) );
MUX2_X1 _11792_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_36 ), .Z(_04137_ ) );
MUX2_X1 _11793_ ( .A(_04136_ ), .B(_04137_ ), .S(_03609_ ), .Z(_04138_ ) );
OAI211_X1 _11794_ ( .A(_03605_ ), .B(_04135_ ), .C1(_04138_ ), .C2(_03618_ ), .ZN(_04139_ ) );
OR2_X1 _11795_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][15] ), .ZN(_04140_ ) );
OAI211_X1 _11796_ ( .A(_04140_ ), .B(fanout_net_40 ), .C1(_03662_ ), .C2(\myreg.Reg[15][15] ), .ZN(_04141_ ) );
OR2_X1 _11797_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[12][15] ), .ZN(_04142_ ) );
OAI211_X1 _11798_ ( .A(_04142_ ), .B(_03609_ ), .C1(_03662_ ), .C2(\myreg.Reg[13][15] ), .ZN(_04143_ ) );
NAND3_X1 _11799_ ( .A1(_04141_ ), .A2(_04143_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04144_ ) );
MUX2_X1 _11800_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_36 ), .Z(_04145_ ) );
MUX2_X1 _11801_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_36 ), .Z(_04146_ ) );
MUX2_X1 _11802_ ( .A(_04145_ ), .B(_04146_ ), .S(fanout_net_40 ), .Z(_04147_ ) );
OAI211_X1 _11803_ ( .A(fanout_net_43 ), .B(_04144_ ), .C1(_04147_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04148_ ) );
NAND2_X1 _11804_ ( .A1(_04139_ ), .A2(_04148_ ), .ZN(_04149_ ) );
OAI21_X1 _11805_ ( .A(_04149_ ), .B1(_03643_ ), .B2(_03648_ ), .ZN(_04150_ ) );
INV_X1 _11806_ ( .A(\EX_LS_result_reg [15] ), .ZN(_04151_ ) );
OR3_X1 _11807_ ( .A1(_03647_ ), .A2(_04151_ ), .A3(_03642_ ), .ZN(_04152_ ) );
AND2_X1 _11808_ ( .A1(_04150_ ), .A2(_04152_ ), .ZN(_04153_ ) );
INV_X1 _11809_ ( .A(_03094_ ), .ZN(_04154_ ) );
XNOR2_X1 _11810_ ( .A(_04153_ ), .B(_04154_ ), .ZN(_04155_ ) );
OR3_X1 _11811_ ( .A1(_03649_ ), .A2(\EX_LS_result_reg [14] ), .A3(_03644_ ), .ZN(_04156_ ) );
OR2_X1 _11812_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[4][14] ), .ZN(_04157_ ) );
OAI211_X1 _11813_ ( .A(_04157_ ), .B(_03677_ ), .C1(_03671_ ), .C2(\myreg.Reg[5][14] ), .ZN(_04158_ ) );
OR2_X1 _11814_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[6][14] ), .ZN(_04159_ ) );
OAI211_X1 _11815_ ( .A(_04159_ ), .B(fanout_net_41 ), .C1(_03671_ ), .C2(\myreg.Reg[7][14] ), .ZN(_04160_ ) );
NAND3_X1 _11816_ ( .A1(_04158_ ), .A2(_04160_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04161_ ) );
MUX2_X1 _11817_ ( .A(\myreg.Reg[2][14] ), .B(\myreg.Reg[3][14] ), .S(fanout_net_36 ), .Z(_04162_ ) );
MUX2_X1 _11818_ ( .A(\myreg.Reg[0][14] ), .B(\myreg.Reg[1][14] ), .S(fanout_net_36 ), .Z(_04163_ ) );
MUX2_X1 _11819_ ( .A(_04162_ ), .B(_04163_ ), .S(_03669_ ), .Z(_04164_ ) );
OAI211_X1 _11820_ ( .A(_03661_ ), .B(_04161_ ), .C1(_04164_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04165_ ) );
NOR2_X1 _11821_ ( .A1(_03664_ ), .A2(\myreg.Reg[11][14] ), .ZN(_04166_ ) );
OAI21_X1 _11822_ ( .A(fanout_net_41 ), .B1(fanout_net_36 ), .B2(\myreg.Reg[10][14] ), .ZN(_04167_ ) );
NOR2_X1 _11823_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[8][14] ), .ZN(_04168_ ) );
OAI21_X1 _11824_ ( .A(_03669_ ), .B1(_03671_ ), .B2(\myreg.Reg[9][14] ), .ZN(_04169_ ) );
OAI221_X1 _11825_ ( .A(_03624_ ), .B1(_04166_ ), .B2(_04167_ ), .C1(_04168_ ), .C2(_04169_ ), .ZN(_04170_ ) );
MUX2_X1 _11826_ ( .A(\myreg.Reg[12][14] ), .B(\myreg.Reg[13][14] ), .S(fanout_net_36 ), .Z(_04171_ ) );
MUX2_X1 _11827_ ( .A(\myreg.Reg[14][14] ), .B(\myreg.Reg[15][14] ), .S(fanout_net_36 ), .Z(_04172_ ) );
MUX2_X1 _11828_ ( .A(_04171_ ), .B(_04172_ ), .S(fanout_net_41 ), .Z(_04173_ ) );
OAI211_X1 _11829_ ( .A(fanout_net_43 ), .B(_04170_ ), .C1(_04173_ ), .C2(_03709_ ), .ZN(_04174_ ) );
OAI211_X1 _11830_ ( .A(_04165_ ), .B(_04174_ ), .C1(_03658_ ), .C2(_03659_ ), .ZN(_04175_ ) );
NAND2_X1 _11831_ ( .A1(_04156_ ), .A2(_04175_ ), .ZN(_04176_ ) );
XOR2_X1 _11832_ ( .A(_04176_ ), .B(_03118_ ), .Z(_04177_ ) );
AND2_X1 _11833_ ( .A1(_04155_ ), .A2(_04177_ ), .ZN(_04178_ ) );
NAND2_X1 _11834_ ( .A1(_03044_ ), .A2(_03046_ ), .ZN(_04179_ ) );
OR3_X1 _11835_ ( .A1(_03651_ ), .A2(\EX_LS_result_reg [13] ), .A3(_03653_ ), .ZN(_04180_ ) );
OR2_X1 _11836_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[4][13] ), .ZN(_04181_ ) );
OAI211_X1 _11837_ ( .A(_04181_ ), .B(_03706_ ), .C1(_03700_ ), .C2(\myreg.Reg[5][13] ), .ZN(_04182_ ) );
OR2_X1 _11838_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[6][13] ), .ZN(_04183_ ) );
OAI211_X1 _11839_ ( .A(_04183_ ), .B(fanout_net_41 ), .C1(_03700_ ), .C2(\myreg.Reg[7][13] ), .ZN(_04184_ ) );
NAND3_X1 _11840_ ( .A1(_04182_ ), .A2(_04184_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04185_ ) );
MUX2_X1 _11841_ ( .A(\myreg.Reg[2][13] ), .B(\myreg.Reg[3][13] ), .S(fanout_net_37 ), .Z(_04186_ ) );
MUX2_X1 _11842_ ( .A(\myreg.Reg[0][13] ), .B(\myreg.Reg[1][13] ), .S(fanout_net_37 ), .Z(_04187_ ) );
MUX2_X1 _11843_ ( .A(_04186_ ), .B(_04187_ ), .S(_03706_ ), .Z(_04188_ ) );
OAI211_X1 _11844_ ( .A(_03606_ ), .B(_04185_ ), .C1(_04188_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04189_ ) );
NOR2_X1 _11845_ ( .A1(_03700_ ), .A2(\myreg.Reg[11][13] ), .ZN(_04190_ ) );
OAI21_X1 _11846_ ( .A(fanout_net_41 ), .B1(fanout_net_37 ), .B2(\myreg.Reg[10][13] ), .ZN(_04191_ ) );
NOR2_X1 _11847_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][13] ), .ZN(_04192_ ) );
OAI21_X1 _11848_ ( .A(_03706_ ), .B1(_03700_ ), .B2(\myreg.Reg[9][13] ), .ZN(_04193_ ) );
OAI221_X1 _11849_ ( .A(_03708_ ), .B1(_04190_ ), .B2(_04191_ ), .C1(_04192_ ), .C2(_04193_ ), .ZN(_04194_ ) );
MUX2_X1 _11850_ ( .A(\myreg.Reg[12][13] ), .B(\myreg.Reg[13][13] ), .S(fanout_net_37 ), .Z(_04195_ ) );
MUX2_X1 _11851_ ( .A(\myreg.Reg[14][13] ), .B(\myreg.Reg[15][13] ), .S(fanout_net_37 ), .Z(_04196_ ) );
MUX2_X1 _11852_ ( .A(_04195_ ), .B(_04196_ ), .S(fanout_net_41 ), .Z(_04197_ ) );
OAI211_X1 _11853_ ( .A(fanout_net_43 ), .B(_04194_ ), .C1(_04197_ ), .C2(_03624_ ), .ZN(_04198_ ) );
OAI211_X1 _11854_ ( .A(_04189_ ), .B(_04198_ ), .C1(_03649_ ), .C2(_03644_ ), .ZN(_04199_ ) );
NAND2_X1 _11855_ ( .A1(_04180_ ), .A2(_04199_ ), .ZN(_04200_ ) );
XOR2_X1 _11856_ ( .A(_04179_ ), .B(_04200_ ), .Z(_04201_ ) );
OR3_X1 _11857_ ( .A1(_03651_ ), .A2(\EX_LS_result_reg [12] ), .A3(_03653_ ), .ZN(_04202_ ) );
OR2_X1 _11858_ ( .A1(_03663_ ), .A2(\myreg.Reg[1][12] ), .ZN(_04203_ ) );
OAI211_X1 _11859_ ( .A(_04203_ ), .B(_03669_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[0][12] ), .ZN(_04204_ ) );
OR2_X1 _11860_ ( .A1(_03663_ ), .A2(\myreg.Reg[3][12] ), .ZN(_04205_ ) );
OAI211_X1 _11861_ ( .A(_04205_ ), .B(fanout_net_41 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[2][12] ), .ZN(_04206_ ) );
NAND3_X1 _11862_ ( .A1(_04204_ ), .A2(_04206_ ), .A3(_03624_ ), .ZN(_04207_ ) );
MUX2_X1 _11863_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_37 ), .Z(_04208_ ) );
MUX2_X1 _11864_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_37 ), .Z(_04209_ ) );
MUX2_X1 _11865_ ( .A(_04208_ ), .B(_04209_ ), .S(_03706_ ), .Z(_04210_ ) );
OAI211_X1 _11866_ ( .A(_03661_ ), .B(_04207_ ), .C1(_04210_ ), .C2(_03709_ ), .ZN(_04211_ ) );
OR2_X1 _11867_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[14][12] ), .ZN(_04212_ ) );
OAI211_X1 _11868_ ( .A(_04212_ ), .B(fanout_net_41 ), .C1(_03664_ ), .C2(\myreg.Reg[15][12] ), .ZN(_04213_ ) );
OR2_X1 _11869_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][12] ), .ZN(_04214_ ) );
OAI211_X1 _11870_ ( .A(_04214_ ), .B(_03706_ ), .C1(_03700_ ), .C2(\myreg.Reg[13][12] ), .ZN(_04215_ ) );
NAND3_X1 _11871_ ( .A1(_04213_ ), .A2(_04215_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04216_ ) );
MUX2_X1 _11872_ ( .A(\myreg.Reg[8][12] ), .B(\myreg.Reg[9][12] ), .S(fanout_net_37 ), .Z(_04217_ ) );
MUX2_X1 _11873_ ( .A(\myreg.Reg[10][12] ), .B(\myreg.Reg[11][12] ), .S(fanout_net_37 ), .Z(_04218_ ) );
MUX2_X1 _11874_ ( .A(_04217_ ), .B(_04218_ ), .S(fanout_net_41 ), .Z(_04219_ ) );
OAI211_X1 _11875_ ( .A(fanout_net_43 ), .B(_04216_ ), .C1(_04219_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04220_ ) );
OAI211_X1 _11876_ ( .A(_04211_ ), .B(_04220_ ), .C1(_03649_ ), .C2(_03644_ ), .ZN(_04221_ ) );
NAND2_X1 _11877_ ( .A1(_04202_ ), .A2(_04221_ ), .ZN(_04222_ ) );
XOR2_X1 _11878_ ( .A(_04222_ ), .B(_03070_ ), .Z(_04223_ ) );
AND3_X1 _11879_ ( .A1(_04178_ ), .A2(_04201_ ), .A3(_04223_ ), .ZN(_04224_ ) );
OR2_X1 _11880_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][11] ), .ZN(_04225_ ) );
OAI211_X1 _11881_ ( .A(_04225_ ), .B(_03609_ ), .C1(_03612_ ), .C2(\myreg.Reg[1][11] ), .ZN(_04226_ ) );
OR2_X1 _11882_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][11] ), .ZN(_04227_ ) );
OAI211_X1 _11883_ ( .A(_04227_ ), .B(fanout_net_41 ), .C1(_03612_ ), .C2(\myreg.Reg[3][11] ), .ZN(_04228_ ) );
NAND3_X1 _11884_ ( .A1(_04226_ ), .A2(_04228_ ), .A3(_03618_ ), .ZN(_04229_ ) );
MUX2_X1 _11885_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_37 ), .Z(_04230_ ) );
MUX2_X1 _11886_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_37 ), .Z(_04231_ ) );
MUX2_X1 _11887_ ( .A(_04230_ ), .B(_04231_ ), .S(_03609_ ), .Z(_04232_ ) );
OAI211_X1 _11888_ ( .A(_03605_ ), .B(_04229_ ), .C1(_04232_ ), .C2(_03618_ ), .ZN(_04233_ ) );
OR2_X1 _11889_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[14][11] ), .ZN(_04234_ ) );
OAI211_X1 _11890_ ( .A(_04234_ ), .B(fanout_net_41 ), .C1(_03612_ ), .C2(\myreg.Reg[15][11] ), .ZN(_04235_ ) );
OR2_X1 _11891_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][11] ), .ZN(_04236_ ) );
OAI211_X1 _11892_ ( .A(_04236_ ), .B(_03609_ ), .C1(_03662_ ), .C2(\myreg.Reg[13][11] ), .ZN(_04237_ ) );
NAND3_X1 _11893_ ( .A1(_04235_ ), .A2(_04237_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04238_ ) );
MUX2_X1 _11894_ ( .A(\myreg.Reg[8][11] ), .B(\myreg.Reg[9][11] ), .S(fanout_net_37 ), .Z(_04239_ ) );
MUX2_X1 _11895_ ( .A(\myreg.Reg[10][11] ), .B(\myreg.Reg[11][11] ), .S(fanout_net_37 ), .Z(_04240_ ) );
MUX2_X1 _11896_ ( .A(_04239_ ), .B(_04240_ ), .S(fanout_net_41 ), .Z(_04241_ ) );
OAI211_X1 _11897_ ( .A(fanout_net_43 ), .B(_04238_ ), .C1(_04241_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04242_ ) );
NAND2_X1 _11898_ ( .A1(_04233_ ), .A2(_04242_ ), .ZN(_04243_ ) );
OAI21_X1 _11899_ ( .A(_04243_ ), .B1(_03643_ ), .B2(_03648_ ), .ZN(_04244_ ) );
INV_X1 _11900_ ( .A(\EX_LS_result_reg [11] ), .ZN(_04245_ ) );
OR3_X1 _11901_ ( .A1(_03647_ ), .A2(_04245_ ), .A3(_03642_ ), .ZN(_04246_ ) );
AND2_X1 _11902_ ( .A1(_04244_ ), .A2(_04246_ ), .ZN(_04247_ ) );
NAND2_X1 _11903_ ( .A1(_02967_ ), .A2(_02987_ ), .ZN(_04248_ ) );
INV_X1 _11904_ ( .A(_04248_ ), .ZN(_04249_ ) );
XNOR2_X1 _11905_ ( .A(_04247_ ), .B(_04249_ ), .ZN(_04250_ ) );
OR3_X1 _11906_ ( .A1(_03649_ ), .A2(\EX_LS_result_reg [10] ), .A3(_03644_ ), .ZN(_04251_ ) );
OR2_X1 _11907_ ( .A1(_03613_ ), .A2(\myreg.Reg[3][10] ), .ZN(_04252_ ) );
OAI211_X1 _11908_ ( .A(_04252_ ), .B(fanout_net_41 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[2][10] ), .ZN(_04253_ ) );
OR2_X1 _11909_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][10] ), .ZN(_04254_ ) );
OAI211_X1 _11910_ ( .A(_04254_ ), .B(_03677_ ), .C1(_03671_ ), .C2(\myreg.Reg[1][10] ), .ZN(_04255_ ) );
NAND3_X1 _11911_ ( .A1(_04253_ ), .A2(_03624_ ), .A3(_04255_ ), .ZN(_04256_ ) );
MUX2_X1 _11912_ ( .A(\myreg.Reg[6][10] ), .B(\myreg.Reg[7][10] ), .S(fanout_net_37 ), .Z(_04257_ ) );
MUX2_X1 _11913_ ( .A(\myreg.Reg[4][10] ), .B(\myreg.Reg[5][10] ), .S(fanout_net_37 ), .Z(_04258_ ) );
MUX2_X1 _11914_ ( .A(_04257_ ), .B(_04258_ ), .S(_03669_ ), .Z(_04259_ ) );
OAI211_X1 _11915_ ( .A(_03661_ ), .B(_04256_ ), .C1(_04259_ ), .C2(_03709_ ), .ZN(_04260_ ) );
OR2_X1 _11916_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[14][10] ), .ZN(_04261_ ) );
OAI211_X1 _11917_ ( .A(_04261_ ), .B(fanout_net_41 ), .C1(_03671_ ), .C2(\myreg.Reg[15][10] ), .ZN(_04262_ ) );
OR2_X1 _11918_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][10] ), .ZN(_04263_ ) );
OAI211_X1 _11919_ ( .A(_04263_ ), .B(_03669_ ), .C1(_03671_ ), .C2(\myreg.Reg[13][10] ), .ZN(_04264_ ) );
NAND3_X1 _11920_ ( .A1(_04262_ ), .A2(_04264_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04265_ ) );
MUX2_X1 _11921_ ( .A(\myreg.Reg[8][10] ), .B(\myreg.Reg[9][10] ), .S(fanout_net_37 ), .Z(_04266_ ) );
MUX2_X1 _11922_ ( .A(\myreg.Reg[10][10] ), .B(\myreg.Reg[11][10] ), .S(fanout_net_37 ), .Z(_04267_ ) );
MUX2_X1 _11923_ ( .A(_04266_ ), .B(_04267_ ), .S(fanout_net_41 ), .Z(_04268_ ) );
OAI211_X1 _11924_ ( .A(fanout_net_43 ), .B(_04265_ ), .C1(_04268_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04269_ ) );
OAI211_X1 _11925_ ( .A(_04260_ ), .B(_04269_ ), .C1(_03658_ ), .C2(_03659_ ), .ZN(_04270_ ) );
NAND2_X1 _11926_ ( .A1(_04251_ ), .A2(_04270_ ), .ZN(_04271_ ) );
XOR2_X1 _11927_ ( .A(_04271_ ), .B(_03012_ ), .Z(_04272_ ) );
AND2_X1 _11928_ ( .A1(_04250_ ), .A2(_04272_ ), .ZN(_04273_ ) );
OR2_X1 _11929_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][9] ), .ZN(_04274_ ) );
OAI211_X1 _11930_ ( .A(_04274_ ), .B(_03610_ ), .C1(_03613_ ), .C2(\myreg.Reg[1][9] ), .ZN(_04275_ ) );
OR2_X1 _11931_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[2][9] ), .ZN(_04276_ ) );
OAI211_X1 _11932_ ( .A(_04276_ ), .B(fanout_net_41 ), .C1(_03613_ ), .C2(\myreg.Reg[3][9] ), .ZN(_04277_ ) );
NAND3_X1 _11933_ ( .A1(_04275_ ), .A2(_04277_ ), .A3(_03619_ ), .ZN(_04278_ ) );
MUX2_X1 _11934_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_38 ), .Z(_04279_ ) );
MUX2_X1 _11935_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_38 ), .Z(_04280_ ) );
MUX2_X1 _11936_ ( .A(_04279_ ), .B(_04280_ ), .S(_03610_ ), .Z(_04281_ ) );
OAI211_X1 _11937_ ( .A(_03606_ ), .B(_04278_ ), .C1(_04281_ ), .C2(_03708_ ), .ZN(_04282_ ) );
OR2_X1 _11938_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[14][9] ), .ZN(_04283_ ) );
OAI211_X1 _11939_ ( .A(_04283_ ), .B(fanout_net_41 ), .C1(_03613_ ), .C2(\myreg.Reg[15][9] ), .ZN(_04284_ ) );
OR2_X1 _11940_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[12][9] ), .ZN(_04285_ ) );
OAI211_X1 _11941_ ( .A(_04285_ ), .B(_03610_ ), .C1(_03613_ ), .C2(\myreg.Reg[13][9] ), .ZN(_04286_ ) );
NAND3_X1 _11942_ ( .A1(_04284_ ), .A2(_04286_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04287_ ) );
MUX2_X1 _11943_ ( .A(\myreg.Reg[8][9] ), .B(\myreg.Reg[9][9] ), .S(fanout_net_38 ), .Z(_04288_ ) );
MUX2_X1 _11944_ ( .A(\myreg.Reg[10][9] ), .B(\myreg.Reg[11][9] ), .S(fanout_net_38 ), .Z(_04289_ ) );
MUX2_X1 _11945_ ( .A(_04288_ ), .B(_04289_ ), .S(fanout_net_41 ), .Z(_04290_ ) );
OAI211_X1 _11946_ ( .A(fanout_net_43 ), .B(_04287_ ), .C1(_04290_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04291_ ) );
NAND2_X1 _11947_ ( .A1(_04282_ ), .A2(_04291_ ), .ZN(_04292_ ) );
OAI21_X1 _11948_ ( .A(_04292_ ), .B1(_03644_ ), .B2(_03649_ ), .ZN(_04293_ ) );
INV_X1 _11949_ ( .A(\EX_LS_result_reg [9] ), .ZN(_04294_ ) );
OR3_X1 _11950_ ( .A1(_03651_ ), .A2(_04294_ ), .A3(_03643_ ), .ZN(_04295_ ) );
AND2_X1 _11951_ ( .A1(_04293_ ), .A2(_04295_ ), .ZN(_04296_ ) );
INV_X1 _11952_ ( .A(_02963_ ), .ZN(_04297_ ) );
XNOR2_X1 _11953_ ( .A(_04296_ ), .B(_04297_ ), .ZN(_04298_ ) );
OR3_X1 _11954_ ( .A1(_03649_ ), .A2(\EX_LS_result_reg [8] ), .A3(_03644_ ), .ZN(_04299_ ) );
OR2_X1 _11955_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[4][8] ), .ZN(_04300_ ) );
OAI211_X1 _11956_ ( .A(_04300_ ), .B(_03669_ ), .C1(_03664_ ), .C2(\myreg.Reg[5][8] ), .ZN(_04301_ ) );
OR2_X1 _11957_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[6][8] ), .ZN(_04302_ ) );
OAI211_X1 _11958_ ( .A(_04302_ ), .B(fanout_net_41 ), .C1(_03664_ ), .C2(\myreg.Reg[7][8] ), .ZN(_04303_ ) );
NAND3_X1 _11959_ ( .A1(_04301_ ), .A2(_04303_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04304_ ) );
MUX2_X1 _11960_ ( .A(\myreg.Reg[2][8] ), .B(\myreg.Reg[3][8] ), .S(fanout_net_38 ), .Z(_04305_ ) );
MUX2_X1 _11961_ ( .A(\myreg.Reg[0][8] ), .B(\myreg.Reg[1][8] ), .S(fanout_net_38 ), .Z(_04306_ ) );
MUX2_X1 _11962_ ( .A(_04305_ ), .B(_04306_ ), .S(_03669_ ), .Z(_04307_ ) );
OAI211_X1 _11963_ ( .A(_03661_ ), .B(_04304_ ), .C1(_04307_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04308_ ) );
NOR2_X1 _11964_ ( .A1(_03700_ ), .A2(\myreg.Reg[11][8] ), .ZN(_04309_ ) );
OAI21_X1 _11965_ ( .A(fanout_net_41 ), .B1(fanout_net_38 ), .B2(\myreg.Reg[10][8] ), .ZN(_04310_ ) );
NOR2_X1 _11966_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[8][8] ), .ZN(_04311_ ) );
OAI21_X1 _11967_ ( .A(_03669_ ), .B1(_03664_ ), .B2(\myreg.Reg[9][8] ), .ZN(_04312_ ) );
OAI221_X1 _11968_ ( .A(_03624_ ), .B1(_04309_ ), .B2(_04310_ ), .C1(_04311_ ), .C2(_04312_ ), .ZN(_04313_ ) );
MUX2_X1 _11969_ ( .A(\myreg.Reg[12][8] ), .B(\myreg.Reg[13][8] ), .S(fanout_net_38 ), .Z(_04314_ ) );
MUX2_X1 _11970_ ( .A(\myreg.Reg[14][8] ), .B(\myreg.Reg[15][8] ), .S(fanout_net_38 ), .Z(_04315_ ) );
MUX2_X1 _11971_ ( .A(_04314_ ), .B(_04315_ ), .S(fanout_net_41 ), .Z(_04316_ ) );
OAI211_X1 _11972_ ( .A(fanout_net_43 ), .B(_04313_ ), .C1(_04316_ ), .C2(_03709_ ), .ZN(_04317_ ) );
OAI211_X1 _11973_ ( .A(_04308_ ), .B(_04317_ ), .C1(_03649_ ), .C2(_03659_ ), .ZN(_04318_ ) );
NAND2_X1 _11974_ ( .A1(_04299_ ), .A2(_04318_ ), .ZN(_04319_ ) );
XOR2_X1 _11975_ ( .A(_04319_ ), .B(_02938_ ), .Z(_04320_ ) );
AND3_X1 _11976_ ( .A1(_04273_ ), .A2(_04298_ ), .A3(_04320_ ), .ZN(_04321_ ) );
OR3_X1 _11977_ ( .A1(_03648_ ), .A2(\EX_LS_result_reg [7] ), .A3(_03643_ ), .ZN(_04322_ ) );
OR2_X1 _11978_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[8][7] ), .ZN(_04323_ ) );
OAI211_X1 _11979_ ( .A(_04323_ ), .B(_03705_ ), .C1(_03699_ ), .C2(\myreg.Reg[9][7] ), .ZN(_04324_ ) );
OR2_X1 _11980_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[10][7] ), .ZN(_04325_ ) );
OAI211_X1 _11981_ ( .A(_04325_ ), .B(fanout_net_41 ), .C1(_03699_ ), .C2(\myreg.Reg[11][7] ), .ZN(_04326_ ) );
NAND3_X1 _11982_ ( .A1(_04324_ ), .A2(_04326_ ), .A3(_03619_ ), .ZN(_04327_ ) );
MUX2_X1 _11983_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_38 ), .Z(_04328_ ) );
MUX2_X1 _11984_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_38 ), .Z(_04329_ ) );
MUX2_X1 _11985_ ( .A(_04328_ ), .B(_04329_ ), .S(_04043_ ), .Z(_04330_ ) );
OAI211_X1 _11986_ ( .A(fanout_net_43 ), .B(_04327_ ), .C1(_04330_ ), .C2(_03708_ ), .ZN(_04331_ ) );
OAI21_X1 _11987_ ( .A(_04043_ ), .B1(_03612_ ), .B2(\myreg.Reg[1][7] ), .ZN(_04332_ ) );
NOR2_X1 _11988_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][7] ), .ZN(_04333_ ) );
NOR2_X1 _11989_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[2][7] ), .ZN(_04334_ ) );
OAI21_X1 _11990_ ( .A(fanout_net_41 ), .B1(_03699_ ), .B2(\myreg.Reg[3][7] ), .ZN(_04335_ ) );
OAI221_X1 _11991_ ( .A(_03618_ ), .B1(_04332_ ), .B2(_04333_ ), .C1(_04334_ ), .C2(_04335_ ), .ZN(_04336_ ) );
MUX2_X1 _11992_ ( .A(\myreg.Reg[6][7] ), .B(\myreg.Reg[7][7] ), .S(fanout_net_38 ), .Z(_04337_ ) );
MUX2_X1 _11993_ ( .A(\myreg.Reg[4][7] ), .B(\myreg.Reg[5][7] ), .S(fanout_net_38 ), .Z(_04338_ ) );
MUX2_X1 _11994_ ( .A(_04337_ ), .B(_04338_ ), .S(_04043_ ), .Z(_04339_ ) );
OAI211_X1 _11995_ ( .A(_03606_ ), .B(_04336_ ), .C1(_04339_ ), .C2(_03708_ ), .ZN(_04340_ ) );
OAI211_X1 _11996_ ( .A(_04331_ ), .B(_04340_ ), .C1(_03651_ ), .C2(_03653_ ), .ZN(_04341_ ) );
NAND2_X2 _11997_ ( .A1(_04322_ ), .A2(_04341_ ), .ZN(_04342_ ) );
XOR2_X1 _11998_ ( .A(_02886_ ), .B(_04342_ ), .Z(_04343_ ) );
OR3_X4 _11999_ ( .A1(_03648_ ), .A2(\EX_LS_result_reg [6] ), .A3(_03643_ ), .ZN(_04344_ ) );
OR2_X1 _12000_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[8][6] ), .ZN(_04345_ ) );
OAI211_X1 _12001_ ( .A(_04345_ ), .B(_03705_ ), .C1(_03663_ ), .C2(\myreg.Reg[9][6] ), .ZN(_04346_ ) );
OR2_X1 _12002_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[10][6] ), .ZN(_04347_ ) );
OAI211_X1 _12003_ ( .A(_04347_ ), .B(fanout_net_41 ), .C1(_03699_ ), .C2(\myreg.Reg[11][6] ), .ZN(_04348_ ) );
NAND3_X1 _12004_ ( .A1(_04346_ ), .A2(_04348_ ), .A3(_03619_ ), .ZN(_04349_ ) );
MUX2_X1 _12005_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(fanout_net_38 ), .Z(_04350_ ) );
MUX2_X1 _12006_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(fanout_net_38 ), .Z(_04351_ ) );
MUX2_X1 _12007_ ( .A(_04350_ ), .B(_04351_ ), .S(_03705_ ), .Z(_04352_ ) );
OAI211_X1 _12008_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04349_ ), .C1(_04352_ ), .C2(_03708_ ), .ZN(_04353_ ) );
OR2_X1 _12009_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][6] ), .ZN(_04354_ ) );
OAI211_X1 _12010_ ( .A(_04354_ ), .B(_03705_ ), .C1(_03699_ ), .C2(\myreg.Reg[1][6] ), .ZN(_04355_ ) );
NOR2_X1 _12011_ ( .A1(_03663_ ), .A2(\myreg.Reg[3][6] ), .ZN(_04356_ ) );
OAI21_X1 _12012_ ( .A(fanout_net_41 ), .B1(fanout_net_38 ), .B2(\myreg.Reg[2][6] ), .ZN(_04357_ ) );
OAI211_X1 _12013_ ( .A(_04355_ ), .B(_03619_ ), .C1(_04356_ ), .C2(_04357_ ), .ZN(_04358_ ) );
MUX2_X1 _12014_ ( .A(\myreg.Reg[6][6] ), .B(\myreg.Reg[7][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04359_ ) );
MUX2_X1 _12015_ ( .A(\myreg.Reg[4][6] ), .B(\myreg.Reg[5][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04360_ ) );
MUX2_X1 _12016_ ( .A(_04359_ ), .B(_04360_ ), .S(_04043_ ), .Z(_04361_ ) );
OAI211_X1 _12017_ ( .A(_03606_ ), .B(_04358_ ), .C1(_04361_ ), .C2(_03708_ ), .ZN(_04362_ ) );
OAI211_X1 _12018_ ( .A(_04353_ ), .B(_04362_ ), .C1(_03651_ ), .C2(_03653_ ), .ZN(_04363_ ) );
NAND2_X2 _12019_ ( .A1(_04344_ ), .A2(_04363_ ), .ZN(_04364_ ) );
NAND2_X1 _12020_ ( .A1(_04364_ ), .A2(_02908_ ), .ZN(_04365_ ) );
NAND4_X1 _12021_ ( .A1(_02888_ ), .A2(_04344_ ), .A3(_02907_ ), .A4(_04363_ ), .ZN(_04366_ ) );
AND2_X1 _12022_ ( .A1(_04365_ ), .A2(_04366_ ), .ZN(_04367_ ) );
AND2_X1 _12023_ ( .A1(_04343_ ), .A2(_04367_ ), .ZN(_04368_ ) );
OR3_X1 _12024_ ( .A1(_03651_ ), .A2(\EX_LS_result_reg [4] ), .A3(_03653_ ), .ZN(_04369_ ) );
OR2_X1 _12025_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[0][4] ), .ZN(_04370_ ) );
OAI211_X1 _12026_ ( .A(_04370_ ), .B(_03706_ ), .C1(_03664_ ), .C2(\myreg.Reg[1][4] ), .ZN(_04371_ ) );
OR2_X1 _12027_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[2][4] ), .ZN(_04372_ ) );
OAI211_X1 _12028_ ( .A(_04372_ ), .B(fanout_net_41 ), .C1(_03700_ ), .C2(\myreg.Reg[3][4] ), .ZN(_04373_ ) );
NAND3_X1 _12029_ ( .A1(_04371_ ), .A2(_04373_ ), .A3(_03624_ ), .ZN(_04374_ ) );
MUX2_X1 _12030_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04375_ ) );
MUX2_X1 _12031_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04376_ ) );
MUX2_X1 _12032_ ( .A(_04375_ ), .B(_04376_ ), .S(_03706_ ), .Z(_04377_ ) );
OAI211_X1 _12033_ ( .A(_03661_ ), .B(_04374_ ), .C1(_04377_ ), .C2(_03709_ ), .ZN(_04378_ ) );
OR2_X1 _12034_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[14][4] ), .ZN(_04379_ ) );
OAI211_X1 _12035_ ( .A(_04379_ ), .B(fanout_net_41 ), .C1(_03700_ ), .C2(\myreg.Reg[15][4] ), .ZN(_04380_ ) );
OR2_X1 _12036_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[12][4] ), .ZN(_04381_ ) );
OAI211_X1 _12037_ ( .A(_04381_ ), .B(_03706_ ), .C1(_03700_ ), .C2(\myreg.Reg[13][4] ), .ZN(_04382_ ) );
NAND3_X1 _12038_ ( .A1(_04380_ ), .A2(_04382_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04383_ ) );
MUX2_X1 _12039_ ( .A(\myreg.Reg[8][4] ), .B(\myreg.Reg[9][4] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04384_ ) );
MUX2_X1 _12040_ ( .A(\myreg.Reg[10][4] ), .B(\myreg.Reg[11][4] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04385_ ) );
MUX2_X1 _12041_ ( .A(_04384_ ), .B(_04385_ ), .S(fanout_net_41 ), .Z(_04386_ ) );
OAI211_X1 _12042_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04383_ ), .C1(_04386_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04387_ ) );
OAI211_X1 _12043_ ( .A(_04378_ ), .B(_04387_ ), .C1(_03649_ ), .C2(_03644_ ), .ZN(_04388_ ) );
NAND2_X1 _12044_ ( .A1(_04369_ ), .A2(_04388_ ), .ZN(_04389_ ) );
XOR2_X1 _12045_ ( .A(_02855_ ), .B(_04389_ ), .Z(_04390_ ) );
OR2_X1 _12046_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04391_ ) );
OAI211_X1 _12047_ ( .A(_04391_ ), .B(_03610_ ), .C1(_03663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04392_ ) );
OR2_X1 _12048_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04393_ ) );
OAI211_X1 _12049_ ( .A(_04393_ ), .B(fanout_net_41 ), .C1(_03663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04394_ ) );
NAND3_X1 _12050_ ( .A1(_04392_ ), .A2(_04394_ ), .A3(_03619_ ), .ZN(_04395_ ) );
MUX2_X1 _12051_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04396_ ) );
MUX2_X1 _12052_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04397_ ) );
MUX2_X1 _12053_ ( .A(_04396_ ), .B(_04397_ ), .S(_03705_ ), .Z(_04398_ ) );
OAI211_X1 _12054_ ( .A(_03606_ ), .B(_04395_ ), .C1(_04398_ ), .C2(_03708_ ), .ZN(_04399_ ) );
OR2_X1 _12055_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04400_ ) );
OAI211_X1 _12056_ ( .A(_04400_ ), .B(fanout_net_41 ), .C1(_03663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04401_ ) );
OR2_X1 _12057_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04402_ ) );
OAI211_X1 _12058_ ( .A(_04402_ ), .B(_03705_ ), .C1(_03699_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04403_ ) );
NAND3_X1 _12059_ ( .A1(_04401_ ), .A2(_04403_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04404_ ) );
MUX2_X1 _12060_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04405_ ) );
MUX2_X1 _12061_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04406_ ) );
MUX2_X1 _12062_ ( .A(_04405_ ), .B(_04406_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04407_ ) );
OAI211_X1 _12063_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04404_ ), .C1(_04407_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04408_ ) );
AOI21_X1 _12064_ ( .A(_03941_ ), .B1(_04399_ ), .B2(_04408_ ), .ZN(_04409_ ) );
AND2_X1 _12065_ ( .A1(_03941_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04410_ ) );
NOR2_X2 _12066_ ( .A1(_04409_ ), .A2(_04410_ ), .ZN(_04411_ ) );
XNOR2_X1 _12067_ ( .A(_04411_ ), .B(_02833_ ), .ZN(_04412_ ) );
AND2_X1 _12068_ ( .A1(_04390_ ), .A2(_04412_ ), .ZN(_04413_ ) );
AND4_X1 _12069_ ( .A1(_04224_ ), .A2(_04321_ ), .A3(_04368_ ), .A4(_04413_ ), .ZN(_04414_ ) );
AND3_X1 _12070_ ( .A1(_04034_ ), .A2(_04130_ ), .A3(_04414_ ), .ZN(_04415_ ) );
AND2_X1 _12071_ ( .A1(fanout_net_5 ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04416_ ) );
INV_X1 _12072_ ( .A(\ID_EX_typ [1] ), .ZN(_04417_ ) );
AND2_X1 _12073_ ( .A1(_04416_ ), .A2(_04417_ ), .ZN(_04418_ ) );
BUF_X4 _12074_ ( .A(_04418_ ), .Z(_04419_ ) );
INV_X1 _12075_ ( .A(_04419_ ), .ZN(_04420_ ) );
AND3_X1 _12076_ ( .A1(_04155_ ), .A2(_03118_ ), .A3(_04176_ ), .ZN(_04421_ ) );
AND2_X1 _12077_ ( .A1(_04179_ ), .A2(_04200_ ), .ZN(_04422_ ) );
AND2_X1 _12078_ ( .A1(_04222_ ), .A2(_03070_ ), .ZN(_04423_ ) );
AOI21_X1 _12079_ ( .A(_04422_ ), .B1(_04201_ ), .B2(_04423_ ), .ZN(_04424_ ) );
INV_X1 _12080_ ( .A(_04424_ ), .ZN(_04425_ ) );
NAND2_X1 _12081_ ( .A1(_04425_ ), .A2(_04178_ ), .ZN(_04426_ ) );
AND2_X1 _12082_ ( .A1(_04319_ ), .A2(_02938_ ), .ZN(_04427_ ) );
AND2_X1 _12083_ ( .A1(_04298_ ), .A2(_04427_ ), .ZN(_04428_ ) );
AOI21_X1 _12084_ ( .A(_04428_ ), .B1(_02963_ ), .B2(_04296_ ), .ZN(_04429_ ) );
INV_X1 _12085_ ( .A(_04429_ ), .ZN(_04430_ ) );
AND2_X1 _12086_ ( .A1(_04430_ ), .A2(_04273_ ), .ZN(_04431_ ) );
AND3_X1 _12087_ ( .A1(_04248_ ), .A2(_04244_ ), .A3(_04246_ ), .ZN(_04432_ ) );
AND3_X1 _12088_ ( .A1(_04250_ ), .A2(_03012_ ), .A3(_04271_ ), .ZN(_04433_ ) );
NOR3_X4 _12089_ ( .A1(_04431_ ), .A2(_04432_ ), .A3(_04433_ ), .ZN(_04434_ ) );
INV_X1 _12090_ ( .A(_04224_ ), .ZN(_04435_ ) );
OAI21_X1 _12091_ ( .A(_04426_ ), .B1(_04434_ ), .B2(_04435_ ), .ZN(_04436_ ) );
AOI211_X1 _12092_ ( .A(_04421_ ), .B(_04436_ ), .C1(_03094_ ), .C2(_04153_ ), .ZN(_04437_ ) );
AND2_X1 _12093_ ( .A1(_04057_ ), .A2(_04082_ ), .ZN(_04438_ ) );
AOI21_X1 _12094_ ( .A(_04438_ ), .B1(_02779_ ), .B2(_04056_ ), .ZN(_04439_ ) );
INV_X1 _12095_ ( .A(_04107_ ), .ZN(_04440_ ) );
INV_X1 _12096_ ( .A(_04129_ ), .ZN(_04441_ ) );
NOR3_X1 _12097_ ( .A1(_04439_ ), .A2(_04440_ ), .A3(_04441_ ), .ZN(_04442_ ) );
AND2_X1 _12098_ ( .A1(_04128_ ), .A2(_02755_ ), .ZN(_04443_ ) );
NAND2_X1 _12099_ ( .A1(_04107_ ), .A2(_04443_ ), .ZN(_04444_ ) );
OAI21_X1 _12100_ ( .A(_04444_ ), .B1(_02810_ ), .B2(_04106_ ), .ZN(_04445_ ) );
OAI211_X1 _12101_ ( .A(_04368_ ), .B(_04413_ ), .C1(_04442_ ), .C2(_04445_ ), .ZN(_04446_ ) );
AND3_X1 _12102_ ( .A1(_04343_ ), .A2(_02908_ ), .A3(_04364_ ), .ZN(_04447_ ) );
AND2_X1 _12103_ ( .A1(_02855_ ), .A2(_04389_ ), .ZN(_04448_ ) );
NAND2_X1 _12104_ ( .A1(_04412_ ), .A2(_04448_ ), .ZN(_04449_ ) );
INV_X1 _12105_ ( .A(_02833_ ), .ZN(_04450_ ) );
OAI21_X1 _12106_ ( .A(_04449_ ), .B1(_04450_ ), .B2(_04411_ ), .ZN(_04451_ ) );
AOI221_X1 _12107_ ( .A(_04447_ ), .B1(_02886_ ), .B2(_04342_ ), .C1(_04368_ ), .C2(_04451_ ), .ZN(_04452_ ) );
AND2_X1 _12108_ ( .A1(_04446_ ), .A2(_04452_ ), .ZN(_04453_ ) );
INV_X2 _12109_ ( .A(_04453_ ), .ZN(_04454_ ) );
NAND3_X1 _12110_ ( .A1(_04454_ ), .A2(_04224_ ), .A3(_04321_ ), .ZN(_04455_ ) );
AND2_X1 _12111_ ( .A1(_04437_ ), .A2(_04455_ ), .ZN(_04456_ ) );
INV_X2 _12112_ ( .A(_04456_ ), .ZN(_04457_ ) );
AND2_X4 _12113_ ( .A1(_04457_ ), .A2(_03841_ ), .ZN(_04458_ ) );
NAND3_X1 _12114_ ( .A1(_03657_ ), .A2(_02626_ ), .A3(_03692_ ), .ZN(_04459_ ) );
INV_X1 _12115_ ( .A(_03655_ ), .ZN(_04460_ ) );
OAI21_X1 _12116_ ( .A(_04459_ ), .B1(_03656_ ), .B2(_04460_ ), .ZN(_04461_ ) );
NOR2_X1 _12117_ ( .A1(_03721_ ), .A2(_02682_ ), .ZN(_04462_ ) );
AND2_X1 _12118_ ( .A1(_03721_ ), .A2(_02682_ ), .ZN(_04463_ ) );
INV_X1 _12119_ ( .A(_04463_ ), .ZN(_04464_ ) );
NAND2_X1 _12120_ ( .A1(_03746_ ), .A2(_02706_ ), .ZN(_04465_ ) );
AOI21_X1 _12121_ ( .A(_04462_ ), .B1(_04464_ ), .B2(_04465_ ), .ZN(_04466_ ) );
AOI21_X1 _12122_ ( .A(_04461_ ), .B1(_04466_ ), .B2(_03694_ ), .ZN(_04467_ ) );
INV_X1 _12123_ ( .A(_03840_ ), .ZN(_04468_ ) );
NOR2_X1 _12124_ ( .A1(_04467_ ), .A2(_04468_ ), .ZN(_04469_ ) );
AND2_X1 _12125_ ( .A1(_03817_ ), .A2(_03839_ ), .ZN(_04470_ ) );
INV_X1 _12126_ ( .A(_04470_ ), .ZN(_04471_ ) );
INV_X1 _12127_ ( .A(_03792_ ), .ZN(_04472_ ) );
AND2_X1 _12128_ ( .A1(_03769_ ), .A2(_02598_ ), .ZN(_04473_ ) );
NAND2_X1 _12129_ ( .A1(_03794_ ), .A2(_04473_ ), .ZN(_04474_ ) );
AOI21_X1 _12130_ ( .A(_04471_ ), .B1(_04472_ ), .B2(_04474_ ), .ZN(_04475_ ) );
OR2_X1 _12131_ ( .A1(_04469_ ), .A2(_04475_ ), .ZN(_04476_ ) );
AND2_X1 _12132_ ( .A1(_02548_ ), .A2(_03816_ ), .ZN(_04477_ ) );
AND2_X1 _12133_ ( .A1(_02522_ ), .A2(_03838_ ), .ZN(_04478_ ) );
AND2_X1 _12134_ ( .A1(_03817_ ), .A2(_04478_ ), .ZN(_04479_ ) );
NOR3_X1 _12135_ ( .A1(_04476_ ), .A2(_04477_ ), .A3(_04479_ ), .ZN(_04480_ ) );
INV_X1 _12136_ ( .A(_04480_ ), .ZN(_04481_ ) );
OAI211_X4 _12137_ ( .A(_03940_ ), .B(_04033_ ), .C1(_04458_ ), .C2(_04481_ ), .ZN(_04482_ ) );
INV_X1 _12138_ ( .A(_03172_ ), .ZN(_04483_ ) );
NOR2_X1 _12139_ ( .A1(_04483_ ), .A2(_03961_ ), .ZN(_04484_ ) );
AOI21_X1 _12140_ ( .A(_03984_ ), .B1(_03178_ ), .B2(_03197_ ), .ZN(_04485_ ) );
NOR2_X1 _12141_ ( .A1(_04484_ ), .A2(_04485_ ), .ZN(_04486_ ) );
NAND2_X1 _12142_ ( .A1(_04010_ ), .A2(_04032_ ), .ZN(_04487_ ) );
INV_X1 _12143_ ( .A(_03198_ ), .ZN(_04488_ ) );
AOI211_X1 _12144_ ( .A(_04486_ ), .B(_04487_ ), .C1(_04488_ ), .C2(_03984_ ), .ZN(_04489_ ) );
INV_X1 _12145_ ( .A(_03987_ ), .ZN(_04490_ ) );
NOR2_X1 _12146_ ( .A1(_04490_ ), .A2(_04009_ ), .ZN(_04491_ ) );
NOR2_X1 _12147_ ( .A1(_03227_ ), .A2(_04031_ ), .ZN(_04492_ ) );
AND2_X1 _12148_ ( .A1(_04010_ ), .A2(_04492_ ), .ZN(_04493_ ) );
NOR3_X1 _12149_ ( .A1(_04489_ ), .A2(_04491_ ), .A3(_04493_ ), .ZN(_04494_ ) );
INV_X1 _12150_ ( .A(_03940_ ), .ZN(_04495_ ) );
NOR2_X1 _12151_ ( .A1(_04494_ ), .A2(_04495_ ), .ZN(_04496_ ) );
INV_X1 _12152_ ( .A(_04496_ ), .ZN(_04497_ ) );
NAND4_X1 _12153_ ( .A1(_03892_ ), .A2(_03253_ ), .A3(_03868_ ), .A4(_03844_ ), .ZN(_04498_ ) );
OAI21_X1 _12154_ ( .A(_04498_ ), .B1(_03282_ ), .B2(_03891_ ), .ZN(_04499_ ) );
AND3_X1 _12155_ ( .A1(_04499_ ), .A2(_03917_ ), .A3(_03939_ ), .ZN(_04500_ ) );
INV_X1 _12156_ ( .A(_04500_ ), .ZN(_04501_ ) );
AOI21_X1 _12157_ ( .A(_03916_ ), .B1(_03335_ ), .B2(_03316_ ), .ZN(_04502_ ) );
NOR2_X1 _12158_ ( .A1(_03310_ ), .A2(_03937_ ), .ZN(_04503_ ) );
AOI21_X1 _12159_ ( .A(_04502_ ), .B1(_04503_ ), .B2(_03917_ ), .ZN(_04504_ ) );
AND3_X1 _12160_ ( .A1(_04497_ ), .A2(_04501_ ), .A3(_04504_ ), .ZN(_04505_ ) );
AND2_X1 _12161_ ( .A1(_04416_ ), .A2(\ID_EX_typ [1] ), .ZN(_04506_ ) );
AND3_X1 _12162_ ( .A1(_04482_ ), .A2(_04505_ ), .A3(_04506_ ), .ZN(_04507_ ) );
INV_X1 _12163_ ( .A(fanout_net_7 ), .ZN(_04508_ ) );
BUF_X4 _12164_ ( .A(_04508_ ), .Z(_04509_ ) );
BUF_X4 _12165_ ( .A(_04509_ ), .Z(_04510_ ) );
BUF_X2 _12166_ ( .A(_04510_ ), .Z(_04511_ ) );
NAND3_X1 _12167_ ( .A1(_03918_ ), .A2(_04511_ ), .A3(_03936_ ), .ZN(_04512_ ) );
NAND2_X1 _12168_ ( .A1(fanout_net_7 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04513_ ) );
AND2_X1 _12169_ ( .A1(_04512_ ), .A2(_04513_ ), .ZN(_04514_ ) );
XNOR2_X1 _12170_ ( .A(_03309_ ), .B(_04514_ ), .ZN(_04515_ ) );
NAND2_X1 _12171_ ( .A1(_03916_ ), .A2(_04511_ ), .ZN(_04516_ ) );
OR2_X1 _12172_ ( .A1(_04511_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04517_ ) );
AND3_X1 _12173_ ( .A1(_04516_ ), .A2(_03336_ ), .A3(_04517_ ), .ZN(_04518_ ) );
AOI21_X1 _12174_ ( .A(_03336_ ), .B1(_04516_ ), .B2(_04517_ ), .ZN(_04519_ ) );
NOR2_X1 _12175_ ( .A1(_04518_ ), .A2(_04519_ ), .ZN(_04520_ ) );
INV_X1 _12176_ ( .A(_04520_ ), .ZN(_04521_ ) );
NAND3_X1 _12177_ ( .A1(_03871_ ), .A2(_04510_ ), .A3(_03890_ ), .ZN(_04522_ ) );
NAND2_X1 _12178_ ( .A1(fanout_net_7 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04523_ ) );
AND2_X2 _12179_ ( .A1(_04522_ ), .A2(_04523_ ), .ZN(_04524_ ) );
XNOR2_X1 _12180_ ( .A(_04524_ ), .B(_03282_ ), .ZN(_04525_ ) );
NOR3_X1 _12181_ ( .A1(_04515_ ), .A2(_04521_ ), .A3(_04525_ ), .ZN(_04526_ ) );
NAND3_X1 _12182_ ( .A1(_03844_ ), .A2(_04511_ ), .A3(_03868_ ), .ZN(_04527_ ) );
NAND2_X1 _12183_ ( .A1(fanout_net_7 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04528_ ) );
AND2_X2 _12184_ ( .A1(_04527_ ), .A2(_04528_ ), .ZN(_04529_ ) );
XOR2_X1 _12185_ ( .A(_03253_ ), .B(_04529_ ), .Z(_04530_ ) );
INV_X1 _12186_ ( .A(_04530_ ), .ZN(_04531_ ) );
NAND2_X1 _12187_ ( .A1(_04526_ ), .A2(_04531_ ), .ZN(_04532_ ) );
NAND3_X1 _12188_ ( .A1(_03818_ ), .A2(_03837_ ), .A3(_04510_ ), .ZN(_04533_ ) );
NAND2_X1 _12189_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [22] ), .ZN(_04534_ ) );
AND2_X2 _12190_ ( .A1(_04533_ ), .A2(_04534_ ), .ZN(_04535_ ) );
XNOR2_X1 _12191_ ( .A(_04535_ ), .B(_02521_ ), .ZN(_04536_ ) );
NAND3_X1 _12192_ ( .A1(_03796_ ), .A2(_04510_ ), .A3(_03815_ ), .ZN(_04537_ ) );
NAND2_X1 _12193_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [23] ), .ZN(_04538_ ) );
AND2_X1 _12194_ ( .A1(_04537_ ), .A2(_04538_ ), .ZN(_04539_ ) );
XNOR2_X1 _12195_ ( .A(_04539_ ), .B(_02547_ ), .ZN(_04540_ ) );
NOR2_X1 _12196_ ( .A1(_04536_ ), .A2(_04540_ ), .ZN(_04541_ ) );
INV_X1 _12197_ ( .A(_04541_ ), .ZN(_04542_ ) );
NAND3_X1 _12198_ ( .A1(_03771_ ), .A2(_04510_ ), .A3(_03790_ ), .ZN(_04543_ ) );
NAND2_X1 _12199_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [21] ), .ZN(_04544_ ) );
AND2_X1 _12200_ ( .A1(_04543_ ), .A2(_04544_ ), .ZN(_04545_ ) );
XNOR2_X1 _12201_ ( .A(_04545_ ), .B(_02575_ ), .ZN(_04546_ ) );
NAND2_X1 _12202_ ( .A1(_03769_ ), .A2(_04510_ ), .ZN(_04547_ ) );
NAND2_X1 _12203_ ( .A1(_02599_ ), .A2(fanout_net_7 ), .ZN(_04548_ ) );
NAND2_X2 _12204_ ( .A1(_04547_ ), .A2(_04548_ ), .ZN(_04549_ ) );
XNOR2_X1 _12205_ ( .A(_04549_ ), .B(_02598_ ), .ZN(_04550_ ) );
NOR3_X4 _12206_ ( .A1(_04542_ ), .A2(_04546_ ), .A3(_04550_ ), .ZN(_04551_ ) );
NAND3_X1 _12207_ ( .A1(_03660_ ), .A2(_04510_ ), .A3(_03691_ ), .ZN(_04552_ ) );
NAND2_X1 _12208_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [18] ), .ZN(_04553_ ) );
AND2_X2 _12209_ ( .A1(_04552_ ), .A2(_04553_ ), .ZN(_04554_ ) );
XNOR2_X1 _12210_ ( .A(_04554_ ), .B(_02626_ ), .ZN(_04555_ ) );
OR2_X1 _12211_ ( .A1(_03655_ ), .A2(fanout_net_7 ), .ZN(_04556_ ) );
NAND2_X1 _12212_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [19] ), .ZN(_04557_ ) );
AND2_X1 _12213_ ( .A1(_04556_ ), .A2(_04557_ ), .ZN(_04558_ ) );
NOR2_X1 _12214_ ( .A1(_04558_ ), .A2(_03656_ ), .ZN(_04559_ ) );
INV_X1 _12215_ ( .A(_04559_ ), .ZN(_04560_ ) );
AND3_X1 _12216_ ( .A1(_04556_ ), .A2(_03656_ ), .A3(_04557_ ), .ZN(_04561_ ) );
INV_X1 _12217_ ( .A(_04561_ ), .ZN(_04562_ ) );
AOI21_X1 _12218_ ( .A(_04555_ ), .B1(_04560_ ), .B2(_04562_ ), .ZN(_04563_ ) );
NAND2_X1 _12219_ ( .A1(_04551_ ), .A2(_04563_ ), .ZN(_04564_ ) );
NAND3_X1 _12220_ ( .A1(_03719_ ), .A2(_03720_ ), .A3(_04509_ ), .ZN(_04565_ ) );
NAND2_X1 _12221_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [17] ), .ZN(_04566_ ) );
AND2_X2 _12222_ ( .A1(_04565_ ), .A2(_04566_ ), .ZN(_04567_ ) );
XNOR2_X1 _12223_ ( .A(_04567_ ), .B(_02682_ ), .ZN(_04568_ ) );
NAND3_X1 _12224_ ( .A1(_03723_ ), .A2(_04510_ ), .A3(_03745_ ), .ZN(_04569_ ) );
NAND2_X1 _12225_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [16] ), .ZN(_04570_ ) );
AND2_X2 _12226_ ( .A1(_04569_ ), .A2(_04570_ ), .ZN(_04571_ ) );
INV_X1 _12227_ ( .A(_02706_ ), .ZN(_04572_ ) );
NOR2_X1 _12228_ ( .A1(_04571_ ), .A2(_04572_ ), .ZN(_04573_ ) );
AND3_X1 _12229_ ( .A1(_04572_ ), .A2(_04570_ ), .A3(_04569_ ), .ZN(_04574_ ) );
NOR2_X1 _12230_ ( .A1(_04573_ ), .A2(_04574_ ), .ZN(_04575_ ) );
NOR3_X1 _12231_ ( .A1(_04564_ ), .A2(_04568_ ), .A3(_04575_ ), .ZN(_04576_ ) );
NAND3_X1 _12232_ ( .A1(_04299_ ), .A2(_04318_ ), .A3(_04510_ ), .ZN(_04577_ ) );
NAND2_X1 _12233_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [8] ), .ZN(_04578_ ) );
AND2_X2 _12234_ ( .A1(_04577_ ), .A2(_04578_ ), .ZN(_04579_ ) );
XNOR2_X1 _12235_ ( .A(_04579_ ), .B(_02938_ ), .ZN(_04580_ ) );
INV_X1 _12236_ ( .A(_04580_ ), .ZN(_04581_ ) );
NAND3_X1 _12237_ ( .A1(_04293_ ), .A2(_04509_ ), .A3(_04295_ ), .ZN(_04582_ ) );
NAND2_X1 _12238_ ( .A1(_02964_ ), .A2(fanout_net_7 ), .ZN(_04583_ ) );
NAND2_X1 _12239_ ( .A1(_04582_ ), .A2(_04583_ ), .ZN(_04584_ ) );
XNOR2_X1 _12240_ ( .A(_04584_ ), .B(_02963_ ), .ZN(_04585_ ) );
INV_X1 _12241_ ( .A(_04585_ ), .ZN(_04586_ ) );
NAND2_X1 _12242_ ( .A1(_04581_ ), .A2(_04586_ ), .ZN(_04587_ ) );
OR2_X1 _12243_ ( .A1(_04153_ ), .A2(fanout_net_7 ), .ZN(_04588_ ) );
NAND2_X1 _12244_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [15] ), .ZN(_04589_ ) );
AND2_X1 _12245_ ( .A1(_04588_ ), .A2(_04589_ ), .ZN(_04590_ ) );
NOR2_X1 _12246_ ( .A1(_04590_ ), .A2(_04154_ ), .ZN(_04591_ ) );
AND3_X1 _12247_ ( .A1(_04588_ ), .A2(_04154_ ), .A3(_04589_ ), .ZN(_04592_ ) );
NOR2_X2 _12248_ ( .A1(_04591_ ), .A2(_04592_ ), .ZN(_04593_ ) );
NAND3_X1 _12249_ ( .A1(_04156_ ), .A2(_04175_ ), .A3(_04509_ ), .ZN(_04594_ ) );
NAND2_X1 _12250_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [14] ), .ZN(_04595_ ) );
AND2_X2 _12251_ ( .A1(_04594_ ), .A2(_04595_ ), .ZN(_04596_ ) );
XNOR2_X1 _12252_ ( .A(_04596_ ), .B(_03118_ ), .ZN(_04597_ ) );
NOR2_X1 _12253_ ( .A1(_04593_ ), .A2(_04597_ ), .ZN(_04598_ ) );
NAND3_X1 _12254_ ( .A1(_04202_ ), .A2(_04509_ ), .A3(_04221_ ), .ZN(_04599_ ) );
NAND2_X1 _12255_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [12] ), .ZN(_04600_ ) );
AND2_X2 _12256_ ( .A1(_04599_ ), .A2(_04600_ ), .ZN(_04601_ ) );
XNOR2_X1 _12257_ ( .A(_04601_ ), .B(_03070_ ), .ZN(_04602_ ) );
INV_X1 _12258_ ( .A(_04602_ ), .ZN(_04603_ ) );
NAND3_X1 _12259_ ( .A1(_04180_ ), .A2(_04509_ ), .A3(_04199_ ), .ZN(_04604_ ) );
NAND2_X1 _12260_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [13] ), .ZN(_04605_ ) );
AND2_X1 _12261_ ( .A1(_04604_ ), .A2(_04605_ ), .ZN(_04606_ ) );
XNOR2_X1 _12262_ ( .A(_04606_ ), .B(_04179_ ), .ZN(_04607_ ) );
INV_X1 _12263_ ( .A(_04607_ ), .ZN(_04608_ ) );
AND3_X1 _12264_ ( .A1(_04598_ ), .A2(_04603_ ), .A3(_04608_ ), .ZN(_04609_ ) );
OR2_X1 _12265_ ( .A1(_04247_ ), .A2(fanout_net_7 ), .ZN(_04610_ ) );
NAND2_X1 _12266_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [11] ), .ZN(_04611_ ) );
AND2_X1 _12267_ ( .A1(_04610_ ), .A2(_04611_ ), .ZN(_04612_ ) );
NOR2_X1 _12268_ ( .A1(_04612_ ), .A2(_04249_ ), .ZN(_04613_ ) );
AND3_X1 _12269_ ( .A1(_04610_ ), .A2(_04249_ ), .A3(_04611_ ), .ZN(_04614_ ) );
NOR2_X2 _12270_ ( .A1(_04613_ ), .A2(_04614_ ), .ZN(_04615_ ) );
INV_X1 _12271_ ( .A(_04615_ ), .ZN(_04616_ ) );
NAND3_X1 _12272_ ( .A1(_04251_ ), .A2(_04509_ ), .A3(_04270_ ), .ZN(_04617_ ) );
NAND2_X1 _12273_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [10] ), .ZN(_04618_ ) );
AND2_X2 _12274_ ( .A1(_04617_ ), .A2(_04618_ ), .ZN(_04619_ ) );
XNOR2_X1 _12275_ ( .A(_04619_ ), .B(_03012_ ), .ZN(_04620_ ) );
INV_X1 _12276_ ( .A(_04620_ ), .ZN(_04621_ ) );
NAND3_X1 _12277_ ( .A1(_04609_ ), .A2(_04616_ ), .A3(_04621_ ), .ZN(_04622_ ) );
NAND2_X1 _12278_ ( .A1(_04411_ ), .A2(_04509_ ), .ZN(_04623_ ) );
NAND2_X1 _12279_ ( .A1(_02862_ ), .A2(fanout_net_7 ), .ZN(_04624_ ) );
NAND2_X2 _12280_ ( .A1(_04623_ ), .A2(_04624_ ), .ZN(_04625_ ) );
XNOR2_X1 _12281_ ( .A(_04625_ ), .B(_04450_ ), .ZN(_04626_ ) );
NAND3_X1 _12282_ ( .A1(_04369_ ), .A2(_04509_ ), .A3(_04388_ ), .ZN(_04627_ ) );
NAND2_X1 _12283_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [4] ), .ZN(_04628_ ) );
AND2_X2 _12284_ ( .A1(_04627_ ), .A2(_04628_ ), .ZN(_04629_ ) );
INV_X1 _12285_ ( .A(_04629_ ), .ZN(_04630_ ) );
NOR3_X1 _12286_ ( .A1(_04626_ ), .A2(_02860_ ), .A3(_04630_ ), .ZN(_04631_ ) );
XNOR2_X1 _12287_ ( .A(_04629_ ), .B(_02855_ ), .ZN(_04632_ ) );
OR2_X1 _12288_ ( .A1(_04106_ ), .A2(fanout_net_7 ), .ZN(_04633_ ) );
NAND2_X1 _12289_ ( .A1(fanout_net_7 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_04634_ ) );
AND2_X2 _12290_ ( .A1(_04633_ ), .A2(_04634_ ), .ZN(_04635_ ) );
XNOR2_X1 _12291_ ( .A(_04635_ ), .B(_02810_ ), .ZN(_04636_ ) );
NAND3_X1 _12292_ ( .A1(_04126_ ), .A2(_04127_ ), .A3(_04508_ ), .ZN(_04637_ ) );
NAND2_X1 _12293_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [2] ), .ZN(_04638_ ) );
AND2_X2 _12294_ ( .A1(_04637_ ), .A2(_04638_ ), .ZN(_04639_ ) );
BUF_X4 _12295_ ( .A(_04639_ ), .Z(_04640_ ) );
INV_X2 _12296_ ( .A(_04640_ ), .ZN(_04641_ ) );
NOR3_X1 _12297_ ( .A1(_04636_ ), .A2(_04108_ ), .A3(_04641_ ), .ZN(_04642_ ) );
INV_X1 _12298_ ( .A(_04635_ ), .ZN(_04643_ ) );
AOI21_X1 _12299_ ( .A(_04642_ ), .B1(_02732_ ), .B2(_04643_ ), .ZN(_04644_ ) );
NAND2_X2 _12300_ ( .A1(_04056_ ), .A2(_04508_ ), .ZN(_04645_ ) );
NAND2_X1 _12301_ ( .A1(_02780_ ), .A2(fanout_net_7 ), .ZN(_04646_ ) );
NAND2_X4 _12302_ ( .A1(_04645_ ), .A2(_04646_ ), .ZN(_04647_ ) );
NAND2_X1 _12303_ ( .A1(_04647_ ), .A2(_02779_ ), .ZN(_04648_ ) );
XNOR2_X2 _12304_ ( .A(_04647_ ), .B(_02779_ ), .ZN(_04649_ ) );
INV_X1 _12305_ ( .A(_04058_ ), .ZN(_04650_ ) );
NAND3_X1 _12306_ ( .A1(_04078_ ), .A2(_04508_ ), .A3(_04080_ ), .ZN(_04651_ ) );
NAND2_X1 _12307_ ( .A1(_02782_ ), .A2(fanout_net_7 ), .ZN(_04652_ ) );
AND3_X1 _12308_ ( .A1(_04650_ ), .A2(_04651_ ), .A3(_04652_ ), .ZN(_04653_ ) );
OAI21_X1 _12309_ ( .A(_04648_ ), .B1(_04649_ ), .B2(_04653_ ), .ZN(_04654_ ) );
XNOR2_X1 _12310_ ( .A(_04639_ ), .B(_02755_ ), .ZN(_04655_ ) );
INV_X1 _12311_ ( .A(_04655_ ), .ZN(_04656_ ) );
AND2_X1 _12312_ ( .A1(_04635_ ), .A2(_02732_ ), .ZN(_04657_ ) );
NOR2_X1 _12313_ ( .A1(_04635_ ), .A2(_02732_ ), .ZN(_04658_ ) );
OAI211_X1 _12314_ ( .A(_04654_ ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_04659_ ) );
AOI211_X1 _12315_ ( .A(_04626_ ), .B(_04632_ ), .C1(_04644_ ), .C2(_04659_ ), .ZN(_04660_ ) );
INV_X1 _12316_ ( .A(_04625_ ), .ZN(_04661_ ) );
AOI211_X1 _12317_ ( .A(_04631_ ), .B(_04660_ ), .C1(_02833_ ), .C2(_04661_ ), .ZN(_04662_ ) );
NAND2_X1 _12318_ ( .A1(_04342_ ), .A2(_04508_ ), .ZN(_04663_ ) );
OR2_X1 _12319_ ( .A1(_04508_ ), .A2(\ID_EX_imm [7] ), .ZN(_04664_ ) );
NAND2_X1 _12320_ ( .A1(_04663_ ), .A2(_04664_ ), .ZN(_04665_ ) );
XNOR2_X2 _12321_ ( .A(_04665_ ), .B(_02886_ ), .ZN(_04666_ ) );
NAND2_X1 _12322_ ( .A1(_04364_ ), .A2(_04509_ ), .ZN(_04667_ ) );
OR2_X1 _12323_ ( .A1(_04508_ ), .A2(\ID_EX_imm [6] ), .ZN(_04668_ ) );
NAND2_X1 _12324_ ( .A1(_04667_ ), .A2(_04668_ ), .ZN(_04669_ ) );
XNOR2_X1 _12325_ ( .A(_04669_ ), .B(_02908_ ), .ZN(_04670_ ) );
OR3_X2 _12326_ ( .A1(_04662_ ), .A2(_04666_ ), .A3(_04670_ ), .ZN(_04671_ ) );
INV_X1 _12327_ ( .A(_04666_ ), .ZN(_04672_ ) );
AND3_X1 _12328_ ( .A1(_04672_ ), .A2(_02908_ ), .A3(_04669_ ), .ZN(_04673_ ) );
AOI21_X1 _12329_ ( .A(_04673_ ), .B1(_02886_ ), .B2(_04665_ ), .ZN(_04674_ ) );
AOI211_X2 _12330_ ( .A(_04587_ ), .B(_04622_ ), .C1(_04671_ ), .C2(_04674_ ), .ZN(_04675_ ) );
NAND3_X1 _12331_ ( .A1(_04616_ ), .A2(_03012_ ), .A3(_04619_ ), .ZN(_04676_ ) );
INV_X1 _12332_ ( .A(_04612_ ), .ZN(_04677_ ) );
OAI21_X1 _12333_ ( .A(_04621_ ), .B1(_04613_ ), .B2(_04614_ ), .ZN(_04678_ ) );
INV_X1 _12334_ ( .A(_02938_ ), .ZN(_04679_ ) );
INV_X1 _12335_ ( .A(_04579_ ), .ZN(_04680_ ) );
NOR3_X1 _12336_ ( .A1(_04585_ ), .A2(_04679_ ), .A3(_04680_ ), .ZN(_04681_ ) );
AOI21_X1 _12337_ ( .A(_04681_ ), .B1(_02963_ ), .B2(_04584_ ), .ZN(_04682_ ) );
OAI221_X1 _12338_ ( .A(_04676_ ), .B1(_04249_ ), .B2(_04677_ ), .C1(_04678_ ), .C2(_04682_ ), .ZN(_04683_ ) );
AND2_X1 _12339_ ( .A1(_04683_ ), .A2(_04609_ ), .ZN(_04684_ ) );
INV_X1 _12340_ ( .A(_03118_ ), .ZN(_04685_ ) );
INV_X1 _12341_ ( .A(_04596_ ), .ZN(_04686_ ) );
NOR3_X1 _12342_ ( .A1(_04593_ ), .A2(_04685_ ), .A3(_04686_ ), .ZN(_04687_ ) );
AND3_X1 _12343_ ( .A1(_04179_ ), .A2(_04605_ ), .A3(_04604_ ), .ZN(_04688_ ) );
AND3_X1 _12344_ ( .A1(_04608_ ), .A2(_03070_ ), .A3(_04601_ ), .ZN(_04689_ ) );
OAI21_X1 _12345_ ( .A(_04598_ ), .B1(_04688_ ), .B2(_04689_ ), .ZN(_04690_ ) );
INV_X1 _12346_ ( .A(_04590_ ), .ZN(_04691_ ) );
OAI21_X1 _12347_ ( .A(_04690_ ), .B1(_04154_ ), .B2(_04691_ ), .ZN(_04692_ ) );
OR3_X4 _12348_ ( .A1(_04684_ ), .A2(_04687_ ), .A3(_04692_ ), .ZN(_04693_ ) );
OAI21_X1 _12349_ ( .A(_04576_ ), .B1(_04675_ ), .B2(_04693_ ), .ZN(_04694_ ) );
INV_X1 _12350_ ( .A(_04540_ ), .ZN(_04695_ ) );
NAND3_X1 _12351_ ( .A1(_04695_ ), .A2(_02522_ ), .A3(_04535_ ), .ZN(_04696_ ) );
INV_X1 _12352_ ( .A(_04545_ ), .ZN(_04697_ ) );
AND2_X1 _12353_ ( .A1(_04697_ ), .A2(_02575_ ), .ZN(_04698_ ) );
NOR2_X1 _12354_ ( .A1(_04697_ ), .A2(_02575_ ), .ZN(_04699_ ) );
OAI211_X1 _12355_ ( .A(_02598_ ), .B(_04549_ ), .C1(_04698_ ), .C2(_04699_ ), .ZN(_04700_ ) );
NAND3_X1 _12356_ ( .A1(_04543_ ), .A2(_02575_ ), .A3(_04544_ ), .ZN(_04701_ ) );
AOI21_X1 _12357_ ( .A(_04542_ ), .B1(_04700_ ), .B2(_04701_ ), .ZN(_04702_ ) );
NOR2_X2 _12358_ ( .A1(_04559_ ), .A2(_04561_ ), .ZN(_04703_ ) );
INV_X1 _12359_ ( .A(_04703_ ), .ZN(_04704_ ) );
NAND3_X1 _12360_ ( .A1(_04704_ ), .A2(_02626_ ), .A3(_04554_ ), .ZN(_04705_ ) );
NAND3_X1 _12361_ ( .A1(_04556_ ), .A2(_02655_ ), .A3(_04557_ ), .ZN(_04706_ ) );
INV_X1 _12362_ ( .A(_04563_ ), .ZN(_04707_ ) );
INV_X1 _12363_ ( .A(_04568_ ), .ZN(_04708_ ) );
AND3_X1 _12364_ ( .A1(_04708_ ), .A2(_02706_ ), .A3(_04571_ ), .ZN(_04709_ ) );
AOI21_X1 _12365_ ( .A(_04709_ ), .B1(_02682_ ), .B2(_04567_ ), .ZN(_04710_ ) );
OAI211_X1 _12366_ ( .A(_04705_ ), .B(_04706_ ), .C1(_04707_ ), .C2(_04710_ ), .ZN(_04711_ ) );
AOI221_X2 _12367_ ( .A(_04702_ ), .B1(_02548_ ), .B2(_04539_ ), .C1(_04711_ ), .C2(_04551_ ), .ZN(_04712_ ) );
NAND3_X1 _12368_ ( .A1(_04694_ ), .A2(_04696_ ), .A3(_04712_ ), .ZN(_04713_ ) );
NAND3_X1 _12369_ ( .A1(_03989_ ), .A2(_04511_ ), .A3(_04008_ ), .ZN(_04714_ ) );
NAND2_X1 _12370_ ( .A1(_02484_ ), .A2(\ID_EX_typ [4] ), .ZN(_04715_ ) );
NAND2_X1 _12371_ ( .A1(_04714_ ), .A2(_04715_ ), .ZN(_04716_ ) );
XNOR2_X1 _12372_ ( .A(_03987_ ), .B(_04716_ ), .ZN(_04717_ ) );
NAND3_X1 _12373_ ( .A1(_04011_ ), .A2(_04510_ ), .A3(_04030_ ), .ZN(_04718_ ) );
INV_X1 _12374_ ( .A(\ID_EX_imm [26] ), .ZN(_04719_ ) );
NAND2_X1 _12375_ ( .A1(_04719_ ), .A2(\ID_EX_typ [4] ), .ZN(_04720_ ) );
NAND2_X1 _12376_ ( .A1(_04718_ ), .A2(_04720_ ), .ZN(_04721_ ) );
NOR2_X1 _12377_ ( .A1(_04721_ ), .A2(_03227_ ), .ZN(_04722_ ) );
AOI21_X1 _12378_ ( .A(_03221_ ), .B1(_04718_ ), .B2(_04720_ ), .ZN(_04723_ ) );
NOR2_X1 _12379_ ( .A1(_04722_ ), .A2(_04723_ ), .ZN(_04724_ ) );
NOR2_X1 _12380_ ( .A1(_04717_ ), .A2(_04724_ ), .ZN(_04725_ ) );
NAND3_X1 _12381_ ( .A1(_03942_ ), .A2(_04511_ ), .A3(_03960_ ), .ZN(_04726_ ) );
NAND2_X1 _12382_ ( .A1(_03173_ ), .A2(\ID_EX_typ [4] ), .ZN(_04727_ ) );
NAND2_X1 _12383_ ( .A1(_04726_ ), .A2(_04727_ ), .ZN(_04728_ ) );
NOR2_X1 _12384_ ( .A1(_04728_ ), .A2(_04483_ ), .ZN(_04729_ ) );
AOI21_X1 _12385_ ( .A(_03172_ ), .B1(_04726_ ), .B2(_04727_ ), .ZN(_04730_ ) );
NOR2_X1 _12386_ ( .A1(_04729_ ), .A2(_04730_ ), .ZN(_04731_ ) );
INV_X1 _12387_ ( .A(_04731_ ), .ZN(_04732_ ) );
NAND3_X1 _12388_ ( .A1(_03964_ ), .A2(_04511_ ), .A3(_03983_ ), .ZN(_04733_ ) );
NAND2_X1 _12389_ ( .A1(_03224_ ), .A2(\ID_EX_typ [4] ), .ZN(_04734_ ) );
NAND2_X1 _12390_ ( .A1(_04733_ ), .A2(_04734_ ), .ZN(_04735_ ) );
NOR2_X1 _12391_ ( .A1(_04735_ ), .A2(_04488_ ), .ZN(_04736_ ) );
AOI21_X1 _12392_ ( .A(_03198_ ), .B1(_04733_ ), .B2(_04734_ ), .ZN(_04737_ ) );
NOR2_X1 _12393_ ( .A1(_04736_ ), .A2(_04737_ ), .ZN(_04738_ ) );
INV_X1 _12394_ ( .A(_04738_ ), .ZN(_04739_ ) );
NAND4_X1 _12395_ ( .A1(_04713_ ), .A2(_04725_ ), .A3(_04732_ ), .A4(_04739_ ), .ZN(_04740_ ) );
INV_X1 _12396_ ( .A(_04728_ ), .ZN(_04741_ ) );
NOR3_X1 _12397_ ( .A1(_04738_ ), .A2(_04483_ ), .A3(_04741_ ), .ZN(_04742_ ) );
AOI22_X1 _12398_ ( .A1(_04733_ ), .A2(_04734_ ), .B1(_03178_ ), .B2(_03197_ ), .ZN(_04743_ ) );
OAI21_X1 _12399_ ( .A(_04725_ ), .B1(_04742_ ), .B2(_04743_ ), .ZN(_04744_ ) );
INV_X1 _12400_ ( .A(_04717_ ), .ZN(_04745_ ) );
NAND3_X1 _12401_ ( .A1(_04745_ ), .A2(_03221_ ), .A3(_04721_ ), .ZN(_04746_ ) );
NAND2_X1 _12402_ ( .A1(_03987_ ), .A2(_04716_ ), .ZN(_04747_ ) );
AND3_X1 _12403_ ( .A1(_04744_ ), .A2(_04746_ ), .A3(_04747_ ), .ZN(_04748_ ) );
AOI21_X2 _12404_ ( .A(_04532_ ), .B1(_04740_ ), .B2(_04748_ ), .ZN(_04749_ ) );
INV_X1 _12405_ ( .A(_03253_ ), .ZN(_04750_ ) );
OR3_X1 _12406_ ( .A1(_04525_ ), .A2(_04750_ ), .A3(_04529_ ), .ZN(_04751_ ) );
OAI21_X1 _12407_ ( .A(_04751_ ), .B1(_03282_ ), .B2(_04524_ ), .ZN(_04752_ ) );
NOR2_X1 _12408_ ( .A1(_04515_ ), .A2(_04521_ ), .ZN(_04753_ ) );
AND2_X1 _12409_ ( .A1(_04752_ ), .A2(_04753_ ), .ZN(_04754_ ) );
INV_X1 _12410_ ( .A(_04754_ ), .ZN(_04755_ ) );
AOI21_X1 _12411_ ( .A(_04514_ ), .B1(_03307_ ), .B2(_03308_ ), .ZN(_04756_ ) );
NAND2_X1 _12412_ ( .A1(_04520_ ), .A2(_04756_ ), .ZN(_04757_ ) );
NAND2_X1 _12413_ ( .A1(_04516_ ), .A2(_04517_ ), .ZN(_04758_ ) );
INV_X1 _12414_ ( .A(_04758_ ), .ZN(_04759_ ) );
OAI211_X1 _12415_ ( .A(_04755_ ), .B(_04757_ ), .C1(_03337_ ), .C2(_04759_ ), .ZN(_04760_ ) );
AND2_X1 _12416_ ( .A1(_03602_ ), .A2(\ID_EX_typ [2] ), .ZN(_04761_ ) );
INV_X1 _12417_ ( .A(_04761_ ), .ZN(_04762_ ) );
OR3_X2 _12418_ ( .A1(_04749_ ), .A2(_04760_ ), .A3(_04762_ ), .ZN(_04763_ ) );
NOR2_X1 _12419_ ( .A1(_02419_ ), .A2(\ID_EX_typ [1] ), .ZN(_04764_ ) );
AND2_X1 _12420_ ( .A1(_04764_ ), .A2(\ID_EX_typ [2] ), .ZN(_04765_ ) );
NAND3_X1 _12421_ ( .A1(_04482_ ), .A2(_04505_ ), .A3(_04765_ ), .ZN(_04766_ ) );
AND2_X2 _12422_ ( .A1(_04763_ ), .A2(_04766_ ), .ZN(_04767_ ) );
INV_X1 _12423_ ( .A(_04506_ ), .ZN(_04768_ ) );
AOI21_X2 _12424_ ( .A(_04507_ ), .B1(_04767_ ), .B2(_04768_ ), .ZN(_04769_ ) );
NOR2_X1 _12425_ ( .A1(_04417_ ), .A2(fanout_net_5 ), .ZN(_04770_ ) );
INV_X1 _12426_ ( .A(\ID_EX_typ [2] ), .ZN(_04771_ ) );
AND2_X1 _12427_ ( .A1(_04770_ ), .A2(_04771_ ), .ZN(_04772_ ) );
OAI21_X1 _12428_ ( .A(_04772_ ), .B1(_04749_ ), .B2(_04760_ ), .ZN(_04773_ ) );
NAND2_X1 _12429_ ( .A1(_04773_ ), .A2(_04420_ ), .ZN(_04774_ ) );
OAI221_X2 _12430_ ( .A(_03604_ ), .B1(_04415_ ), .B2(_04420_ ), .C1(_04769_ ), .C2(_04774_ ), .ZN(_04775_ ) );
OR2_X2 _12431_ ( .A1(_04415_ ), .A2(_03604_ ), .ZN(_04776_ ) );
AND2_X4 _12432_ ( .A1(_04775_ ), .A2(_04776_ ), .ZN(_04777_ ) );
BUF_X16 _12433_ ( .A(_04777_ ), .Z(_04778_ ) );
MUX2_X1 _12434_ ( .A(_03600_ ), .B(_03601_ ), .S(_04778_ ), .Z(_04779_ ) );
OAI21_X1 _12435_ ( .A(_03581_ ), .B1(_04779_ ), .B2(fanout_net_6 ), .ZN(_04780_ ) );
MUX2_X2 _12436_ ( .A(_03519_ ), .B(_04780_ ), .S(_02411_ ), .Z(_04781_ ) );
INV_X1 _12437_ ( .A(_02415_ ), .ZN(_04782_ ) );
BUF_X4 _12438_ ( .A(_04782_ ), .Z(_04783_ ) );
AOI211_X1 _12439_ ( .A(_03406_ ), .B(_03518_ ), .C1(_04781_ ), .C2(_04783_ ), .ZN(_04784_ ) );
BUF_X2 _12440_ ( .A(_02419_ ), .Z(_04785_ ) );
OR3_X4 _12441_ ( .A1(_03347_ ), .A2(_04785_ ), .A3(_04782_ ), .ZN(_04786_ ) );
AND2_X1 _12442_ ( .A1(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .A2(_02403_ ), .ZN(\myidu.state_$_ANDNOT__A_Y ) );
INV_X1 _12443_ ( .A(\myidu.state_$_ANDNOT__A_Y ), .ZN(_04787_ ) );
BUF_X4 _12444_ ( .A(_04787_ ), .Z(_04788_ ) );
BUF_X2 _12445_ ( .A(_03401_ ), .Z(_04789_ ) );
NAND3_X1 _12446_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [30] ), .ZN(_04790_ ) );
AOI22_X1 _12447_ ( .A1(_04784_ ), .A2(_04786_ ), .B1(_04788_ ), .B2(_04790_ ), .ZN(_00123_ ) );
NAND2_X1 _12448_ ( .A1(_03508_ ), .A2(_03509_ ), .ZN(_04791_ ) );
XOR2_X1 _12449_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .Z(_04792_ ) );
XNOR2_X1 _12450_ ( .A(_04791_ ), .B(_04792_ ), .ZN(_04793_ ) );
NOR2_X1 _12451_ ( .A1(_04793_ ), .A2(_02420_ ), .ZN(_04794_ ) );
NOR2_X1 _12452_ ( .A1(_02396_ ), .A2(fanout_net_16 ), .ZN(_04795_ ) );
BUF_X4 _12453_ ( .A(_03560_ ), .Z(_04796_ ) );
NAND3_X1 _12454_ ( .A1(_03557_ ), .A2(\mepc [29] ), .A3(_04796_ ), .ZN(_04797_ ) );
BUF_X2 _12455_ ( .A(_03562_ ), .Z(_04798_ ) );
BUF_X4 _12456_ ( .A(_03565_ ), .Z(_04799_ ) );
BUF_X2 _12457_ ( .A(_03559_ ), .Z(_04800_ ) );
NAND4_X1 _12458_ ( .A1(_04798_ ), .A2(_04799_ ), .A3(\mycsreg.CSReg[3][29] ), .A4(_04800_ ), .ZN(_04801_ ) );
NAND4_X1 _12459_ ( .A1(_03569_ ), .A2(\mtvec [29] ), .A3(_04800_ ), .A4(_03574_ ), .ZN(_04802_ ) );
NAND4_X1 _12460_ ( .A1(_03552_ ), .A2(_04797_ ), .A3(_04801_ ), .A4(_04802_ ), .ZN(_04803_ ) );
AND4_X1 _12461_ ( .A1(\mycsreg.CSReg[0][29] ), .A2(_03573_ ), .A3(_04800_ ), .A4(_03574_ ), .ZN(_04804_ ) );
OAI22_X1 _12462_ ( .A1(_03540_ ), .A2(_03542_ ), .B1(_04803_ ), .B2(_04804_ ), .ZN(_04805_ ) );
NAND3_X1 _12463_ ( .A1(_03539_ ), .A2(\EX_LS_result_csreg_mem [29] ), .A3(_03577_ ), .ZN(_04806_ ) );
NAND2_X1 _12464_ ( .A1(_04805_ ), .A2(_04806_ ), .ZN(_04807_ ) );
AND2_X1 _12465_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_04808_ ) );
NAND3_X1 _12466_ ( .A1(_04808_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_04809_ ) );
NAND4_X1 _12467_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_04810_ ) );
NOR2_X1 _12468_ ( .A1(_04809_ ), .A2(_04810_ ), .ZN(_04811_ ) );
AND2_X1 _12469_ ( .A1(_03588_ ), .A2(_04811_ ), .ZN(_04812_ ) );
AND4_X1 _12470_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_04813_ ) );
AND2_X1 _12471_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_04814_ ) );
AND4_X1 _12472_ ( .A1(\ID_EX_pc [21] ), .A2(_04813_ ), .A3(\ID_EX_pc [20] ), .A4(_04814_ ), .ZN(_04815_ ) );
NAND2_X1 _12473_ ( .A1(_04812_ ), .A2(_04815_ ), .ZN(_04816_ ) );
INV_X1 _12474_ ( .A(\ID_EX_pc [27] ), .ZN(_04817_ ) );
INV_X1 _12475_ ( .A(\ID_EX_pc [26] ), .ZN(_04818_ ) );
NOR3_X1 _12476_ ( .A1(_04816_ ), .A2(_04817_ ), .A3(_04818_ ), .ZN(_04819_ ) );
NAND2_X1 _12477_ ( .A1(_04819_ ), .A2(\ID_EX_pc [28] ), .ZN(_04820_ ) );
XNOR2_X1 _12478_ ( .A(_04820_ ), .B(\ID_EX_pc [29] ), .ZN(_04821_ ) );
AOI21_X1 _12479_ ( .A(_04821_ ), .B1(_04775_ ), .B2(_04776_ ), .ZN(_04822_ ) );
AOI21_X2 _12480_ ( .A(_04822_ ), .B1(_04778_ ), .B2(_04793_ ), .ZN(_04823_ ) );
MUX2_X2 _12481_ ( .A(_04807_ ), .B(_04823_ ), .S(_03580_ ), .Z(_04824_ ) );
MUX2_X2 _12482_ ( .A(_04795_ ), .B(_04824_ ), .S(_02411_ ), .Z(_04825_ ) );
AOI211_X2 _12483_ ( .A(_03406_ ), .B(_04794_ ), .C1(_04825_ ), .C2(_04783_ ), .ZN(_04826_ ) );
NAND2_X1 _12484_ ( .A1(_02415_ ), .A2(fanout_net_5 ), .ZN(_04827_ ) );
BUF_X2 _12485_ ( .A(_04827_ ), .Z(_04828_ ) );
OR2_X1 _12486_ ( .A1(_03381_ ), .A2(_04828_ ), .ZN(_04829_ ) );
NAND3_X1 _12487_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [29] ), .ZN(_04830_ ) );
AOI22_X1 _12488_ ( .A1(_04826_ ), .A2(_04829_ ), .B1(_04788_ ), .B2(_04830_ ), .ZN(_00124_ ) );
BUF_X4 _12489_ ( .A(_04782_ ), .Z(_04831_ ) );
BUF_X4 _12490_ ( .A(_04831_ ), .Z(_04832_ ) );
BUF_X2 _12491_ ( .A(_03560_ ), .Z(_04833_ ) );
NAND3_X1 _12492_ ( .A1(_03557_ ), .A2(\mepc [20] ), .A3(_04833_ ), .ZN(_04834_ ) );
AND4_X1 _12493_ ( .A1(\ID_EX_csr [4] ), .A2(_03545_ ), .A3(_03546_ ), .A4(_03564_ ), .ZN(_04835_ ) );
NAND2_X1 _12494_ ( .A1(_04835_ ), .A2(_03551_ ), .ZN(_04836_ ) );
AND2_X1 _12495_ ( .A1(_03552_ ), .A2(_04836_ ), .ZN(_04837_ ) );
BUF_X4 _12496_ ( .A(_03562_ ), .Z(_04838_ ) );
NAND4_X1 _12497_ ( .A1(_04838_ ), .A2(_04799_ ), .A3(\mycsreg.CSReg[3][20] ), .A4(_04796_ ), .ZN(_04839_ ) );
NAND4_X1 _12498_ ( .A1(_03569_ ), .A2(\mtvec [20] ), .A3(_04796_ ), .A4(_03574_ ), .ZN(_04840_ ) );
AND4_X1 _12499_ ( .A1(_04834_ ), .A2(_04837_ ), .A3(_04839_ ), .A4(_04840_ ), .ZN(_04841_ ) );
BUF_X2 _12500_ ( .A(_03573_ ), .Z(_04842_ ) );
BUF_X2 _12501_ ( .A(_04842_ ), .Z(_04843_ ) );
BUF_X4 _12502_ ( .A(_03560_ ), .Z(_04844_ ) );
BUF_X2 _12503_ ( .A(_04844_ ), .Z(_04845_ ) );
BUF_X4 _12504_ ( .A(_03574_ ), .Z(_04846_ ) );
BUF_X4 _12505_ ( .A(_04846_ ), .Z(_04847_ ) );
NAND4_X1 _12506_ ( .A1(_04843_ ), .A2(_04845_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][20] ), .ZN(_04848_ ) );
BUF_X2 _12507_ ( .A(_03539_ ), .Z(_04849_ ) );
AOI22_X1 _12508_ ( .A1(_04841_ ), .A2(_04848_ ), .B1(_03577_ ), .B2(_04849_ ), .ZN(_04850_ ) );
AND3_X1 _12509_ ( .A1(_04849_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_03577_ ), .ZN(_04851_ ) );
NOR2_X1 _12510_ ( .A1(_04850_ ), .A2(_04851_ ), .ZN(_04852_ ) );
BUF_X4 _12511_ ( .A(_03580_ ), .Z(_04853_ ) );
NOR2_X1 _12512_ ( .A1(_04852_ ), .A2(_04853_ ), .ZN(_04854_ ) );
NAND3_X1 _12513_ ( .A1(_03588_ ), .A2(_04811_ ), .A3(_04814_ ), .ZN(_04855_ ) );
XNOR2_X1 _12514_ ( .A(_04855_ ), .B(\ID_EX_pc [20] ), .ZN(_04856_ ) );
XOR2_X1 _12515_ ( .A(_03481_ ), .B(_03486_ ), .Z(_04857_ ) );
BUF_X8 _12516_ ( .A(_04778_ ), .Z(_04858_ ) );
MUX2_X1 _12517_ ( .A(_04856_ ), .B(_04857_ ), .S(_04858_ ), .Z(_04859_ ) );
BUF_X4 _12518_ ( .A(_04853_ ), .Z(_04860_ ) );
AOI21_X1 _12519_ ( .A(_04854_ ), .B1(_04859_ ), .B2(_04860_ ), .ZN(_04861_ ) );
BUF_X4 _12520_ ( .A(_02421_ ), .Z(_04862_ ) );
NOR2_X1 _12521_ ( .A1(_04861_ ), .A2(_04862_ ), .ZN(_04863_ ) );
BUF_X2 _12522_ ( .A(_02421_ ), .Z(_04864_ ) );
AND3_X1 _12523_ ( .A1(_04864_ ), .A2(_03402_ ), .A3(\myexu.pc_jump [20] ), .ZN(_04865_ ) );
OAI21_X1 _12524_ ( .A(_04832_ ), .B1(_04863_ ), .B2(_04865_ ), .ZN(_04866_ ) );
NOR2_X1 _12525_ ( .A1(_03355_ ), .A2(_04828_ ), .ZN(_04867_ ) );
BUF_X4 _12526_ ( .A(_03405_ ), .Z(_04868_ ) );
CLKBUF_X2 _12527_ ( .A(_02419_ ), .Z(_04869_ ) );
CLKBUF_X2 _12528_ ( .A(_02415_ ), .Z(_04870_ ) );
AND3_X1 _12529_ ( .A1(_04857_ ), .A2(_04869_ ), .A3(_04870_ ), .ZN(_04871_ ) );
NOR3_X1 _12530_ ( .A1(_04867_ ), .A2(_04868_ ), .A3(_04871_ ), .ZN(_04872_ ) );
NAND3_X1 _12531_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [20] ), .ZN(_04873_ ) );
AOI22_X1 _12532_ ( .A1(_04866_ ), .A2(_04872_ ), .B1(_04788_ ), .B2(_04873_ ), .ZN(_00125_ ) );
BUF_X2 _12533_ ( .A(_02421_ ), .Z(_04874_ ) );
INV_X4 _12534_ ( .A(_04778_ ), .ZN(_04875_ ) );
NAND3_X1 _12535_ ( .A1(_03588_ ), .A2(\ID_EX_pc [18] ), .A3(_04811_ ), .ZN(_04876_ ) );
XNOR2_X1 _12536_ ( .A(_04876_ ), .B(\ID_EX_pc [19] ), .ZN(_04877_ ) );
AND2_X1 _12537_ ( .A1(_04875_ ), .A2(_04877_ ), .ZN(_04878_ ) );
BUF_X4 _12538_ ( .A(_04778_ ), .Z(_04879_ ) );
INV_X1 _12539_ ( .A(_03467_ ), .ZN(_04880_ ) );
OAI21_X1 _12540_ ( .A(_03471_ ), .B1(_03456_ ), .B2(_03464_ ), .ZN(_04881_ ) );
AOI21_X1 _12541_ ( .A(_04880_ ), .B1(_04881_ ), .B2(_03478_ ), .ZN(_04882_ ) );
NOR2_X1 _12542_ ( .A1(_04882_ ), .A2(_03473_ ), .ZN(_04883_ ) );
XNOR2_X1 _12543_ ( .A(_04883_ ), .B(_03466_ ), .ZN(_04884_ ) );
AOI211_X1 _12544_ ( .A(fanout_net_6 ), .B(_04878_ ), .C1(_04879_ ), .C2(_04884_ ), .ZN(_04885_ ) );
AND3_X1 _12545_ ( .A1(_03538_ ), .A2(_03577_ ), .A3(_03521_ ), .ZN(_04886_ ) );
NAND3_X1 _12546_ ( .A1(_04886_ ), .A2(_03524_ ), .A3(_03530_ ), .ZN(_04887_ ) );
CLKBUF_X2 _12547_ ( .A(_04887_ ), .Z(_04888_ ) );
NAND3_X1 _12548_ ( .A1(_03527_ ), .A2(_03535_ ), .A3(_03533_ ), .ZN(_04889_ ) );
CLKBUF_X2 _12549_ ( .A(_04889_ ), .Z(_04890_ ) );
OR3_X1 _12550_ ( .A1(_04888_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_04890_ ), .ZN(_04891_ ) );
AND3_X2 _12551_ ( .A1(_03551_ ), .A2(\ID_EX_csr [4] ), .A3(_03545_ ), .ZN(_04892_ ) );
AND2_X2 _12552_ ( .A1(_04892_ ), .A2(_03565_ ), .ZN(_04893_ ) );
INV_X1 _12553_ ( .A(_04893_ ), .ZN(_04894_ ) );
BUF_X4 _12554_ ( .A(_04798_ ), .Z(_04895_ ) );
BUF_X2 _12555_ ( .A(_04895_ ), .Z(_04896_ ) );
BUF_X2 _12556_ ( .A(_04799_ ), .Z(_04897_ ) );
BUF_X4 _12557_ ( .A(_04844_ ), .Z(_04898_ ) );
BUF_X4 _12558_ ( .A(_04898_ ), .Z(_04899_ ) );
NAND4_X1 _12559_ ( .A1(_04896_ ), .A2(_04897_ ), .A3(\mycsreg.CSReg[3][19] ), .A4(_04899_ ), .ZN(_04900_ ) );
NAND4_X1 _12560_ ( .A1(_03548_ ), .A2(_03567_ ), .A3(_03543_ ), .A4(_03555_ ), .ZN(_04901_ ) );
NAND3_X1 _12561_ ( .A1(_03550_ ), .A2(_03558_ ), .A3(\ID_EX_csr [2] ), .ZN(_04902_ ) );
NOR2_X1 _12562_ ( .A1(_04901_ ), .A2(_04902_ ), .ZN(_04903_ ) );
BUF_X2 _12563_ ( .A(_04903_ ), .Z(_04904_ ) );
NAND2_X1 _12564_ ( .A1(_04904_ ), .A2(\mtvec [19] ), .ZN(_04905_ ) );
NAND3_X1 _12565_ ( .A1(_04894_ ), .A2(_04900_ ), .A3(_04905_ ), .ZN(_04906_ ) );
BUF_X4 _12566_ ( .A(_03557_ ), .Z(_04907_ ) );
BUF_X2 _12567_ ( .A(_04796_ ), .Z(_04908_ ) );
NAND3_X1 _12568_ ( .A1(_04907_ ), .A2(\mepc [19] ), .A3(_04908_ ), .ZN(_04909_ ) );
NAND4_X1 _12569_ ( .A1(_04843_ ), .A2(_04908_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][19] ), .ZN(_04910_ ) );
AND2_X1 _12570_ ( .A1(_04909_ ), .A2(_04910_ ), .ZN(_04911_ ) );
BUF_X2 _12571_ ( .A(_04887_ ), .Z(_04912_ ) );
BUF_X2 _12572_ ( .A(_04889_ ), .Z(_04913_ ) );
BUF_X2 _12573_ ( .A(_04913_ ), .Z(_04914_ ) );
OAI21_X1 _12574_ ( .A(_04911_ ), .B1(_04912_ ), .B2(_04914_ ), .ZN(_04915_ ) );
OAI21_X1 _12575_ ( .A(_04891_ ), .B1(_04906_ ), .B2(_04915_ ), .ZN(_04916_ ) );
AOI211_X1 _12576_ ( .A(_04874_ ), .B(_04885_ ), .C1(fanout_net_6 ), .C2(_04916_ ), .ZN(_04917_ ) );
INV_X1 _12577_ ( .A(\myexu.pc_jump [19] ), .ZN(_04918_ ) );
BUF_X4 _12578_ ( .A(_02408_ ), .Z(_04919_ ) );
BUF_X4 _12579_ ( .A(_02409_ ), .Z(_04920_ ) );
AOI211_X1 _12580_ ( .A(fanout_net_16 ), .B(_04918_ ), .C1(_04919_ ), .C2(_04920_ ), .ZN(_04921_ ) );
OAI21_X1 _12581_ ( .A(_04832_ ), .B1(_04917_ ), .B2(_04921_ ), .ZN(_04922_ ) );
NOR2_X1 _12582_ ( .A1(_03363_ ), .A2(_04828_ ), .ZN(_04923_ ) );
AND3_X1 _12583_ ( .A1(_04884_ ), .A2(_04869_ ), .A3(_04870_ ), .ZN(_04924_ ) );
NOR3_X1 _12584_ ( .A1(_04923_ ), .A2(_04868_ ), .A3(_04924_ ), .ZN(_04925_ ) );
NAND3_X1 _12585_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [19] ), .ZN(_04926_ ) );
AOI22_X1 _12586_ ( .A1(_04922_ ), .A2(_04925_ ), .B1(_04788_ ), .B2(_04926_ ), .ZN(_00126_ ) );
XNOR2_X1 _12587_ ( .A(_04812_ ), .B(\ID_EX_pc [18] ), .ZN(_04927_ ) );
AOI21_X1 _12588_ ( .A(_04927_ ), .B1(_04775_ ), .B2(_04776_ ), .ZN(_04928_ ) );
AND3_X1 _12589_ ( .A1(_04881_ ), .A2(_04880_ ), .A3(_03478_ ), .ZN(_04929_ ) );
NOR2_X1 _12590_ ( .A1(_04929_ ), .A2(_04882_ ), .ZN(_04930_ ) );
AOI211_X1 _12591_ ( .A(fanout_net_6 ), .B(_04928_ ), .C1(_04879_ ), .C2(_04930_ ), .ZN(_04931_ ) );
AND4_X1 _12592_ ( .A1(\mycsreg.CSReg[3][18] ), .A2(_04798_ ), .A3(_04799_ ), .A4(_04800_ ), .ZN(_04932_ ) );
AND2_X1 _12593_ ( .A1(_03548_ ), .A2(_03546_ ), .ZN(_04933_ ) );
BUF_X2 _12594_ ( .A(_04933_ ), .Z(_04934_ ) );
AND4_X1 _12595_ ( .A1(\mepc [18] ), .A2(_04934_ ), .A3(_04798_ ), .A4(_04800_ ), .ZN(_04935_ ) );
NOR3_X1 _12596_ ( .A1(_04893_ ), .A2(_04932_ ), .A3(_04935_ ), .ZN(_04936_ ) );
INV_X1 _12597_ ( .A(\ID_EX_csr [4] ), .ZN(_04937_ ) );
AND3_X2 _12598_ ( .A1(_03559_ ), .A2(_04937_ ), .A3(_03545_ ), .ZN(_04938_ ) );
BUF_X4 _12599_ ( .A(_04938_ ), .Z(_04939_ ) );
BUF_X4 _12600_ ( .A(_03569_ ), .Z(_04940_ ) );
NAND3_X1 _12601_ ( .A1(_04939_ ), .A2(\mtvec [18] ), .A3(_04940_ ), .ZN(_04941_ ) );
BUF_X4 _12602_ ( .A(_03573_ ), .Z(_04942_ ) );
NAND3_X1 _12603_ ( .A1(_04939_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_04942_ ), .ZN(_04943_ ) );
AND2_X1 _12604_ ( .A1(_04941_ ), .A2(_04943_ ), .ZN(_04944_ ) );
INV_X1 _12605_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_04945_ ) );
OAI221_X1 _12606_ ( .A(_03536_ ), .B1(\EX_LS_dest_csreg_mem [3] ), .B2(_03567_ ), .C1(_04945_ ), .C2(\ID_EX_csr [9] ), .ZN(_04946_ ) );
INV_X1 _12607_ ( .A(\EX_LS_dest_csreg_mem [4] ), .ZN(_04947_ ) );
AOI22_X1 _12608_ ( .A1(_04947_ ), .A2(\ID_EX_csr [4] ), .B1(_03567_ ), .B2(\EX_LS_dest_csreg_mem [3] ), .ZN(_04948_ ) );
OAI221_X1 _12609_ ( .A(_04948_ ), .B1(\EX_LS_dest_csreg_mem [1] ), .B2(_03563_ ), .C1(_04947_ ), .C2(\ID_EX_csr [4] ), .ZN(_04949_ ) );
INV_X1 _12610_ ( .A(\EX_LS_dest_csreg_mem [5] ), .ZN(_04950_ ) );
AOI22_X1 _12611_ ( .A1(\EX_LS_dest_csreg_mem [1] ), .A2(_03563_ ), .B1(_04950_ ), .B2(\ID_EX_csr [5] ), .ZN(_04951_ ) );
OAI221_X1 _12612_ ( .A(_04951_ ), .B1(fanout_net_4 ), .B2(_03547_ ), .C1(_04950_ ), .C2(\ID_EX_csr [5] ), .ZN(_04952_ ) );
NOR3_X1 _12613_ ( .A1(_04946_ ), .A2(_04949_ ), .A3(_04952_ ), .ZN(_04953_ ) );
INV_X1 _12614_ ( .A(\EX_LS_dest_csreg_mem [7] ), .ZN(_04954_ ) );
AOI22_X1 _12615_ ( .A1(_04945_ ), .A2(\ID_EX_csr [9] ), .B1(_04954_ ), .B2(\ID_EX_csr [7] ), .ZN(_04955_ ) );
INV_X1 _12616_ ( .A(\ID_EX_csr [7] ), .ZN(_04956_ ) );
AOI22_X1 _12617_ ( .A1(fanout_net_4 ), .A2(_03547_ ), .B1(_04956_ ), .B2(\EX_LS_dest_csreg_mem [7] ), .ZN(_04957_ ) );
NAND4_X1 _12618_ ( .A1(_04955_ ), .A2(_03535_ ), .A3(_03531_ ), .A4(_04957_ ), .ZN(_04958_ ) );
NOR4_X1 _12619_ ( .A1(_04958_ ), .A2(_03541_ ), .A3(_03520_ ), .A4(_03525_ ), .ZN(_04959_ ) );
AOI22_X1 _12620_ ( .A1(_04936_ ), .A2(_04944_ ), .B1(_04953_ ), .B2(_04959_ ), .ZN(_04960_ ) );
AND3_X1 _12621_ ( .A1(_04953_ ), .A2(_04959_ ), .A3(\EX_LS_result_csreg_mem [18] ), .ZN(_04961_ ) );
NOR2_X1 _12622_ ( .A1(_04960_ ), .A2(_04961_ ), .ZN(_04962_ ) );
AOI211_X1 _12623_ ( .A(_04874_ ), .B(_04931_ ), .C1(fanout_net_6 ), .C2(_04962_ ), .ZN(_04963_ ) );
AND3_X1 _12624_ ( .A1(_04864_ ), .A2(_03402_ ), .A3(\myexu.pc_jump [18] ), .ZN(_04964_ ) );
OAI21_X1 _12625_ ( .A(_04832_ ), .B1(_04963_ ), .B2(_04964_ ), .ZN(_04965_ ) );
NOR2_X1 _12626_ ( .A1(_03364_ ), .A2(_04828_ ), .ZN(_04966_ ) );
NOR3_X1 _12627_ ( .A1(_04929_ ), .A2(_04882_ ), .A3(_02420_ ), .ZN(_04967_ ) );
NOR3_X1 _12628_ ( .A1(_04966_ ), .A2(_04868_ ), .A3(_04967_ ), .ZN(_04968_ ) );
NAND3_X1 _12629_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [18] ), .ZN(_04969_ ) );
AOI22_X1 _12630_ ( .A1(_04965_ ), .A2(_04968_ ), .B1(_04788_ ), .B2(_04969_ ), .ZN(_00127_ ) );
BUF_X4 _12631_ ( .A(_04875_ ), .Z(_04970_ ) );
INV_X1 _12632_ ( .A(_03588_ ), .ZN(_04971_ ) );
NOR2_X1 _12633_ ( .A1(_04971_ ), .A2(_04809_ ), .ZN(_04972_ ) );
NAND3_X1 _12634_ ( .A1(_04972_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_04973_ ) );
INV_X1 _12635_ ( .A(\ID_EX_pc [16] ), .ZN(_04974_ ) );
NOR2_X1 _12636_ ( .A1(_04973_ ), .A2(_04974_ ), .ZN(_04975_ ) );
XNOR2_X1 _12637_ ( .A(_04975_ ), .B(\ID_EX_pc [17] ), .ZN(_04976_ ) );
NAND2_X1 _12638_ ( .A1(_04970_ ), .A2(_04976_ ), .ZN(_04977_ ) );
BUF_X4 _12639_ ( .A(_03580_ ), .Z(_04978_ ) );
AND2_X1 _12640_ ( .A1(_03465_ ), .A2(_03469_ ), .ZN(_04979_ ) );
NOR2_X1 _12641_ ( .A1(_04979_ ), .A2(_03476_ ), .ZN(_04980_ ) );
XNOR2_X1 _12642_ ( .A(_04980_ ), .B(_03470_ ), .ZN(_04981_ ) );
OAI211_X1 _12643_ ( .A(_04977_ ), .B(_04978_ ), .C1(_04970_ ), .C2(_04981_ ), .ZN(_04982_ ) );
NAND3_X1 _12644_ ( .A1(_03557_ ), .A2(\mepc [17] ), .A3(_03560_ ), .ZN(_04983_ ) );
BUF_X4 _12645_ ( .A(_04838_ ), .Z(_04984_ ) );
BUF_X4 _12646_ ( .A(_04844_ ), .Z(_04985_ ) );
NAND4_X1 _12647_ ( .A1(_04984_ ), .A2(_04897_ ), .A3(\mycsreg.CSReg[3][17] ), .A4(_04985_ ), .ZN(_04986_ ) );
BUF_X4 _12648_ ( .A(_03569_ ), .Z(_04987_ ) );
BUF_X2 _12649_ ( .A(_03574_ ), .Z(_04988_ ) );
NAND4_X1 _12650_ ( .A1(_04987_ ), .A2(\mtvec [17] ), .A3(_04985_ ), .A4(_04988_ ), .ZN(_04989_ ) );
AND4_X1 _12651_ ( .A1(_04837_ ), .A2(_04983_ ), .A3(_04986_ ), .A4(_04989_ ), .ZN(_04990_ ) );
BUF_X2 _12652_ ( .A(_04843_ ), .Z(_04991_ ) );
BUF_X2 _12653_ ( .A(_04845_ ), .Z(_04992_ ) );
BUF_X4 _12654_ ( .A(_04847_ ), .Z(_04993_ ) );
NAND4_X1 _12655_ ( .A1(_04991_ ), .A2(_04992_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][17] ), .ZN(_04994_ ) );
BUF_X2 _12656_ ( .A(_03577_ ), .Z(_04995_ ) );
CLKBUF_X2 _12657_ ( .A(_03539_ ), .Z(_04996_ ) );
AOI22_X1 _12658_ ( .A1(_04990_ ), .A2(_04994_ ), .B1(_04995_ ), .B2(_04996_ ), .ZN(_04997_ ) );
BUF_X4 _12659_ ( .A(_03577_ ), .Z(_04998_ ) );
AND3_X1 _12660_ ( .A1(_04849_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_04998_ ), .ZN(_04999_ ) );
OAI21_X1 _12661_ ( .A(fanout_net_6 ), .B1(_04997_ ), .B2(_04999_ ), .ZN(_05000_ ) );
AOI21_X1 _12662_ ( .A(_04862_ ), .B1(_04982_ ), .B2(_05000_ ), .ZN(_05001_ ) );
INV_X1 _12663_ ( .A(\myexu.pc_jump [17] ), .ZN(_05002_ ) );
AOI211_X1 _12664_ ( .A(fanout_net_16 ), .B(_05002_ ), .C1(_04919_ ), .C2(_04920_ ), .ZN(_05003_ ) );
OAI21_X1 _12665_ ( .A(_04832_ ), .B1(_05001_ ), .B2(_05003_ ), .ZN(_05004_ ) );
NOR2_X1 _12666_ ( .A1(_03366_ ), .A2(_04828_ ), .ZN(_05005_ ) );
AND3_X1 _12667_ ( .A1(_04981_ ), .A2(_04869_ ), .A3(_04870_ ), .ZN(_05006_ ) );
NOR3_X1 _12668_ ( .A1(_05005_ ), .A2(_04868_ ), .A3(_05006_ ), .ZN(_05007_ ) );
NAND3_X1 _12669_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [17] ), .ZN(_05008_ ) );
AOI22_X1 _12670_ ( .A1(_05004_ ), .A2(_05007_ ), .B1(_04788_ ), .B2(_05008_ ), .ZN(_00128_ ) );
XNOR2_X1 _12671_ ( .A(_04973_ ), .B(_04974_ ), .ZN(_05009_ ) );
AOI21_X1 _12672_ ( .A(_05009_ ), .B1(_04775_ ), .B2(_04776_ ), .ZN(_05010_ ) );
XOR2_X1 _12673_ ( .A(_03465_ ), .B(_03469_ ), .Z(_05011_ ) );
AOI211_X1 _12674_ ( .A(fanout_net_6 ), .B(_05010_ ), .C1(_04879_ ), .C2(_05011_ ), .ZN(_05012_ ) );
AND2_X2 _12675_ ( .A1(_04892_ ), .A2(_04933_ ), .ZN(_05013_ ) );
NOR2_X1 _12676_ ( .A1(_05013_ ), .A2(_04893_ ), .ZN(_05014_ ) );
AND4_X2 _12677_ ( .A1(_03546_ ), .A2(_03564_ ), .A3(_03550_ ), .A4(_03558_ ), .ZN(_05015_ ) );
BUF_X2 _12678_ ( .A(_05015_ ), .Z(_05016_ ) );
NAND3_X1 _12679_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_04895_ ), .ZN(_05017_ ) );
NAND3_X1 _12680_ ( .A1(_04907_ ), .A2(\mepc [16] ), .A3(_04908_ ), .ZN(_05018_ ) );
NAND2_X1 _12681_ ( .A1(_04903_ ), .A2(\mtvec [16] ), .ZN(_05019_ ) );
NAND4_X1 _12682_ ( .A1(_05014_ ), .A2(_05017_ ), .A3(_05018_ ), .A4(_05019_ ), .ZN(_05020_ ) );
NAND4_X1 _12683_ ( .A1(_04843_ ), .A2(_04908_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][16] ), .ZN(_05021_ ) );
BUF_X2 _12684_ ( .A(_04887_ ), .Z(_05022_ ) );
OAI21_X1 _12685_ ( .A(_05021_ ), .B1(_05022_ ), .B2(_04913_ ), .ZN(_05023_ ) );
NOR2_X1 _12686_ ( .A1(_05020_ ), .A2(_05023_ ), .ZN(_05024_ ) );
NOR3_X1 _12687_ ( .A1(_04888_ ), .A2(\EX_LS_result_csreg_mem [16] ), .A3(_04890_ ), .ZN(_05025_ ) );
NOR2_X1 _12688_ ( .A1(_05024_ ), .A2(_05025_ ), .ZN(_05026_ ) );
INV_X1 _12689_ ( .A(_05026_ ), .ZN(_05027_ ) );
AOI211_X1 _12690_ ( .A(_04874_ ), .B(_05012_ ), .C1(fanout_net_6 ), .C2(_05027_ ), .ZN(_05028_ ) );
AND3_X1 _12691_ ( .A1(_04864_ ), .A2(_03402_ ), .A3(\myexu.pc_jump [16] ), .ZN(_05029_ ) );
OAI21_X1 _12692_ ( .A(_04832_ ), .B1(_05028_ ), .B2(_05029_ ), .ZN(_05030_ ) );
NOR3_X1 _12693_ ( .A1(_03367_ ), .A2(_03357_ ), .A3(_04827_ ), .ZN(_05031_ ) );
AND3_X1 _12694_ ( .A1(_05011_ ), .A2(_04869_ ), .A3(_04870_ ), .ZN(_05032_ ) );
NOR3_X1 _12695_ ( .A1(_05031_ ), .A2(_04868_ ), .A3(_05032_ ), .ZN(_05033_ ) );
NAND3_X1 _12696_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [16] ), .ZN(_05034_ ) );
AOI22_X1 _12697_ ( .A1(_05030_ ), .A2(_05033_ ), .B1(_04788_ ), .B2(_05034_ ), .ZN(_00129_ ) );
INV_X1 _12698_ ( .A(\ID_EX_pc [14] ), .ZN(_05035_ ) );
NOR3_X1 _12699_ ( .A1(_04971_ ), .A2(_05035_ ), .A3(_04809_ ), .ZN(_05036_ ) );
INV_X1 _12700_ ( .A(\ID_EX_pc [15] ), .ZN(_05037_ ) );
XNOR2_X1 _12701_ ( .A(_05036_ ), .B(_05037_ ), .ZN(_05038_ ) );
OR2_X1 _12702_ ( .A1(_04858_ ), .A2(_05038_ ), .ZN(_05039_ ) );
INV_X1 _12703_ ( .A(_03450_ ), .ZN(_05040_ ) );
OAI21_X1 _12704_ ( .A(_03455_ ), .B1(_03439_ ), .B2(_03447_ ), .ZN(_05041_ ) );
AOI21_X1 _12705_ ( .A(_05040_ ), .B1(_05041_ ), .B2(_03463_ ), .ZN(_05042_ ) );
NOR2_X1 _12706_ ( .A1(_05042_ ), .A2(_03457_ ), .ZN(_05043_ ) );
XNOR2_X1 _12707_ ( .A(_05043_ ), .B(_03449_ ), .ZN(_05044_ ) );
OAI211_X1 _12708_ ( .A(_05039_ ), .B(_04978_ ), .C1(_04970_ ), .C2(_05044_ ), .ZN(_05045_ ) );
BUF_X2 _12709_ ( .A(_04849_ ), .Z(_05046_ ) );
AND3_X1 _12710_ ( .A1(_05046_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_04995_ ), .ZN(_05047_ ) );
BUF_X4 _12711_ ( .A(_04998_ ), .Z(_05048_ ) );
BUF_X4 _12712_ ( .A(_03557_ ), .Z(_05049_ ) );
NAND3_X1 _12713_ ( .A1(_05049_ ), .A2(\mepc [15] ), .A3(_04985_ ), .ZN(_05050_ ) );
BUF_X4 _12714_ ( .A(_04799_ ), .Z(_05051_ ) );
BUF_X4 _12715_ ( .A(_04796_ ), .Z(_05052_ ) );
NAND4_X1 _12716_ ( .A1(_04895_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][15] ), .A4(_05052_ ), .ZN(_05053_ ) );
BUF_X4 _12717_ ( .A(_03569_ ), .Z(_05054_ ) );
BUF_X4 _12718_ ( .A(_04800_ ), .Z(_05055_ ) );
BUF_X4 _12719_ ( .A(_03574_ ), .Z(_05056_ ) );
NAND4_X1 _12720_ ( .A1(_05054_ ), .A2(\mtvec [15] ), .A3(_05055_ ), .A4(_05056_ ), .ZN(_05057_ ) );
AND4_X1 _12721_ ( .A1(_04836_ ), .A2(_05050_ ), .A3(_05053_ ), .A4(_05057_ ), .ZN(_05058_ ) );
BUF_X4 _12722_ ( .A(_04942_ ), .Z(_05059_ ) );
NAND4_X1 _12723_ ( .A1(_05059_ ), .A2(_04899_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][15] ), .ZN(_05060_ ) );
AOI22_X1 _12724_ ( .A1(_05046_ ), .A2(_05048_ ), .B1(_05058_ ), .B2(_05060_ ), .ZN(_05061_ ) );
OAI21_X1 _12725_ ( .A(fanout_net_6 ), .B1(_05047_ ), .B2(_05061_ ), .ZN(_05062_ ) );
AOI21_X1 _12726_ ( .A(_04862_ ), .B1(_05045_ ), .B2(_05062_ ), .ZN(_05063_ ) );
INV_X1 _12727_ ( .A(\myexu.pc_jump [15] ), .ZN(_05064_ ) );
AOI211_X1 _12728_ ( .A(fanout_net_16 ), .B(_05064_ ), .C1(_04919_ ), .C2(_04920_ ), .ZN(_05065_ ) );
OAI21_X1 _12729_ ( .A(_04832_ ), .B1(_05063_ ), .B2(_05065_ ), .ZN(_05066_ ) );
NOR2_X1 _12730_ ( .A1(_03374_ ), .A2(_04828_ ), .ZN(_05067_ ) );
AND3_X1 _12731_ ( .A1(_05044_ ), .A2(_04869_ ), .A3(_04870_ ), .ZN(_05068_ ) );
NOR3_X1 _12732_ ( .A1(_05067_ ), .A2(_04868_ ), .A3(_05068_ ), .ZN(_05069_ ) );
NAND3_X1 _12733_ ( .A1(_02041_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [15] ), .ZN(_05070_ ) );
AOI22_X1 _12734_ ( .A1(_05066_ ), .A2(_05069_ ), .B1(_04788_ ), .B2(_05070_ ), .ZN(_00130_ ) );
XNOR2_X1 _12735_ ( .A(_04972_ ), .B(\ID_EX_pc [14] ), .ZN(_05071_ ) );
NAND2_X1 _12736_ ( .A1(_04875_ ), .A2(_05071_ ), .ZN(_05072_ ) );
AND3_X1 _12737_ ( .A1(_05041_ ), .A2(_05040_ ), .A3(_03463_ ), .ZN(_05073_ ) );
NOR2_X1 _12738_ ( .A1(_05073_ ), .A2(_05042_ ), .ZN(_05074_ ) );
OAI211_X1 _12739_ ( .A(_05072_ ), .B(_04978_ ), .C1(_04970_ ), .C2(_05074_ ), .ZN(_05075_ ) );
BUF_X2 _12740_ ( .A(_03560_ ), .Z(_05076_ ) );
NAND3_X1 _12741_ ( .A1(_05049_ ), .A2(\mepc [14] ), .A3(_05076_ ), .ZN(_05077_ ) );
NAND4_X1 _12742_ ( .A1(_04984_ ), .A2(_04897_ ), .A3(\mycsreg.CSReg[3][14] ), .A4(_04985_ ), .ZN(_05078_ ) );
NAND4_X1 _12743_ ( .A1(_05054_ ), .A2(\mtvec [14] ), .A3(_04985_ ), .A4(_04988_ ), .ZN(_05079_ ) );
AND4_X1 _12744_ ( .A1(_04837_ ), .A2(_05077_ ), .A3(_05078_ ), .A4(_05079_ ), .ZN(_05080_ ) );
NAND4_X1 _12745_ ( .A1(_04991_ ), .A2(_04899_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][14] ), .ZN(_05081_ ) );
AOI22_X1 _12746_ ( .A1(_05080_ ), .A2(_05081_ ), .B1(_04995_ ), .B2(_04996_ ), .ZN(_05082_ ) );
AND3_X1 _12747_ ( .A1(_04849_ ), .A2(\EX_LS_result_csreg_mem [14] ), .A3(_04998_ ), .ZN(_05083_ ) );
OAI21_X1 _12748_ ( .A(fanout_net_6 ), .B1(_05082_ ), .B2(_05083_ ), .ZN(_05084_ ) );
AOI21_X1 _12749_ ( .A(_04862_ ), .B1(_05075_ ), .B2(_05084_ ), .ZN(_05085_ ) );
AND3_X1 _12750_ ( .A1(_04874_ ), .A2(_03402_ ), .A3(\myexu.pc_jump [14] ), .ZN(_05086_ ) );
OAI21_X1 _12751_ ( .A(_04832_ ), .B1(_05085_ ), .B2(_05086_ ), .ZN(_05087_ ) );
AND2_X1 _12752_ ( .A1(_02415_ ), .A2(fanout_net_5 ), .ZN(_05088_ ) );
NAND3_X1 _12753_ ( .A1(_03375_ ), .A2(_05088_ ), .A3(_03371_ ), .ZN(_05089_ ) );
OR3_X1 _12754_ ( .A1(_05073_ ), .A2(_05042_ ), .A3(_02420_ ), .ZN(_05090_ ) );
AND3_X1 _12755_ ( .A1(_05089_ ), .A2(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_05090_ ), .ZN(_05091_ ) );
BUF_X4 _12756_ ( .A(_01773_ ), .Z(_05092_ ) );
NAND3_X1 _12757_ ( .A1(_05092_ ), .A2(_04789_ ), .A3(\myexu.pc_jump [14] ), .ZN(_05093_ ) );
AOI22_X1 _12758_ ( .A1(_05087_ ), .A2(_05091_ ), .B1(_04788_ ), .B2(_05093_ ), .ZN(_00131_ ) );
NAND3_X1 _12759_ ( .A1(_03587_ ), .A2(\ID_EX_pc [9] ), .A3(_04808_ ), .ZN(_05094_ ) );
INV_X1 _12760_ ( .A(\ID_EX_pc [12] ), .ZN(_05095_ ) );
NOR2_X1 _12761_ ( .A1(_05094_ ), .A2(_05095_ ), .ZN(_05096_ ) );
XNOR2_X1 _12762_ ( .A(_05096_ ), .B(\ID_EX_pc [13] ), .ZN(_05097_ ) );
AOI21_X1 _12763_ ( .A(_05097_ ), .B1(_04775_ ), .B2(_04776_ ), .ZN(_05098_ ) );
OAI21_X1 _12764_ ( .A(_03452_ ), .B1(_03439_ ), .B2(_03447_ ), .ZN(_05099_ ) );
NAND2_X1 _12765_ ( .A1(_05099_ ), .A2(_03461_ ), .ZN(_05100_ ) );
XNOR2_X1 _12766_ ( .A(_05100_ ), .B(_03454_ ), .ZN(_05101_ ) );
AOI211_X1 _12767_ ( .A(fanout_net_6 ), .B(_05098_ ), .C1(_04879_ ), .C2(_05101_ ), .ZN(_05102_ ) );
AND2_X2 _12768_ ( .A1(_04953_ ), .A2(_04959_ ), .ZN(_05103_ ) );
NAND3_X1 _12769_ ( .A1(_04939_ ), .A2(\mtvec [13] ), .A3(_04940_ ), .ZN(_05104_ ) );
NAND3_X1 _12770_ ( .A1(_04938_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_04842_ ), .ZN(_05105_ ) );
NAND3_X1 _12771_ ( .A1(_05015_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_04838_ ), .ZN(_05106_ ) );
NAND4_X1 _12772_ ( .A1(_04934_ ), .A2(_04798_ ), .A3(\mepc [13] ), .A4(_04796_ ), .ZN(_05107_ ) );
NAND4_X1 _12773_ ( .A1(_05104_ ), .A2(_05105_ ), .A3(_05106_ ), .A4(_05107_ ), .ZN(_05108_ ) );
NOR3_X1 _12774_ ( .A1(_05103_ ), .A2(_05013_ ), .A3(_05108_ ), .ZN(_05109_ ) );
INV_X1 _12775_ ( .A(\EX_LS_result_csreg_mem [13] ), .ZN(_05110_ ) );
AND3_X1 _12776_ ( .A1(_04953_ ), .A2(_04959_ ), .A3(_05110_ ), .ZN(_05111_ ) );
NOR2_X1 _12777_ ( .A1(_05109_ ), .A2(_05111_ ), .ZN(_05112_ ) );
INV_X1 _12778_ ( .A(_05112_ ), .ZN(_05113_ ) );
AOI211_X1 _12779_ ( .A(_04874_ ), .B(_05102_ ), .C1(fanout_net_6 ), .C2(_05113_ ), .ZN(_05114_ ) );
AND3_X1 _12780_ ( .A1(_04874_ ), .A2(_03402_ ), .A3(\myexu.pc_jump [13] ), .ZN(_05115_ ) );
OAI21_X1 _12781_ ( .A(_04832_ ), .B1(_05114_ ), .B2(_05115_ ), .ZN(_05116_ ) );
NOR2_X1 _12782_ ( .A1(_03378_ ), .A2(_04828_ ), .ZN(_05117_ ) );
BUF_X4 _12783_ ( .A(_03406_ ), .Z(_05118_ ) );
AND3_X1 _12784_ ( .A1(_05101_ ), .A2(_04869_ ), .A3(_04870_ ), .ZN(_05119_ ) );
NOR3_X1 _12785_ ( .A1(_05117_ ), .A2(_05118_ ), .A3(_05119_ ), .ZN(_05120_ ) );
BUF_X4 _12786_ ( .A(_03402_ ), .Z(_05121_ ) );
NAND3_X1 _12787_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [13] ), .ZN(_05122_ ) );
AOI22_X1 _12788_ ( .A1(_05116_ ), .A2(_05120_ ), .B1(_04788_ ), .B2(_05122_ ), .ZN(_00132_ ) );
BUF_X4 _12789_ ( .A(_03542_ ), .Z(_05123_ ) );
NAND3_X1 _12790_ ( .A1(_05049_ ), .A2(\mepc [12] ), .A3(_05076_ ), .ZN(_05124_ ) );
NAND4_X1 _12791_ ( .A1(_04984_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][12] ), .A4(_05052_ ), .ZN(_05125_ ) );
BUF_X2 _12792_ ( .A(_04796_ ), .Z(_05126_ ) );
BUF_X4 _12793_ ( .A(_04846_ ), .Z(_05127_ ) );
NAND4_X1 _12794_ ( .A1(_05054_ ), .A2(\mtvec [12] ), .A3(_05126_ ), .A4(_05127_ ), .ZN(_05128_ ) );
NAND4_X1 _12795_ ( .A1(_04837_ ), .A2(_05124_ ), .A3(_05125_ ), .A4(_05128_ ), .ZN(_05129_ ) );
AND4_X1 _12796_ ( .A1(\mycsreg.CSReg[0][12] ), .A2(_04843_ ), .A3(_04908_ ), .A4(_04988_ ), .ZN(_05130_ ) );
OAI22_X1 _12797_ ( .A1(_03540_ ), .A2(_05123_ ), .B1(_05129_ ), .B2(_05130_ ), .ZN(_05131_ ) );
NAND3_X1 _12798_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [12] ), .A3(_04998_ ), .ZN(_05132_ ) );
AOI21_X1 _12799_ ( .A(_04853_ ), .B1(_05131_ ), .B2(_05132_ ), .ZN(_05133_ ) );
XNOR2_X1 _12800_ ( .A(_05094_ ), .B(\ID_EX_pc [12] ), .ZN(_05134_ ) );
XNOR2_X1 _12801_ ( .A(_03448_ ), .B(_03453_ ), .ZN(_05135_ ) );
MUX2_X1 _12802_ ( .A(_05134_ ), .B(_05135_ ), .S(_04858_ ), .Z(_05136_ ) );
AOI21_X1 _12803_ ( .A(_05133_ ), .B1(_05136_ ), .B2(_04860_ ), .ZN(_05137_ ) );
NOR2_X1 _12804_ ( .A1(_05137_ ), .A2(_04862_ ), .ZN(_05138_ ) );
INV_X1 _12805_ ( .A(\myexu.pc_jump [12] ), .ZN(_05139_ ) );
AOI211_X1 _12806_ ( .A(fanout_net_16 ), .B(_05139_ ), .C1(_04919_ ), .C2(_04920_ ), .ZN(_05140_ ) );
OAI21_X1 _12807_ ( .A(_04832_ ), .B1(_05138_ ), .B2(_05140_ ), .ZN(_05141_ ) );
NOR2_X1 _12808_ ( .A1(_03379_ ), .A2(_04828_ ), .ZN(_05142_ ) );
AND3_X1 _12809_ ( .A1(_05135_ ), .A2(_04869_ ), .A3(_04870_ ), .ZN(_05143_ ) );
NOR3_X1 _12810_ ( .A1(_05142_ ), .A2(_05118_ ), .A3(_05143_ ), .ZN(_05144_ ) );
BUF_X4 _12811_ ( .A(_04787_ ), .Z(_05145_ ) );
NAND3_X1 _12812_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [12] ), .ZN(_05146_ ) );
AOI22_X1 _12813_ ( .A1(_05141_ ), .A2(_05144_ ), .B1(_05145_ ), .B2(_05146_ ), .ZN(_00133_ ) );
BUF_X4 _12814_ ( .A(_04831_ ), .Z(_05147_ ) );
AND2_X1 _12815_ ( .A1(_03588_ ), .A2(\ID_EX_pc [10] ), .ZN(_05148_ ) );
INV_X1 _12816_ ( .A(\ID_EX_pc [11] ), .ZN(_05149_ ) );
XNOR2_X1 _12817_ ( .A(_05148_ ), .B(_05149_ ), .ZN(_05150_ ) );
OR2_X1 _12818_ ( .A1(_04858_ ), .A2(_05150_ ), .ZN(_05151_ ) );
INV_X1 _12819_ ( .A(_03434_ ), .ZN(_05152_ ) );
OAI21_X1 _12820_ ( .A(_03438_ ), .B1(_03430_ ), .B2(_03431_ ), .ZN(_05153_ ) );
AOI21_X1 _12821_ ( .A(_05152_ ), .B1(_05153_ ), .B2(_03445_ ), .ZN(_05154_ ) );
OR2_X1 _12822_ ( .A1(_05154_ ), .A2(_03440_ ), .ZN(_05155_ ) );
XNOR2_X1 _12823_ ( .A(_05155_ ), .B(_03433_ ), .ZN(_05156_ ) );
AOI21_X1 _12824_ ( .A(fanout_net_6 ), .B1(_04879_ ), .B2(_05156_ ), .ZN(_05157_ ) );
NAND3_X1 _12825_ ( .A1(_03557_ ), .A2(\mepc [11] ), .A3(_04833_ ), .ZN(_05158_ ) );
NAND4_X1 _12826_ ( .A1(_04838_ ), .A2(_04799_ ), .A3(\mycsreg.CSReg[3][11] ), .A4(_04796_ ), .ZN(_05159_ ) );
NAND4_X1 _12827_ ( .A1(_03569_ ), .A2(\mtvec [11] ), .A3(_04796_ ), .A4(_03574_ ), .ZN(_05160_ ) );
AND4_X1 _12828_ ( .A1(_04837_ ), .A2(_05158_ ), .A3(_05159_ ), .A4(_05160_ ), .ZN(_05161_ ) );
NAND4_X1 _12829_ ( .A1(_05059_ ), .A2(_04845_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][11] ), .ZN(_05162_ ) );
AOI22_X1 _12830_ ( .A1(_05161_ ), .A2(_05162_ ), .B1(_04998_ ), .B2(_04849_ ), .ZN(_05163_ ) );
AND3_X1 _12831_ ( .A1(_03539_ ), .A2(\EX_LS_result_csreg_mem [11] ), .A3(_03577_ ), .ZN(_05164_ ) );
OR2_X1 _12832_ ( .A1(_05163_ ), .A2(_05164_ ), .ZN(_05165_ ) );
AOI22_X1 _12833_ ( .A1(_05151_ ), .A2(_05157_ ), .B1(fanout_net_6 ), .B2(_05165_ ), .ZN(_05166_ ) );
NOR2_X1 _12834_ ( .A1(_05166_ ), .A2(_04862_ ), .ZN(_05167_ ) );
INV_X1 _12835_ ( .A(\myexu.pc_jump [11] ), .ZN(_05168_ ) );
AOI211_X1 _12836_ ( .A(fanout_net_16 ), .B(_05168_ ), .C1(_04919_ ), .C2(_04920_ ), .ZN(_05169_ ) );
OAI21_X1 _12837_ ( .A(_05147_ ), .B1(_05167_ ), .B2(_05169_ ), .ZN(_05170_ ) );
AND2_X1 _12838_ ( .A1(_02940_ ), .A2(_02965_ ), .ZN(_05171_ ) );
OAI21_X1 _12839_ ( .A(_05171_ ), .B1(_02911_ ), .B2(_02916_ ), .ZN(_05172_ ) );
AOI21_X1 _12840_ ( .A(_03013_ ), .B1(_05172_ ), .B2(_03019_ ), .ZN(_05173_ ) );
NOR2_X1 _12841_ ( .A1(_05173_ ), .A2(_03021_ ), .ZN(_05174_ ) );
XNOR2_X1 _12842_ ( .A(_05174_ ), .B(_02991_ ), .ZN(_05175_ ) );
NOR2_X1 _12843_ ( .A1(_05175_ ), .A2(_04828_ ), .ZN(_05176_ ) );
NOR2_X1 _12844_ ( .A1(_05156_ ), .A2(_02420_ ), .ZN(_05177_ ) );
NOR3_X1 _12845_ ( .A1(_05176_ ), .A2(_05118_ ), .A3(_05177_ ), .ZN(_05178_ ) );
NAND3_X1 _12846_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [11] ), .ZN(_05179_ ) );
AOI22_X1 _12847_ ( .A1(_05170_ ), .A2(_05178_ ), .B1(_05145_ ), .B2(_05179_ ), .ZN(_00134_ ) );
BUF_X2 _12848_ ( .A(_02415_ ), .Z(_05180_ ) );
INV_X1 _12849_ ( .A(\ID_EX_pc [28] ), .ZN(_05181_ ) );
XNOR2_X1 _12850_ ( .A(_04819_ ), .B(_05181_ ), .ZN(_05182_ ) );
XOR2_X1 _12851_ ( .A(_03506_ ), .B(_03507_ ), .Z(_05183_ ) );
MUX2_X1 _12852_ ( .A(_05182_ ), .B(_05183_ ), .S(_04778_ ), .Z(_05184_ ) );
AND2_X1 _12853_ ( .A1(_05184_ ), .A2(_03580_ ), .ZN(_05185_ ) );
NAND3_X1 _12854_ ( .A1(_05049_ ), .A2(\mepc [28] ), .A3(_05126_ ), .ZN(_05186_ ) );
NAND4_X1 _12855_ ( .A1(_04895_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][28] ), .A4(_05052_ ), .ZN(_05187_ ) );
NAND4_X1 _12856_ ( .A1(_05054_ ), .A2(\mtvec [28] ), .A3(_05052_ ), .A4(_05056_ ), .ZN(_05188_ ) );
NAND4_X1 _12857_ ( .A1(_03552_ ), .A2(_05186_ ), .A3(_05187_ ), .A4(_05188_ ), .ZN(_05189_ ) );
BUF_X2 _12858_ ( .A(_03573_ ), .Z(_05190_ ) );
AND4_X1 _12859_ ( .A1(\mycsreg.CSReg[0][28] ), .A2(_05190_ ), .A3(_05126_ ), .A4(_04988_ ), .ZN(_05191_ ) );
OAI22_X1 _12860_ ( .A1(_03540_ ), .A2(_03542_ ), .B1(_05189_ ), .B2(_05191_ ), .ZN(_05192_ ) );
NAND3_X1 _12861_ ( .A1(_04849_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_04998_ ), .ZN(_05193_ ) );
AOI21_X1 _12862_ ( .A(_03580_ ), .B1(_05192_ ), .B2(_05193_ ), .ZN(_05194_ ) );
OAI21_X1 _12863_ ( .A(_02411_ ), .B1(_05185_ ), .B2(_05194_ ), .ZN(_05195_ ) );
NAND3_X1 _12864_ ( .A1(_02421_ ), .A2(_03401_ ), .A3(\myexu.pc_jump [28] ), .ZN(_05196_ ) );
AOI21_X1 _12865_ ( .A(_05180_ ), .B1(_05195_ ), .B2(_05196_ ), .ZN(_05197_ ) );
AND3_X1 _12866_ ( .A1(_05183_ ), .A2(_04785_ ), .A3(_04870_ ), .ZN(_05198_ ) );
NOR3_X1 _12867_ ( .A1(_05197_ ), .A2(_04868_ ), .A3(_05198_ ), .ZN(_05199_ ) );
OR2_X1 _12868_ ( .A1(_03383_ ), .A2(_04828_ ), .ZN(_05200_ ) );
NAND3_X1 _12869_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [28] ), .ZN(_05201_ ) );
AOI22_X1 _12870_ ( .A1(_05199_ ), .A2(_05200_ ), .B1(_05145_ ), .B2(_05201_ ), .ZN(_00135_ ) );
INV_X1 _12871_ ( .A(\ID_EX_pc [10] ), .ZN(_05202_ ) );
XNOR2_X1 _12872_ ( .A(_03588_ ), .B(_05202_ ), .ZN(_05203_ ) );
AND2_X1 _12873_ ( .A1(_04875_ ), .A2(_05203_ ), .ZN(_05204_ ) );
AND3_X1 _12874_ ( .A1(_05153_ ), .A2(_05152_ ), .A3(_03445_ ), .ZN(_05205_ ) );
NOR2_X1 _12875_ ( .A1(_05205_ ), .A2(_05154_ ), .ZN(_05206_ ) );
AOI211_X1 _12876_ ( .A(fanout_net_6 ), .B(_05204_ ), .C1(_04879_ ), .C2(_05206_ ), .ZN(_05207_ ) );
NAND2_X1 _12877_ ( .A1(_04903_ ), .A2(\mtvec [10] ), .ZN(_05208_ ) );
OAI21_X1 _12878_ ( .A(_05208_ ), .B1(_05022_ ), .B2(_04913_ ), .ZN(_05209_ ) );
BUF_X2 _12879_ ( .A(_03562_ ), .Z(_05210_ ) );
AND4_X1 _12880_ ( .A1(\mycsreg.CSReg[3][10] ), .A2(_05210_ ), .A3(_04799_ ), .A4(_05076_ ), .ZN(_05211_ ) );
NAND3_X1 _12881_ ( .A1(_05049_ ), .A2(\mepc [10] ), .A3(_05055_ ), .ZN(_05212_ ) );
NAND4_X1 _12882_ ( .A1(_04942_ ), .A2(_05076_ ), .A3(_05056_ ), .A4(\mycsreg.CSReg[0][10] ), .ZN(_05213_ ) );
NAND2_X1 _12883_ ( .A1(_05212_ ), .A2(_05213_ ), .ZN(_05214_ ) );
NOR4_X1 _12884_ ( .A1(_05209_ ), .A2(_04893_ ), .A3(_05211_ ), .A4(_05214_ ), .ZN(_05215_ ) );
BUF_X2 _12885_ ( .A(_04889_ ), .Z(_05216_ ) );
NOR3_X1 _12886_ ( .A1(_04912_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_05216_ ), .ZN(_05217_ ) );
OR2_X1 _12887_ ( .A1(_05215_ ), .A2(_05217_ ), .ZN(_05218_ ) );
AOI211_X1 _12888_ ( .A(_04874_ ), .B(_05207_ ), .C1(fanout_net_6 ), .C2(_05218_ ), .ZN(_05219_ ) );
INV_X1 _12889_ ( .A(\myexu.pc_jump [10] ), .ZN(_05220_ ) );
AOI211_X1 _12890_ ( .A(fanout_net_16 ), .B(_05220_ ), .C1(_04919_ ), .C2(_04920_ ), .ZN(_05221_ ) );
OAI21_X1 _12891_ ( .A(_05147_ ), .B1(_05219_ ), .B2(_05221_ ), .ZN(_05222_ ) );
AND3_X1 _12892_ ( .A1(_05172_ ), .A2(_03013_ ), .A3(_03019_ ), .ZN(_05223_ ) );
NOR3_X1 _12893_ ( .A1(_05223_ ), .A2(_05173_ ), .A3(_04827_ ), .ZN(_05224_ ) );
NOR3_X1 _12894_ ( .A1(_05205_ ), .A2(_05154_ ), .A3(_02420_ ), .ZN(_05225_ ) );
NOR3_X1 _12895_ ( .A1(_05224_ ), .A2(_05118_ ), .A3(_05225_ ), .ZN(_05226_ ) );
NAND3_X1 _12896_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [10] ), .ZN(_05227_ ) );
AOI22_X1 _12897_ ( .A1(_05222_ ), .A2(_05226_ ), .B1(_05145_ ), .B2(_05227_ ), .ZN(_00136_ ) );
XNOR2_X1 _12898_ ( .A(_03587_ ), .B(\ID_EX_pc [9] ), .ZN(_05228_ ) );
NAND2_X1 _12899_ ( .A1(_04875_ ), .A2(_05228_ ), .ZN(_05229_ ) );
AND2_X1 _12900_ ( .A1(_03432_ ), .A2(_03436_ ), .ZN(_05230_ ) );
NOR2_X1 _12901_ ( .A1(_05230_ ), .A2(_03443_ ), .ZN(_05231_ ) );
XNOR2_X1 _12902_ ( .A(_05231_ ), .B(_03437_ ), .ZN(_05232_ ) );
OAI211_X1 _12903_ ( .A(_05229_ ), .B(_04978_ ), .C1(_04970_ ), .C2(_05232_ ), .ZN(_05233_ ) );
AND3_X1 _12904_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_04995_ ), .ZN(_05234_ ) );
NAND3_X1 _12905_ ( .A1(_04907_ ), .A2(\mepc [9] ), .A3(_04908_ ), .ZN(_05235_ ) );
NAND4_X1 _12906_ ( .A1(_04895_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][9] ), .A4(_05055_ ), .ZN(_05236_ ) );
NAND4_X1 _12907_ ( .A1(_04940_ ), .A2(\mtvec [9] ), .A3(_05055_ ), .A4(_05056_ ), .ZN(_05237_ ) );
AND4_X1 _12908_ ( .A1(_04836_ ), .A2(_05235_ ), .A3(_05236_ ), .A4(_05237_ ), .ZN(_05238_ ) );
NAND4_X1 _12909_ ( .A1(_05059_ ), .A2(_04899_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][9] ), .ZN(_05239_ ) );
AOI22_X1 _12910_ ( .A1(_05046_ ), .A2(_05048_ ), .B1(_05238_ ), .B2(_05239_ ), .ZN(_05240_ ) );
OAI21_X1 _12911_ ( .A(fanout_net_6 ), .B1(_05234_ ), .B2(_05240_ ), .ZN(_05241_ ) );
AOI21_X1 _12912_ ( .A(_04864_ ), .B1(_05233_ ), .B2(_05241_ ), .ZN(_05242_ ) );
INV_X1 _12913_ ( .A(\myexu.pc_jump [9] ), .ZN(_05243_ ) );
AOI211_X1 _12914_ ( .A(fanout_net_16 ), .B(_05243_ ), .C1(_04919_ ), .C2(_04920_ ), .ZN(_05244_ ) );
OAI21_X1 _12915_ ( .A(_05147_ ), .B1(_05242_ ), .B2(_05244_ ), .ZN(_05245_ ) );
INV_X1 _12916_ ( .A(_02940_ ), .ZN(_05246_ ) );
NOR2_X1 _12917_ ( .A1(_02917_ ), .A2(_05246_ ), .ZN(_05247_ ) );
OR2_X1 _12918_ ( .A1(_05247_ ), .A2(_03017_ ), .ZN(_05248_ ) );
XNOR2_X1 _12919_ ( .A(_05248_ ), .B(_02965_ ), .ZN(_05249_ ) );
BUF_X4 _12920_ ( .A(_04827_ ), .Z(_05250_ ) );
NOR2_X1 _12921_ ( .A1(_05249_ ), .A2(_05250_ ), .ZN(_05251_ ) );
AND3_X1 _12922_ ( .A1(_05232_ ), .A2(_04869_ ), .A3(_03517_ ), .ZN(_05252_ ) );
NOR3_X1 _12923_ ( .A1(_05251_ ), .A2(_05118_ ), .A3(_05252_ ), .ZN(_05253_ ) );
NAND3_X1 _12924_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [9] ), .ZN(_05254_ ) );
AOI22_X1 _12925_ ( .A1(_05245_ ), .A2(_05253_ ), .B1(_05145_ ), .B2(_05254_ ), .ZN(_00137_ ) );
NAND3_X1 _12926_ ( .A1(_04907_ ), .A2(\mepc [8] ), .A3(_04898_ ), .ZN(_05255_ ) );
NAND4_X1 _12927_ ( .A1(_04895_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][8] ), .A4(_05052_ ), .ZN(_05256_ ) );
NAND4_X1 _12928_ ( .A1(_05054_ ), .A2(\mtvec [8] ), .A3(_05126_ ), .A4(_05127_ ), .ZN(_05257_ ) );
NAND4_X1 _12929_ ( .A1(_04837_ ), .A2(_05255_ ), .A3(_05256_ ), .A4(_05257_ ), .ZN(_05258_ ) );
AND4_X1 _12930_ ( .A1(\mycsreg.CSReg[0][8] ), .A2(_04843_ ), .A3(_04908_ ), .A4(_04988_ ), .ZN(_05259_ ) );
OAI22_X1 _12931_ ( .A1(_03540_ ), .A2(_03542_ ), .B1(_05258_ ), .B2(_05259_ ), .ZN(_05260_ ) );
NAND3_X1 _12932_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [8] ), .A3(_04998_ ), .ZN(_05261_ ) );
AOI21_X1 _12933_ ( .A(_04853_ ), .B1(_05260_ ), .B2(_05261_ ), .ZN(_05262_ ) );
INV_X1 _12934_ ( .A(\ID_EX_pc [8] ), .ZN(_05263_ ) );
XNOR2_X1 _12935_ ( .A(_03586_ ), .B(_05263_ ), .ZN(_05264_ ) );
XOR2_X1 _12936_ ( .A(_03432_ ), .B(_03436_ ), .Z(_05265_ ) );
MUX2_X1 _12937_ ( .A(_05264_ ), .B(_05265_ ), .S(_04778_ ), .Z(_05266_ ) );
AOI21_X1 _12938_ ( .A(_05262_ ), .B1(_05266_ ), .B2(_04860_ ), .ZN(_05267_ ) );
NOR2_X1 _12939_ ( .A1(_05267_ ), .A2(_04862_ ), .ZN(_05268_ ) );
INV_X1 _12940_ ( .A(\myexu.pc_jump [8] ), .ZN(_05269_ ) );
BUF_X4 _12941_ ( .A(_02409_ ), .Z(_05270_ ) );
AOI211_X1 _12942_ ( .A(fanout_net_16 ), .B(_05269_ ), .C1(_04919_ ), .C2(_05270_ ), .ZN(_05271_ ) );
OAI21_X1 _12943_ ( .A(_05147_ ), .B1(_05268_ ), .B2(_05271_ ), .ZN(_05272_ ) );
XNOR2_X1 _12944_ ( .A(_02917_ ), .B(_05246_ ), .ZN(_05273_ ) );
NOR2_X1 _12945_ ( .A1(_05273_ ), .A2(_05250_ ), .ZN(_05274_ ) );
AND3_X1 _12946_ ( .A1(_05265_ ), .A2(_04869_ ), .A3(_03517_ ), .ZN(_05275_ ) );
NOR3_X1 _12947_ ( .A1(_05274_ ), .A2(_05118_ ), .A3(_05275_ ), .ZN(_05276_ ) );
NAND3_X1 _12948_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [8] ), .ZN(_05277_ ) );
AOI22_X1 _12949_ ( .A1(_05272_ ), .A2(_05276_ ), .B1(_05145_ ), .B2(_05277_ ), .ZN(_00138_ ) );
BUF_X4 _12950_ ( .A(_04938_ ), .Z(_05278_ ) );
NAND3_X1 _12951_ ( .A1(_05278_ ), .A2(\mtvec [7] ), .A3(_04940_ ), .ZN(_05279_ ) );
NAND3_X1 _12952_ ( .A1(_04939_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_04942_ ), .ZN(_05280_ ) );
NAND3_X1 _12953_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_05210_ ), .ZN(_05281_ ) );
NAND4_X1 _12954_ ( .A1(_04934_ ), .A2(_05210_ ), .A3(\mepc [7] ), .A4(_04833_ ), .ZN(_05282_ ) );
NAND4_X1 _12955_ ( .A1(_05279_ ), .A2(_05280_ ), .A3(_05281_ ), .A4(_05282_ ), .ZN(_05283_ ) );
OR4_X1 _12956_ ( .A1(_03542_ ), .A2(_04958_ ), .A3(_03520_ ), .A4(_03525_ ), .ZN(_05284_ ) );
OR3_X1 _12957_ ( .A1(_04946_ ), .A2(_04949_ ), .A3(_04952_ ), .ZN(_05285_ ) );
OAI21_X1 _12958_ ( .A(_05283_ ), .B1(_05284_ ), .B2(_05285_ ), .ZN(_05286_ ) );
NAND3_X1 _12959_ ( .A1(_04953_ ), .A2(_04959_ ), .A3(\EX_LS_result_csreg_mem [7] ), .ZN(_05287_ ) );
AND2_X1 _12960_ ( .A1(_05286_ ), .A2(_05287_ ), .ZN(_05288_ ) );
OR2_X1 _12961_ ( .A1(_05288_ ), .A2(_04853_ ), .ZN(_05289_ ) );
NAND2_X1 _12962_ ( .A1(_03428_ ), .A2(_03429_ ), .ZN(_05290_ ) );
NOR2_X1 _12963_ ( .A1(_03431_ ), .A2(_03409_ ), .ZN(_05291_ ) );
XOR2_X1 _12964_ ( .A(_05290_ ), .B(_05291_ ), .Z(_05292_ ) );
OAI21_X1 _12965_ ( .A(_04860_ ), .B1(_04970_ ), .B2(_05292_ ), .ZN(_05293_ ) );
INV_X1 _12966_ ( .A(\ID_EX_pc [7] ), .ZN(_05294_ ) );
XNOR2_X1 _12967_ ( .A(_03585_ ), .B(_05294_ ), .ZN(_05295_ ) );
AOI21_X1 _12968_ ( .A(_05295_ ), .B1(_04775_ ), .B2(_04776_ ), .ZN(_05296_ ) );
OAI211_X1 _12969_ ( .A(_02411_ ), .B(_05289_ ), .C1(_05293_ ), .C2(_05296_ ), .ZN(_05297_ ) );
AND2_X1 _12970_ ( .A1(_03401_ ), .A2(\myexu.pc_jump [7] ), .ZN(_05298_ ) );
OR2_X1 _12971_ ( .A1(_02411_ ), .A2(_05298_ ), .ZN(_05299_ ) );
NAND3_X1 _12972_ ( .A1(_05297_ ), .A2(_04832_ ), .A3(_05299_ ), .ZN(_05300_ ) );
OAI21_X1 _12973_ ( .A(_02909_ ), .B1(_02859_ ), .B2(_02864_ ), .ZN(_05301_ ) );
AND2_X1 _12974_ ( .A1(_05301_ ), .A2(_02915_ ), .ZN(_05302_ ) );
XNOR2_X1 _12975_ ( .A(_05302_ ), .B(_02887_ ), .ZN(_05303_ ) );
NOR2_X1 _12976_ ( .A1(_05303_ ), .A2(_05250_ ), .ZN(_05304_ ) );
CLKBUF_X2 _12977_ ( .A(_02419_ ), .Z(_05305_ ) );
AND3_X1 _12978_ ( .A1(_05292_ ), .A2(_05305_ ), .A3(_03517_ ), .ZN(_05306_ ) );
NOR3_X1 _12979_ ( .A1(_05304_ ), .A2(_05118_ ), .A3(_05306_ ), .ZN(_05307_ ) );
NAND3_X1 _12980_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [7] ), .ZN(_05308_ ) );
AOI22_X1 _12981_ ( .A1(_05300_ ), .A2(_05307_ ), .B1(_05145_ ), .B2(_05308_ ), .ZN(_00139_ ) );
NAND3_X1 _12982_ ( .A1(_04907_ ), .A2(\mepc [6] ), .A3(_04908_ ), .ZN(_05309_ ) );
NAND4_X1 _12983_ ( .A1(_04895_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][6] ), .A4(_05052_ ), .ZN(_05310_ ) );
NAND4_X1 _12984_ ( .A1(_05054_ ), .A2(\mtvec [6] ), .A3(_05126_ ), .A4(_05127_ ), .ZN(_05311_ ) );
NAND4_X1 _12985_ ( .A1(_03552_ ), .A2(_05309_ ), .A3(_05310_ ), .A4(_05311_ ), .ZN(_05312_ ) );
AND4_X1 _12986_ ( .A1(\mycsreg.CSReg[0][6] ), .A2(_04843_ ), .A3(_04908_ ), .A4(_04988_ ), .ZN(_05313_ ) );
OAI22_X1 _12987_ ( .A1(_03540_ ), .A2(_03542_ ), .B1(_05312_ ), .B2(_05313_ ), .ZN(_05314_ ) );
NAND3_X1 _12988_ ( .A1(_04849_ ), .A2(\EX_LS_result_csreg_mem [6] ), .A3(_04998_ ), .ZN(_05315_ ) );
AOI21_X1 _12989_ ( .A(_04853_ ), .B1(_05314_ ), .B2(_05315_ ), .ZN(_05316_ ) );
INV_X1 _12990_ ( .A(\ID_EX_pc [6] ), .ZN(_05317_ ) );
XNOR2_X1 _12991_ ( .A(_03584_ ), .B(_05317_ ), .ZN(_05318_ ) );
OR3_X1 _12992_ ( .A1(_03426_ ), .A2(_03410_ ), .A3(_03427_ ), .ZN(_05319_ ) );
AND2_X1 _12993_ ( .A1(_05319_ ), .A2(_03428_ ), .ZN(_05320_ ) );
MUX2_X1 _12994_ ( .A(_05318_ ), .B(_05320_ ), .S(_04778_ ), .Z(_05321_ ) );
AOI21_X1 _12995_ ( .A(_05316_ ), .B1(_05321_ ), .B2(_04860_ ), .ZN(_05322_ ) );
NOR2_X1 _12996_ ( .A1(_05322_ ), .A2(_04862_ ), .ZN(_05323_ ) );
AND2_X1 _12997_ ( .A1(_03401_ ), .A2(\myexu.pc_jump [6] ), .ZN(_05324_ ) );
AND2_X1 _12998_ ( .A1(_04864_ ), .A2(_05324_ ), .ZN(_05325_ ) );
OAI21_X1 _12999_ ( .A(_05147_ ), .B1(_05323_ ), .B2(_05325_ ), .ZN(_05326_ ) );
XNOR2_X1 _13000_ ( .A(_02865_ ), .B(_02910_ ), .ZN(_05327_ ) );
NOR2_X1 _13001_ ( .A1(_05327_ ), .A2(_05250_ ), .ZN(_05328_ ) );
AND4_X1 _13002_ ( .A1(_05305_ ), .A2(_05319_ ), .A3(_03517_ ), .A4(_03428_ ), .ZN(_05329_ ) );
NOR3_X1 _13003_ ( .A1(_05328_ ), .A2(_05118_ ), .A3(_05329_ ), .ZN(_05330_ ) );
NAND3_X1 _13004_ ( .A1(_05092_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [6] ), .ZN(_05331_ ) );
AOI22_X1 _13005_ ( .A1(_05326_ ), .A2(_05330_ ), .B1(_05145_ ), .B2(_05331_ ), .ZN(_00140_ ) );
XNOR2_X1 _13006_ ( .A(_03583_ ), .B(\ID_EX_pc [5] ), .ZN(_05332_ ) );
NAND2_X1 _13007_ ( .A1(_04875_ ), .A2(_05332_ ), .ZN(_05333_ ) );
NAND2_X1 _13008_ ( .A1(_03424_ ), .A2(_03425_ ), .ZN(_05334_ ) );
NOR2_X1 _13009_ ( .A1(_03427_ ), .A2(_03411_ ), .ZN(_05335_ ) );
XOR2_X1 _13010_ ( .A(_05334_ ), .B(_05335_ ), .Z(_05336_ ) );
OAI211_X1 _13011_ ( .A(_05333_ ), .B(_04978_ ), .C1(_04970_ ), .C2(_05336_ ), .ZN(_05337_ ) );
NAND3_X1 _13012_ ( .A1(_04907_ ), .A2(\mepc [5] ), .A3(_04898_ ), .ZN(_05338_ ) );
NAND4_X1 _13013_ ( .A1(_04984_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][5] ), .A4(_05126_ ), .ZN(_05339_ ) );
NAND4_X1 _13014_ ( .A1(_05054_ ), .A2(\mtvec [5] ), .A3(_05126_ ), .A4(_05127_ ), .ZN(_05340_ ) );
AND4_X1 _13015_ ( .A1(_03552_ ), .A2(_05338_ ), .A3(_05339_ ), .A4(_05340_ ), .ZN(_05341_ ) );
NAND4_X1 _13016_ ( .A1(_04991_ ), .A2(_04899_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][5] ), .ZN(_05342_ ) );
AOI22_X1 _13017_ ( .A1(_05046_ ), .A2(_05048_ ), .B1(_05341_ ), .B2(_05342_ ), .ZN(_05343_ ) );
AND3_X1 _13018_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [5] ), .A3(_04995_ ), .ZN(_05344_ ) );
OAI21_X1 _13019_ ( .A(fanout_net_6 ), .B1(_05343_ ), .B2(_05344_ ), .ZN(_05345_ ) );
AOI21_X1 _13020_ ( .A(_04864_ ), .B1(_05337_ ), .B2(_05345_ ), .ZN(_05346_ ) );
INV_X1 _13021_ ( .A(\myexu.pc_jump [5] ), .ZN(_05347_ ) );
AOI211_X1 _13022_ ( .A(fanout_net_16 ), .B(_05347_ ), .C1(_04919_ ), .C2(_05270_ ), .ZN(_05348_ ) );
OAI21_X1 _13023_ ( .A(_05147_ ), .B1(_05346_ ), .B2(_05348_ ), .ZN(_05349_ ) );
AND3_X1 _13024_ ( .A1(_05336_ ), .A2(_03516_ ), .A3(_02415_ ), .ZN(_05350_ ) );
NOR2_X1 _13025_ ( .A1(_02812_ ), .A2(_02858_ ), .ZN(_05351_ ) );
AND2_X1 _13026_ ( .A1(_02855_ ), .A2(\ID_EX_imm [4] ), .ZN(_05352_ ) );
NOR2_X1 _13027_ ( .A1(_05351_ ), .A2(_05352_ ), .ZN(_05353_ ) );
XOR2_X1 _13028_ ( .A(_05353_ ), .B(_02834_ ), .Z(_05354_ ) );
AOI211_X1 _13029_ ( .A(_03406_ ), .B(_05350_ ), .C1(_05354_ ), .C2(_05088_ ), .ZN(_05355_ ) );
BUF_X4 _13030_ ( .A(_01773_ ), .Z(_05356_ ) );
NAND3_X1 _13031_ ( .A1(_05356_ ), .A2(_05121_ ), .A3(\myexu.pc_jump [5] ), .ZN(_05357_ ) );
AOI22_X1 _13032_ ( .A1(_05349_ ), .A2(_05355_ ), .B1(_05145_ ), .B2(_05357_ ), .ZN(_00141_ ) );
NAND3_X1 _13033_ ( .A1(_05278_ ), .A2(\mtvec [4] ), .A3(_04940_ ), .ZN(_05358_ ) );
NAND3_X1 _13034_ ( .A1(_05278_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_04942_ ), .ZN(_05359_ ) );
NAND3_X1 _13035_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_05210_ ), .ZN(_05360_ ) );
NAND4_X1 _13036_ ( .A1(_04934_ ), .A2(_05210_ ), .A3(\mepc [4] ), .A4(_05076_ ), .ZN(_05361_ ) );
NAND4_X1 _13037_ ( .A1(_05358_ ), .A2(_05359_ ), .A3(_05360_ ), .A4(_05361_ ), .ZN(_05362_ ) );
NOR3_X1 _13038_ ( .A1(_05103_ ), .A2(_05013_ ), .A3(_05362_ ), .ZN(_05363_ ) );
BUF_X2 _13039_ ( .A(_04953_ ), .Z(_05364_ ) );
BUF_X2 _13040_ ( .A(_04959_ ), .Z(_05365_ ) );
INV_X1 _13041_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_05366_ ) );
AND3_X1 _13042_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_05366_ ), .ZN(_05367_ ) );
NOR2_X1 _13043_ ( .A1(_05363_ ), .A2(_05367_ ), .ZN(_05368_ ) );
OAI21_X1 _13044_ ( .A(_02411_ ), .B1(_05368_ ), .B2(_04978_ ), .ZN(_05369_ ) );
XNOR2_X1 _13045_ ( .A(_03582_ ), .B(\ID_EX_pc [4] ), .ZN(_05370_ ) );
XOR2_X1 _13046_ ( .A(_03422_ ), .B(_03423_ ), .Z(_05371_ ) );
INV_X1 _13047_ ( .A(_05371_ ), .ZN(_05372_ ) );
MUX2_X1 _13048_ ( .A(_05370_ ), .B(_05372_ ), .S(_04858_ ), .Z(_05373_ ) );
AOI21_X1 _13049_ ( .A(_05369_ ), .B1(_05373_ ), .B2(_04860_ ), .ZN(_05374_ ) );
AND3_X1 _13050_ ( .A1(_04874_ ), .A2(_03401_ ), .A3(\myexu.pc_jump [4] ), .ZN(_05375_ ) );
OAI21_X1 _13051_ ( .A(_05147_ ), .B1(_05374_ ), .B2(_05375_ ), .ZN(_05376_ ) );
XNOR2_X1 _13052_ ( .A(_02812_ ), .B(_02858_ ), .ZN(_05377_ ) );
NOR2_X1 _13053_ ( .A1(_05377_ ), .A2(_05250_ ), .ZN(_05378_ ) );
AND3_X1 _13054_ ( .A1(_05371_ ), .A2(_05305_ ), .A3(_03517_ ), .ZN(_05379_ ) );
NOR3_X1 _13055_ ( .A1(_05378_ ), .A2(_05118_ ), .A3(_05379_ ), .ZN(_05380_ ) );
BUF_X4 _13056_ ( .A(_03402_ ), .Z(_05381_ ) );
NAND3_X1 _13057_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [4] ), .ZN(_05382_ ) );
AOI22_X1 _13058_ ( .A1(_05376_ ), .A2(_05380_ ), .B1(_05145_ ), .B2(_05382_ ), .ZN(_00142_ ) );
XNOR2_X1 _13059_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .ZN(_05383_ ) );
AOI21_X1 _13060_ ( .A(_05383_ ), .B1(_04775_ ), .B2(_04776_ ), .ZN(_05384_ ) );
OAI21_X1 _13061_ ( .A(_03416_ ), .B1(_03419_ ), .B2(_03420_ ), .ZN(_05385_ ) );
INV_X1 _13062_ ( .A(_05385_ ), .ZN(_05386_ ) );
NOR2_X1 _13063_ ( .A1(_05386_ ), .A2(_03413_ ), .ZN(_05387_ ) );
XNOR2_X1 _13064_ ( .A(_05387_ ), .B(_03412_ ), .ZN(_05388_ ) );
AOI211_X1 _13065_ ( .A(fanout_net_6 ), .B(_05384_ ), .C1(_04879_ ), .C2(_05388_ ), .ZN(_05389_ ) );
NOR2_X1 _13066_ ( .A1(_04887_ ), .A2(_04889_ ), .ZN(_05390_ ) );
AND2_X1 _13067_ ( .A1(_05015_ ), .A2(_04798_ ), .ZN(_05391_ ) );
AOI22_X1 _13068_ ( .A1(_05391_ ), .A2(\mycsreg.CSReg[3][3] ), .B1(_04892_ ), .B2(_04934_ ), .ZN(_05392_ ) );
NAND3_X1 _13069_ ( .A1(_05049_ ), .A2(\mepc [3] ), .A3(_05076_ ), .ZN(_05393_ ) );
NAND4_X1 _13070_ ( .A1(_04842_ ), .A2(_04833_ ), .A3(_04846_ ), .A4(\mycsreg.CSReg[0][3] ), .ZN(_05394_ ) );
AND2_X1 _13071_ ( .A1(_05393_ ), .A2(_05394_ ), .ZN(_05395_ ) );
NAND2_X1 _13072_ ( .A1(_05392_ ), .A2(_05395_ ), .ZN(_05396_ ) );
AND2_X1 _13073_ ( .A1(_04904_ ), .A2(\mtvec [3] ), .ZN(_05397_ ) );
NOR3_X1 _13074_ ( .A1(_05390_ ), .A2(_05396_ ), .A3(_05397_ ), .ZN(_05398_ ) );
NOR3_X1 _13075_ ( .A1(_04912_ ), .A2(\EX_LS_result_csreg_mem [3] ), .A3(_05216_ ), .ZN(_05399_ ) );
NOR2_X1 _13076_ ( .A1(_05398_ ), .A2(_05399_ ), .ZN(_05400_ ) );
INV_X1 _13077_ ( .A(_05400_ ), .ZN(_05401_ ) );
AOI211_X1 _13078_ ( .A(_02421_ ), .B(_05389_ ), .C1(fanout_net_6 ), .C2(_05401_ ), .ZN(_05402_ ) );
INV_X1 _13079_ ( .A(\myexu.pc_jump [3] ), .ZN(_05403_ ) );
AOI211_X1 _13080_ ( .A(fanout_net_16 ), .B(_05403_ ), .C1(_04919_ ), .C2(_05270_ ), .ZN(_05404_ ) );
OAI21_X1 _13081_ ( .A(_05147_ ), .B1(_05402_ ), .B2(_05404_ ), .ZN(_05405_ ) );
OR3_X1 _13082_ ( .A1(_02807_ ), .A2(_02734_ ), .A3(_02808_ ), .ZN(_05406_ ) );
NAND3_X1 _13083_ ( .A1(_05406_ ), .A2(_05088_ ), .A3(_02809_ ), .ZN(_05407_ ) );
NAND3_X1 _13084_ ( .A1(_05388_ ), .A2(_04785_ ), .A3(_05180_ ), .ZN(_05408_ ) );
AND3_X1 _13085_ ( .A1(_05407_ ), .A2(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_05408_ ), .ZN(_05409_ ) );
BUF_X4 _13086_ ( .A(_04787_ ), .Z(_05410_ ) );
NAND3_X1 _13087_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [3] ), .ZN(_05411_ ) );
AOI22_X1 _13088_ ( .A1(_05405_ ), .A2(_05409_ ), .B1(_05410_ ), .B2(_05411_ ), .ZN(_00143_ ) );
OR2_X1 _13089_ ( .A1(_04858_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05412_ ) );
AOI211_X1 _13090_ ( .A(_03420_ ), .B(_03416_ ), .C1(_03418_ ), .C2(_03417_ ), .ZN(_05413_ ) );
NOR2_X1 _13091_ ( .A1(_05386_ ), .A2(_05413_ ), .ZN(_05414_ ) );
OAI211_X1 _13092_ ( .A(_05412_ ), .B(_04978_ ), .C1(_04970_ ), .C2(_05414_ ), .ZN(_05415_ ) );
AND3_X1 _13093_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_04995_ ), .ZN(_05416_ ) );
NAND3_X1 _13094_ ( .A1(_04907_ ), .A2(\mepc [2] ), .A3(_04908_ ), .ZN(_05417_ ) );
NAND4_X1 _13095_ ( .A1(_04895_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][2] ), .A4(_05055_ ), .ZN(_05418_ ) );
NAND4_X1 _13096_ ( .A1(_04940_ ), .A2(\mtvec [2] ), .A3(_05055_ ), .A4(_05056_ ), .ZN(_05419_ ) );
AND4_X1 _13097_ ( .A1(_04836_ ), .A2(_05417_ ), .A3(_05418_ ), .A4(_05419_ ), .ZN(_05420_ ) );
NAND4_X1 _13098_ ( .A1(_05059_ ), .A2(_04899_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][2] ), .ZN(_05421_ ) );
AOI22_X1 _13099_ ( .A1(_05046_ ), .A2(_05048_ ), .B1(_05420_ ), .B2(_05421_ ), .ZN(_05422_ ) );
OAI21_X1 _13100_ ( .A(fanout_net_6 ), .B1(_05416_ ), .B2(_05422_ ), .ZN(_05423_ ) );
AOI21_X1 _13101_ ( .A(_04864_ ), .B1(_05415_ ), .B2(_05423_ ), .ZN(_05424_ ) );
INV_X1 _13102_ ( .A(\myexu.pc_jump [2] ), .ZN(_05425_ ) );
AOI211_X1 _13103_ ( .A(fanout_net_16 ), .B(_05425_ ), .C1(_02408_ ), .C2(_05270_ ), .ZN(_05426_ ) );
OAI21_X1 _13104_ ( .A(_05147_ ), .B1(_05424_ ), .B2(_05426_ ), .ZN(_05427_ ) );
AND3_X1 _13105_ ( .A1(_02804_ ), .A2(_02806_ ), .A3(_02758_ ), .ZN(_05428_ ) );
NOR3_X1 _13106_ ( .A1(_05428_ ), .A2(_02807_ ), .A3(_04827_ ), .ZN(_05429_ ) );
NOR3_X1 _13107_ ( .A1(_05386_ ), .A2(_02420_ ), .A3(_05413_ ), .ZN(_05430_ ) );
NOR3_X1 _13108_ ( .A1(_05429_ ), .A2(_05118_ ), .A3(_05430_ ), .ZN(_05431_ ) );
NAND3_X1 _13109_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [2] ), .ZN(_05432_ ) );
AOI22_X1 _13110_ ( .A1(_05427_ ), .A2(_05431_ ), .B1(_05410_ ), .B2(_05432_ ), .ZN(_00144_ ) );
OR2_X1 _13111_ ( .A1(_04858_ ), .A2(\ID_EX_pc [1] ), .ZN(_05433_ ) );
XOR2_X1 _13112_ ( .A(_03417_ ), .B(_03418_ ), .Z(_05434_ ) );
OAI211_X1 _13113_ ( .A(_05433_ ), .B(_04978_ ), .C1(_04970_ ), .C2(_05434_ ), .ZN(_05435_ ) );
AND3_X1 _13114_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_04995_ ), .ZN(_05436_ ) );
NAND3_X1 _13115_ ( .A1(_04907_ ), .A2(\mepc [1] ), .A3(_04898_ ), .ZN(_05437_ ) );
NAND4_X1 _13116_ ( .A1(_04984_ ), .A2(_04897_ ), .A3(\mycsreg.CSReg[3][1] ), .A4(_04898_ ), .ZN(_05438_ ) );
NAND4_X1 _13117_ ( .A1(_05054_ ), .A2(\mtvec [1] ), .A3(_05126_ ), .A4(_04988_ ), .ZN(_05439_ ) );
NAND4_X1 _13118_ ( .A1(_05190_ ), .A2(_04985_ ), .A3(_05127_ ), .A4(\mycsreg.CSReg[0][1] ), .ZN(_05440_ ) );
AND4_X1 _13119_ ( .A1(_05437_ ), .A2(_05438_ ), .A3(_05439_ ), .A4(_05440_ ), .ZN(_05441_ ) );
AOI21_X1 _13120_ ( .A(_05441_ ), .B1(_05046_ ), .B2(_05048_ ), .ZN(_05442_ ) );
OAI21_X1 _13121_ ( .A(fanout_net_6 ), .B1(_05436_ ), .B2(_05442_ ), .ZN(_05443_ ) );
AOI21_X1 _13122_ ( .A(_04864_ ), .B1(_05435_ ), .B2(_05443_ ), .ZN(_05444_ ) );
INV_X1 _13123_ ( .A(\myexu.pc_jump [1] ), .ZN(_05445_ ) );
AOI211_X1 _13124_ ( .A(fanout_net_16 ), .B(_05445_ ), .C1(_02408_ ), .C2(_05270_ ), .ZN(_05446_ ) );
OAI21_X1 _13125_ ( .A(_05147_ ), .B1(_05444_ ), .B2(_05446_ ), .ZN(_05447_ ) );
XNOR2_X1 _13126_ ( .A(_02781_ ), .B(_02803_ ), .ZN(_05448_ ) );
NOR2_X1 _13127_ ( .A1(_05448_ ), .A2(_05250_ ), .ZN(_05449_ ) );
AND3_X1 _13128_ ( .A1(_05434_ ), .A2(_05305_ ), .A3(_03517_ ), .ZN(_05450_ ) );
NOR3_X1 _13129_ ( .A1(_05449_ ), .A2(_03406_ ), .A3(_05450_ ), .ZN(_05451_ ) );
NAND3_X1 _13130_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [1] ), .ZN(_05452_ ) );
AOI22_X1 _13131_ ( .A1(_05447_ ), .A2(_05451_ ), .B1(_05410_ ), .B2(_05452_ ), .ZN(_00145_ ) );
BUF_X4 _13132_ ( .A(_04831_ ), .Z(_05453_ ) );
NAND4_X1 _13133_ ( .A1(_04843_ ), .A2(_04845_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][27] ), .ZN(_05454_ ) );
OAI21_X1 _13134_ ( .A(_05454_ ), .B1(_04888_ ), .B2(_04890_ ), .ZN(_05455_ ) );
BUF_X2 _13135_ ( .A(_04934_ ), .Z(_05456_ ) );
AOI22_X1 _13136_ ( .A1(_05391_ ), .A2(\mycsreg.CSReg[3][27] ), .B1(_04892_ ), .B2(_05456_ ), .ZN(_05457_ ) );
NAND3_X1 _13137_ ( .A1(_04907_ ), .A2(\mepc [27] ), .A3(_04845_ ), .ZN(_05458_ ) );
NAND2_X1 _13138_ ( .A1(_04904_ ), .A2(\mtvec [27] ), .ZN(_05459_ ) );
NAND3_X1 _13139_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(_05459_ ), .ZN(_05460_ ) );
NOR2_X1 _13140_ ( .A1(_05455_ ), .A2(_05460_ ), .ZN(_05461_ ) );
NOR3_X1 _13141_ ( .A1(_04912_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_05216_ ), .ZN(_05462_ ) );
NOR2_X1 _13142_ ( .A1(_05461_ ), .A2(_05462_ ), .ZN(_05463_ ) );
OAI21_X1 _13143_ ( .A(_02411_ ), .B1(_05463_ ), .B2(_04978_ ), .ZN(_05464_ ) );
NAND3_X1 _13144_ ( .A1(_04812_ ), .A2(\ID_EX_pc [26] ), .A3(_04815_ ), .ZN(_05465_ ) );
XNOR2_X1 _13145_ ( .A(_05465_ ), .B(_04817_ ), .ZN(_05466_ ) );
NAND2_X1 _13146_ ( .A1(_03500_ ), .A2(_03502_ ), .ZN(_05467_ ) );
NAND2_X1 _13147_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_05468_ ) );
NAND2_X1 _13148_ ( .A1(_05467_ ), .A2(_05468_ ), .ZN(_05469_ ) );
XNOR2_X1 _13149_ ( .A(_05469_ ), .B(_03501_ ), .ZN(_05470_ ) );
MUX2_X1 _13150_ ( .A(_05466_ ), .B(_05470_ ), .S(_04858_ ), .Z(_05471_ ) );
AOI21_X1 _13151_ ( .A(_05464_ ), .B1(_05471_ ), .B2(_04860_ ), .ZN(_05472_ ) );
INV_X1 _13152_ ( .A(\myexu.pc_jump [27] ), .ZN(_05473_ ) );
AOI211_X1 _13153_ ( .A(fanout_net_16 ), .B(_05473_ ), .C1(_02408_ ), .C2(_05270_ ), .ZN(_05474_ ) );
OAI21_X1 _13154_ ( .A(_05453_ ), .B1(_05472_ ), .B2(_05474_ ), .ZN(_05475_ ) );
NOR3_X1 _13155_ ( .A1(_03386_ ), .A2(_04785_ ), .A3(_04831_ ), .ZN(_05476_ ) );
NOR2_X1 _13156_ ( .A1(_05470_ ), .A2(_02420_ ), .ZN(_05477_ ) );
NOR3_X1 _13157_ ( .A1(_05476_ ), .A2(_03406_ ), .A3(_05477_ ), .ZN(_05478_ ) );
NAND3_X1 _13158_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [27] ), .ZN(_05479_ ) );
AOI22_X1 _13159_ ( .A1(_05475_ ), .A2(_05478_ ), .B1(_05410_ ), .B2(_05479_ ), .ZN(_00146_ ) );
NAND3_X1 _13160_ ( .A1(_03557_ ), .A2(\mepc [0] ), .A3(_04833_ ), .ZN(_05480_ ) );
NAND4_X1 _13161_ ( .A1(_04838_ ), .A2(_04799_ ), .A3(\mycsreg.CSReg[3][0] ), .A4(_04844_ ), .ZN(_05481_ ) );
NAND4_X1 _13162_ ( .A1(_03569_ ), .A2(\mtvec [0] ), .A3(_04844_ ), .A4(_04846_ ), .ZN(_05482_ ) );
NAND4_X1 _13163_ ( .A1(_04836_ ), .A2(_05480_ ), .A3(_05481_ ), .A4(_05482_ ), .ZN(_05483_ ) );
AND4_X1 _13164_ ( .A1(\mycsreg.CSReg[0][0] ), .A2(_04842_ ), .A3(_04833_ ), .A4(_04846_ ), .ZN(_05484_ ) );
OAI22_X1 _13165_ ( .A1(_03540_ ), .A2(_03542_ ), .B1(_05483_ ), .B2(_05484_ ), .ZN(_05485_ ) );
NAND3_X1 _13166_ ( .A1(_04849_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_03577_ ), .ZN(_05486_ ) );
AND2_X1 _13167_ ( .A1(_05485_ ), .A2(_05486_ ), .ZN(_05487_ ) );
INV_X1 _13168_ ( .A(\ID_EX_pc [0] ), .ZN(_05488_ ) );
XNOR2_X1 _13169_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .ZN(_05489_ ) );
MUX2_X1 _13170_ ( .A(_05488_ ), .B(_05489_ ), .S(_04778_ ), .Z(_05490_ ) );
MUX2_X1 _13171_ ( .A(_05487_ ), .B(_05490_ ), .S(_04853_ ), .Z(_05491_ ) );
NOR2_X1 _13172_ ( .A1(_05491_ ), .A2(_04862_ ), .ZN(_05492_ ) );
AND3_X1 _13173_ ( .A1(_04874_ ), .A2(_03401_ ), .A3(\myexu.pc_jump [0] ), .ZN(_05493_ ) );
OAI21_X1 _13174_ ( .A(_05453_ ), .B1(_05492_ ), .B2(_05493_ ), .ZN(_05494_ ) );
INV_X1 _13175_ ( .A(_02413_ ), .ZN(_05495_ ) );
NOR3_X1 _13176_ ( .A1(_05489_ ), .A2(_05495_ ), .A3(_02406_ ), .ZN(_05496_ ) );
AOI21_X1 _13177_ ( .A(_04868_ ), .B1(_05496_ ), .B2(\myexu.pc_jump_$_SDFF_PP0__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_05497_ ) );
NAND3_X1 _13178_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [0] ), .ZN(_05498_ ) );
AOI22_X1 _13179_ ( .A1(_05494_ ), .A2(_05497_ ), .B1(_05410_ ), .B2(_05498_ ), .ZN(_00147_ ) );
XOR2_X1 _13180_ ( .A(_03500_ ), .B(_03502_ ), .Z(_05499_ ) );
INV_X1 _13181_ ( .A(_05499_ ), .ZN(_05500_ ) );
AOI21_X1 _13182_ ( .A(fanout_net_6 ), .B1(_04879_ ), .B2(_05500_ ), .ZN(_05501_ ) );
XNOR2_X1 _13183_ ( .A(_04816_ ), .B(\ID_EX_pc [26] ), .ZN(_05502_ ) );
OAI21_X1 _13184_ ( .A(_05501_ ), .B1(_04879_ ), .B2(_05502_ ), .ZN(_05503_ ) );
AND3_X1 _13185_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_04995_ ), .ZN(_05504_ ) );
NAND3_X1 _13186_ ( .A1(_04907_ ), .A2(\mepc [26] ), .A3(_04898_ ), .ZN(_05505_ ) );
NAND4_X1 _13187_ ( .A1(_04984_ ), .A2(_04897_ ), .A3(\mycsreg.CSReg[3][26] ), .A4(_04985_ ), .ZN(_05506_ ) );
NAND4_X1 _13188_ ( .A1(_05054_ ), .A2(\mtvec [26] ), .A3(_05126_ ), .A4(_04988_ ), .ZN(_05507_ ) );
NAND4_X1 _13189_ ( .A1(_05190_ ), .A2(_04985_ ), .A3(_05127_ ), .A4(\mycsreg.CSReg[0][26] ), .ZN(_05508_ ) );
AND4_X1 _13190_ ( .A1(_05505_ ), .A2(_05506_ ), .A3(_05507_ ), .A4(_05508_ ), .ZN(_05509_ ) );
AOI21_X1 _13191_ ( .A(_05509_ ), .B1(_05046_ ), .B2(_05048_ ), .ZN(_05510_ ) );
OAI21_X1 _13192_ ( .A(fanout_net_6 ), .B1(_05504_ ), .B2(_05510_ ), .ZN(_05511_ ) );
AOI21_X1 _13193_ ( .A(_04864_ ), .B1(_05503_ ), .B2(_05511_ ), .ZN(_05512_ ) );
AOI211_X1 _13194_ ( .A(fanout_net_16 ), .B(_02391_ ), .C1(_02408_ ), .C2(_05270_ ), .ZN(_05513_ ) );
OAI21_X1 _13195_ ( .A(_05453_ ), .B1(_05512_ ), .B2(_05513_ ), .ZN(_05514_ ) );
NOR2_X1 _13196_ ( .A1(_03388_ ), .A2(_05250_ ), .ZN(_05515_ ) );
AND3_X1 _13197_ ( .A1(_05499_ ), .A2(_05305_ ), .A3(_03517_ ), .ZN(_05516_ ) );
NOR3_X1 _13198_ ( .A1(_05515_ ), .A2(_03406_ ), .A3(_05516_ ), .ZN(_05517_ ) );
NAND3_X1 _13199_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [26] ), .ZN(_05518_ ) );
AOI22_X1 _13200_ ( .A1(_05514_ ), .A2(_05517_ ), .B1(_05410_ ), .B2(_05518_ ), .ZN(_00148_ ) );
AND3_X1 _13201_ ( .A1(_04814_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05519_ ) );
AND2_X1 _13202_ ( .A1(_04812_ ), .A2(_05519_ ), .ZN(_05520_ ) );
NAND3_X1 _13203_ ( .A1(_05520_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05521_ ) );
INV_X1 _13204_ ( .A(\ID_EX_pc [24] ), .ZN(_05522_ ) );
NOR2_X1 _13205_ ( .A1(_05521_ ), .A2(_05522_ ), .ZN(_05523_ ) );
INV_X1 _13206_ ( .A(\ID_EX_pc [25] ), .ZN(_05524_ ) );
XNOR2_X1 _13207_ ( .A(_05523_ ), .B(_05524_ ), .ZN(_05525_ ) );
NAND2_X1 _13208_ ( .A1(_04875_ ), .A2(_05525_ ), .ZN(_05526_ ) );
OR2_X1 _13209_ ( .A1(_03488_ ), .A2(_03495_ ), .ZN(_05527_ ) );
AND2_X1 _13210_ ( .A1(_05527_ ), .A2(_03408_ ), .ZN(_05528_ ) );
OR2_X1 _13211_ ( .A1(_05528_ ), .A2(_03497_ ), .ZN(_05529_ ) );
XNOR2_X1 _13212_ ( .A(_05529_ ), .B(_03407_ ), .ZN(_05530_ ) );
OAI211_X1 _13213_ ( .A(_05526_ ), .B(_04853_ ), .C1(_04970_ ), .C2(_05530_ ), .ZN(_05531_ ) );
OR3_X1 _13214_ ( .A1(_05022_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_04913_ ), .ZN(_05532_ ) );
NAND3_X1 _13215_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_05210_ ), .ZN(_05533_ ) );
NAND2_X1 _13216_ ( .A1(_04903_ ), .A2(\mtvec [25] ), .ZN(_05534_ ) );
NAND3_X1 _13217_ ( .A1(_05049_ ), .A2(\mepc [25] ), .A3(_05076_ ), .ZN(_05535_ ) );
NAND4_X1 _13218_ ( .A1(_04842_ ), .A2(_04833_ ), .A3(_04846_ ), .A4(\mycsreg.CSReg[0][25] ), .ZN(_05536_ ) );
AND4_X1 _13219_ ( .A1(_05533_ ), .A2(_05534_ ), .A3(_05535_ ), .A4(_05536_ ), .ZN(_05537_ ) );
OAI21_X1 _13220_ ( .A(_05537_ ), .B1(_04888_ ), .B2(_05216_ ), .ZN(_05538_ ) );
NAND2_X1 _13221_ ( .A1(_05532_ ), .A2(_05538_ ), .ZN(_05539_ ) );
AOI21_X1 _13222_ ( .A(_02421_ ), .B1(_05539_ ), .B2(fanout_net_6 ), .ZN(_05540_ ) );
AND2_X1 _13223_ ( .A1(_05531_ ), .A2(_05540_ ), .ZN(_05541_ ) );
AOI211_X1 _13224_ ( .A(fanout_net_16 ), .B(_02392_ ), .C1(_02408_ ), .C2(_05270_ ), .ZN(_05542_ ) );
OAI21_X1 _13225_ ( .A(_05453_ ), .B1(_05541_ ), .B2(_05542_ ), .ZN(_05543_ ) );
NOR2_X1 _13226_ ( .A1(_03390_ ), .A2(_05250_ ), .ZN(_05544_ ) );
NOR2_X1 _13227_ ( .A1(_05530_ ), .A2(_02420_ ), .ZN(_05545_ ) );
NOR3_X1 _13228_ ( .A1(_05544_ ), .A2(_03406_ ), .A3(_05545_ ), .ZN(_05546_ ) );
NAND3_X1 _13229_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [25] ), .ZN(_05547_ ) );
AOI22_X1 _13230_ ( .A1(_05543_ ), .A2(_05546_ ), .B1(_05410_ ), .B2(_05547_ ), .ZN(_00149_ ) );
NAND3_X1 _13231_ ( .A1(_05049_ ), .A2(\mepc [24] ), .A3(_04898_ ), .ZN(_05548_ ) );
NAND4_X1 _13232_ ( .A1(_04895_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][24] ), .A4(_05052_ ), .ZN(_05549_ ) );
NAND4_X1 _13233_ ( .A1(_05054_ ), .A2(\mtvec [24] ), .A3(_05052_ ), .A4(_05127_ ), .ZN(_05550_ ) );
NAND4_X1 _13234_ ( .A1(_04837_ ), .A2(_05548_ ), .A3(_05549_ ), .A4(_05550_ ), .ZN(_05551_ ) );
AND4_X1 _13235_ ( .A1(\mycsreg.CSReg[0][24] ), .A2(_05190_ ), .A3(_04898_ ), .A4(_04988_ ), .ZN(_05552_ ) );
OAI22_X1 _13236_ ( .A1(_03540_ ), .A2(_03542_ ), .B1(_05551_ ), .B2(_05552_ ), .ZN(_05553_ ) );
NAND3_X1 _13237_ ( .A1(_04849_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_04998_ ), .ZN(_05554_ ) );
AOI21_X1 _13238_ ( .A(_04853_ ), .B1(_05553_ ), .B2(_05554_ ), .ZN(_05555_ ) );
XNOR2_X1 _13239_ ( .A(_05521_ ), .B(\ID_EX_pc [24] ), .ZN(_05556_ ) );
XOR2_X1 _13240_ ( .A(_05527_ ), .B(_03408_ ), .Z(_05557_ ) );
MUX2_X1 _13241_ ( .A(_05556_ ), .B(_05557_ ), .S(_04778_ ), .Z(_05558_ ) );
AOI21_X1 _13242_ ( .A(_05555_ ), .B1(_05558_ ), .B2(_04860_ ), .ZN(_05559_ ) );
NOR2_X1 _13243_ ( .A1(_05559_ ), .A2(_04862_ ), .ZN(_05560_ ) );
INV_X1 _13244_ ( .A(\myexu.pc_jump [24] ), .ZN(_05561_ ) );
AOI211_X1 _13245_ ( .A(fanout_net_16 ), .B(_05561_ ), .C1(_02408_ ), .C2(_05270_ ), .ZN(_05562_ ) );
OAI21_X1 _13246_ ( .A(_05453_ ), .B1(_05560_ ), .B2(_05562_ ), .ZN(_05563_ ) );
NOR2_X1 _13247_ ( .A1(_03391_ ), .A2(_05250_ ), .ZN(_05564_ ) );
AND3_X1 _13248_ ( .A1(_05557_ ), .A2(_05305_ ), .A3(_03517_ ), .ZN(_05565_ ) );
NOR3_X1 _13249_ ( .A1(_05564_ ), .A2(_03406_ ), .A3(_05565_ ), .ZN(_05566_ ) );
NAND3_X1 _13250_ ( .A1(_05356_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [24] ), .ZN(_05567_ ) );
AOI22_X1 _13251_ ( .A1(_05563_ ), .A2(_05566_ ), .B1(_05410_ ), .B2(_05567_ ), .ZN(_00150_ ) );
NAND3_X1 _13252_ ( .A1(_04812_ ), .A2(\ID_EX_pc [22] ), .A3(_05519_ ), .ZN(_05568_ ) );
XNOR2_X1 _13253_ ( .A(_05568_ ), .B(\ID_EX_pc [23] ), .ZN(_05569_ ) );
AND2_X2 _13254_ ( .A1(_04875_ ), .A2(_05569_ ), .ZN(_05570_ ) );
INV_X1 _13255_ ( .A(_03483_ ), .ZN(_05571_ ) );
OAI21_X1 _13256_ ( .A(_03487_ ), .B1(_03472_ ), .B2(_03480_ ), .ZN(_05572_ ) );
AOI21_X1 _13257_ ( .A(_05571_ ), .B1(_05572_ ), .B2(_03493_ ), .ZN(_05573_ ) );
NOR2_X1 _13258_ ( .A1(_05573_ ), .A2(_03489_ ), .ZN(_05574_ ) );
XNOR2_X1 _13259_ ( .A(_05574_ ), .B(_03482_ ), .ZN(_05575_ ) );
AOI211_X1 _13260_ ( .A(fanout_net_6 ), .B(_05570_ ), .C1(_04858_ ), .C2(_05575_ ), .ZN(_05576_ ) );
OR3_X1 _13261_ ( .A1(_04888_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_04890_ ), .ZN(_05577_ ) );
NAND3_X1 _13262_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_04984_ ), .ZN(_05578_ ) );
NAND2_X1 _13263_ ( .A1(_04903_ ), .A2(\mtvec [23] ), .ZN(_05579_ ) );
NAND3_X1 _13264_ ( .A1(_05049_ ), .A2(\mepc [23] ), .A3(_04898_ ), .ZN(_05580_ ) );
NAND4_X1 _13265_ ( .A1(_05190_ ), .A2(_05052_ ), .A3(_05056_ ), .A4(\mycsreg.CSReg[0][23] ), .ZN(_05581_ ) );
AND4_X1 _13266_ ( .A1(_05578_ ), .A2(_05579_ ), .A3(_05580_ ), .A4(_05581_ ), .ZN(_05582_ ) );
BUF_X2 _13267_ ( .A(_05022_ ), .Z(_05583_ ) );
OAI21_X1 _13268_ ( .A(_05582_ ), .B1(_05583_ ), .B2(_04914_ ), .ZN(_05584_ ) );
NAND2_X1 _13269_ ( .A1(_05577_ ), .A2(_05584_ ), .ZN(_05585_ ) );
AOI211_X1 _13270_ ( .A(_02421_ ), .B(_05576_ ), .C1(fanout_net_6 ), .C2(_05585_ ), .ZN(_05586_ ) );
INV_X1 _13271_ ( .A(\myexu.pc_jump [23] ), .ZN(_05587_ ) );
AOI211_X1 _13272_ ( .A(fanout_net_16 ), .B(_05587_ ), .C1(_02408_ ), .C2(_05270_ ), .ZN(_05588_ ) );
OAI21_X1 _13273_ ( .A(_05453_ ), .B1(_05586_ ), .B2(_05588_ ), .ZN(_05589_ ) );
OAI21_X1 _13274_ ( .A(_05088_ ), .B1(_03396_ ), .B2(_03397_ ), .ZN(_05590_ ) );
NAND3_X1 _13275_ ( .A1(_05575_ ), .A2(_04785_ ), .A3(_05180_ ), .ZN(_05591_ ) );
AND3_X1 _13276_ ( .A1(_05590_ ), .A2(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_05591_ ), .ZN(_05592_ ) );
NAND3_X1 _13277_ ( .A1(_01886_ ), .A2(_05381_ ), .A3(\myexu.pc_jump [23] ), .ZN(_05593_ ) );
AOI22_X1 _13278_ ( .A1(_05589_ ), .A2(_05592_ ), .B1(_05410_ ), .B2(_05593_ ), .ZN(_00151_ ) );
NAND3_X1 _13279_ ( .A1(_05015_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_04798_ ), .ZN(_05594_ ) );
NAND3_X1 _13280_ ( .A1(_03557_ ), .A2(\mepc [22] ), .A3(_04844_ ), .ZN(_05595_ ) );
NAND2_X1 _13281_ ( .A1(_04903_ ), .A2(\mtvec [22] ), .ZN(_05596_ ) );
NAND4_X1 _13282_ ( .A1(_05014_ ), .A2(_05594_ ), .A3(_05595_ ), .A4(_05596_ ), .ZN(_05597_ ) );
NAND4_X1 _13283_ ( .A1(_04842_ ), .A2(_04844_ ), .A3(_04846_ ), .A4(\mycsreg.CSReg[0][22] ), .ZN(_05598_ ) );
OAI21_X1 _13284_ ( .A(_05598_ ), .B1(_04887_ ), .B2(_04889_ ), .ZN(_05599_ ) );
NOR2_X1 _13285_ ( .A1(_05597_ ), .A2(_05599_ ), .ZN(_05600_ ) );
NOR3_X1 _13286_ ( .A1(_04887_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_04889_ ), .ZN(_05601_ ) );
NOR2_X1 _13287_ ( .A1(_05600_ ), .A2(_05601_ ), .ZN(_05602_ ) );
OAI21_X1 _13288_ ( .A(_02411_ ), .B1(_05602_ ), .B2(_04853_ ), .ZN(_05603_ ) );
XNOR2_X1 _13289_ ( .A(_05520_ ), .B(\ID_EX_pc [22] ), .ZN(_05604_ ) );
NAND2_X1 _13290_ ( .A1(_05572_ ), .A2(_03493_ ), .ZN(_05605_ ) );
XNOR2_X1 _13291_ ( .A(_05605_ ), .B(_05571_ ), .ZN(_05606_ ) );
INV_X1 _13292_ ( .A(_05606_ ), .ZN(_05607_ ) );
MUX2_X1 _13293_ ( .A(_05604_ ), .B(_05607_ ), .S(_04858_ ), .Z(_05608_ ) );
AOI21_X1 _13294_ ( .A(_05603_ ), .B1(_05608_ ), .B2(_04860_ ), .ZN(_05609_ ) );
AND3_X1 _13295_ ( .A1(_04874_ ), .A2(_03401_ ), .A3(\myexu.pc_jump [22] ), .ZN(_05610_ ) );
OAI21_X1 _13296_ ( .A(_05453_ ), .B1(_05609_ ), .B2(_05610_ ), .ZN(_05611_ ) );
NAND3_X1 _13297_ ( .A1(_03399_ ), .A2(_05088_ ), .A3(_03393_ ), .ZN(_05612_ ) );
NAND3_X1 _13298_ ( .A1(_05606_ ), .A2(_04785_ ), .A3(_05180_ ), .ZN(_05613_ ) );
AND3_X1 _13299_ ( .A1(_05612_ ), .A2(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_05613_ ), .ZN(_05614_ ) );
NAND3_X1 _13300_ ( .A1(_01886_ ), .A2(_03402_ ), .A3(\myexu.pc_jump [22] ), .ZN(_05615_ ) );
AOI22_X1 _13301_ ( .A1(_05611_ ), .A2(_05614_ ), .B1(_05410_ ), .B2(_05615_ ), .ZN(_00152_ ) );
OAI21_X1 _13302_ ( .A(_03486_ ), .B1(_03472_ ), .B2(_03480_ ), .ZN(_05616_ ) );
NAND2_X1 _13303_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_05617_ ) );
NAND2_X1 _13304_ ( .A1(_05616_ ), .A2(_05617_ ), .ZN(_05618_ ) );
XNOR2_X1 _13305_ ( .A(_05618_ ), .B(_03485_ ), .ZN(_05619_ ) );
NAND3_X1 _13306_ ( .A1(_04775_ ), .A2(_04776_ ), .A3(_05619_ ), .ZN(_05620_ ) );
INV_X1 _13307_ ( .A(\ID_EX_pc [20] ), .ZN(_05621_ ) );
NOR2_X1 _13308_ ( .A1(_04855_ ), .A2(_05621_ ), .ZN(_05622_ ) );
INV_X1 _13309_ ( .A(\ID_EX_pc [21] ), .ZN(_05623_ ) );
XNOR2_X1 _13310_ ( .A(_05622_ ), .B(_05623_ ), .ZN(_05624_ ) );
OAI211_X1 _13311_ ( .A(_04978_ ), .B(_05620_ ), .C1(_04879_ ), .C2(_05624_ ), .ZN(_05625_ ) );
AND3_X1 _13312_ ( .A1(_04996_ ), .A2(\EX_LS_result_csreg_mem [21] ), .A3(_04995_ ), .ZN(_05626_ ) );
NAND3_X1 _13313_ ( .A1(_05049_ ), .A2(\mepc [21] ), .A3(_05055_ ), .ZN(_05627_ ) );
NAND4_X1 _13314_ ( .A1(_05210_ ), .A2(_05051_ ), .A3(\mycsreg.CSReg[3][21] ), .A4(_05055_ ), .ZN(_05628_ ) );
NAND4_X1 _13315_ ( .A1(_04940_ ), .A2(\mtvec [21] ), .A3(_05055_ ), .A4(_05056_ ), .ZN(_05629_ ) );
AND4_X1 _13316_ ( .A1(_03552_ ), .A2(_05627_ ), .A3(_05628_ ), .A4(_05629_ ), .ZN(_05630_ ) );
NAND4_X1 _13317_ ( .A1(_05059_ ), .A2(_04899_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][21] ), .ZN(_05631_ ) );
AOI22_X1 _13318_ ( .A1(_05046_ ), .A2(_05048_ ), .B1(_05630_ ), .B2(_05631_ ), .ZN(_05632_ ) );
OAI21_X1 _13319_ ( .A(fanout_net_6 ), .B1(_05626_ ), .B2(_05632_ ), .ZN(_05633_ ) );
AOI21_X1 _13320_ ( .A(_04864_ ), .B1(_05625_ ), .B2(_05633_ ), .ZN(_05634_ ) );
INV_X1 _13321_ ( .A(\myexu.pc_jump [21] ), .ZN(_05635_ ) );
AOI211_X1 _13322_ ( .A(fanout_net_16 ), .B(_05635_ ), .C1(_02408_ ), .C2(_02409_ ), .ZN(_05636_ ) );
OAI21_X1 _13323_ ( .A(_05453_ ), .B1(_05634_ ), .B2(_05636_ ), .ZN(_05637_ ) );
NOR2_X1 _13324_ ( .A1(_03354_ ), .A2(_05250_ ), .ZN(_05638_ ) );
NOR2_X1 _13325_ ( .A1(_05619_ ), .A2(_02420_ ), .ZN(_05639_ ) );
NOR3_X1 _13326_ ( .A1(_05638_ ), .A2(_03406_ ), .A3(_05639_ ), .ZN(_05640_ ) );
NAND3_X1 _13327_ ( .A1(_01886_ ), .A2(_03402_ ), .A3(\myexu.pc_jump [21] ), .ZN(_05641_ ) );
AOI22_X1 _13328_ ( .A1(_05637_ ), .A2(_05640_ ), .B1(_04787_ ), .B2(_05641_ ), .ZN(_00153_ ) );
OAI21_X1 _13329_ ( .A(_03514_ ), .B1(_03511_ ), .B2(_03512_ ), .ZN(_05642_ ) );
NAND2_X1 _13330_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_05643_ ) );
NAND2_X1 _13331_ ( .A1(_05642_ ), .A2(_05643_ ), .ZN(_05644_ ) );
XNOR2_X1 _13332_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_05645_ ) );
XNOR2_X1 _13333_ ( .A(_05644_ ), .B(_05645_ ), .ZN(_05646_ ) );
OAI21_X1 _13334_ ( .A(_03517_ ), .B1(_05646_ ), .B2(fanout_net_5 ), .ZN(_05647_ ) );
AOI21_X1 _13335_ ( .A(_05647_ ), .B1(_03339_ ), .B2(fanout_net_5 ), .ZN(_05648_ ) );
NAND2_X1 _13336_ ( .A1(_03401_ ), .A2(_02394_ ), .ZN(_05649_ ) );
NAND3_X1 _13337_ ( .A1(_03557_ ), .A2(\mepc [31] ), .A3(_04833_ ), .ZN(_05650_ ) );
NAND4_X1 _13338_ ( .A1(_03569_ ), .A2(\mtvec [31] ), .A3(_04844_ ), .A4(_04846_ ), .ZN(_05651_ ) );
NAND4_X1 _13339_ ( .A1(_04838_ ), .A2(_04799_ ), .A3(\mycsreg.CSReg[3][31] ), .A4(_04796_ ), .ZN(_05652_ ) );
NAND4_X1 _13340_ ( .A1(_04842_ ), .A2(_04844_ ), .A3(_03574_ ), .A4(\mycsreg.CSReg[0][31] ), .ZN(_05653_ ) );
NAND4_X1 _13341_ ( .A1(_05650_ ), .A2(_05651_ ), .A3(_05652_ ), .A4(_05653_ ), .ZN(_05654_ ) );
OAI21_X1 _13342_ ( .A(_05654_ ), .B1(_03540_ ), .B2(_03542_ ), .ZN(_05655_ ) );
NAND3_X1 _13343_ ( .A1(_03539_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_03577_ ), .ZN(_05656_ ) );
NAND2_X1 _13344_ ( .A1(_05655_ ), .A2(_05656_ ), .ZN(_05657_ ) );
NOR2_X1 _13345_ ( .A1(_03598_ ), .A2(_03599_ ), .ZN(_05658_ ) );
XNOR2_X1 _13346_ ( .A(_05658_ ), .B(_03404_ ), .ZN(_05659_ ) );
MUX2_X1 _13347_ ( .A(_05659_ ), .B(_05646_ ), .S(_04777_ ), .Z(_05660_ ) );
MUX2_X1 _13348_ ( .A(_05657_ ), .B(_05660_ ), .S(_03580_ ), .Z(_05661_ ) );
MUX2_X2 _13349_ ( .A(_05649_ ), .B(_05661_ ), .S(_02411_ ), .Z(_05662_ ) );
BUF_X4 _13350_ ( .A(_04831_ ), .Z(_05663_ ) );
AOI21_X1 _13351_ ( .A(_05648_ ), .B1(_05662_ ), .B2(_05663_ ), .ZN(_05664_ ) );
NOR3_X1 _13352_ ( .A1(fanout_net_2 ), .A2(fanout_net_16 ), .A3(\myexu.pc_jump [31] ), .ZN(_05665_ ) );
OAI22_X1 _13353_ ( .A1(_05664_ ), .A2(_04868_ ), .B1(\myidu.state_$_ANDNOT__A_Y ), .B2(_05665_ ), .ZN(_00154_ ) );
NOR3_X1 _13354_ ( .A1(_03599_ ), .A2(fanout_net_2 ), .A3(fanout_net_16 ), .ZN(_00155_ ) );
NOR3_X1 _13355_ ( .A1(_05623_ ), .A2(fanout_net_2 ), .A3(fanout_net_16 ), .ZN(_00156_ ) );
NOR3_X1 _13356_ ( .A1(_05621_ ), .A2(fanout_net_2 ), .A3(fanout_net_16 ), .ZN(_00157_ ) );
INV_X1 _13357_ ( .A(\ID_EX_pc [19] ), .ZN(_05666_ ) );
NOR3_X1 _13358_ ( .A1(_05666_ ), .A2(fanout_net_2 ), .A3(fanout_net_16 ), .ZN(_00158_ ) );
INV_X1 _13359_ ( .A(\ID_EX_pc [18] ), .ZN(_05667_ ) );
NOR3_X1 _13360_ ( .A1(_05667_ ), .A2(fanout_net_2 ), .A3(fanout_net_16 ), .ZN(_00159_ ) );
AND3_X1 _13361_ ( .A1(_01914_ ), .A2(_03403_ ), .A3(\ID_EX_pc [17] ), .ZN(_00160_ ) );
NOR3_X1 _13362_ ( .A1(_04974_ ), .A2(fanout_net_2 ), .A3(fanout_net_16 ), .ZN(_00161_ ) );
NOR3_X1 _13363_ ( .A1(_05037_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00162_ ) );
NOR3_X1 _13364_ ( .A1(_05035_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00163_ ) );
AND3_X1 _13365_ ( .A1(_01914_ ), .A2(_03403_ ), .A3(\ID_EX_pc [13] ), .ZN(_00164_ ) );
NOR3_X1 _13366_ ( .A1(_05095_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00165_ ) );
NOR3_X1 _13367_ ( .A1(_03510_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00166_ ) );
NOR3_X1 _13368_ ( .A1(_05149_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00167_ ) );
NOR3_X1 _13369_ ( .A1(_05202_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00168_ ) );
INV_X1 _13370_ ( .A(\ID_EX_pc [9] ), .ZN(_05668_ ) );
NOR3_X1 _13371_ ( .A1(_05668_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00169_ ) );
NOR3_X1 _13372_ ( .A1(_05263_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00170_ ) );
NOR3_X1 _13373_ ( .A1(_05294_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00171_ ) );
NOR3_X1 _13374_ ( .A1(_05317_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00172_ ) );
AND3_X1 _13375_ ( .A1(_01914_ ), .A2(_03403_ ), .A3(\ID_EX_pc [5] ), .ZN(_00173_ ) );
AND3_X1 _13376_ ( .A1(_01914_ ), .A2(_03403_ ), .A3(\ID_EX_pc [4] ), .ZN(_00174_ ) );
AND3_X1 _13377_ ( .A1(_01914_ ), .A2(_03403_ ), .A3(\ID_EX_pc [3] ), .ZN(_00175_ ) );
INV_X1 _13378_ ( .A(\ID_EX_pc [2] ), .ZN(_05669_ ) );
NOR3_X1 _13379_ ( .A1(_05669_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00176_ ) );
NOR3_X1 _13380_ ( .A1(_05181_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00177_ ) );
INV_X1 _13381_ ( .A(\ID_EX_pc [1] ), .ZN(_05670_ ) );
NOR3_X1 _13382_ ( .A1(_05670_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00178_ ) );
NOR3_X1 _13383_ ( .A1(_05488_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00179_ ) );
NOR3_X1 _13384_ ( .A1(_04817_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00180_ ) );
NOR3_X1 _13385_ ( .A1(_04818_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00181_ ) );
NOR3_X1 _13386_ ( .A1(_05524_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00182_ ) );
NOR3_X1 _13387_ ( .A1(_05522_ ), .A2(fanout_net_2 ), .A3(excp_written ), .ZN(_00183_ ) );
INV_X1 _13388_ ( .A(\ID_EX_pc [23] ), .ZN(_05671_ ) );
NOR3_X1 _13389_ ( .A1(_05671_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00184_ ) );
AND3_X1 _13390_ ( .A1(_01914_ ), .A2(_04789_ ), .A3(\ID_EX_pc [22] ), .ZN(_00185_ ) );
BUF_X4 _13391_ ( .A(_02406_ ), .Z(_05672_ ) );
NOR3_X1 _13392_ ( .A1(_05672_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00186_ ) );
AND3_X1 _13393_ ( .A1(_02296_ ), .A2(\myclint.rvalid ), .A3(_02316_ ), .ZN(_05673_ ) );
INV_X1 _13394_ ( .A(_05673_ ), .ZN(_05674_ ) );
OAI21_X1 _13395_ ( .A(_05674_ ), .B1(_02317_ ), .B2(io_master_arready ), .ZN(_05675_ ) );
INV_X2 _13396_ ( .A(_02270_ ), .ZN(_05676_ ) );
NOR2_X1 _13397_ ( .A1(_05675_ ), .A2(_05676_ ), .ZN(_05677_ ) );
BUF_X2 _13398_ ( .A(_02272_ ), .Z(_05678_ ) );
BUF_X4 _13399_ ( .A(_02327_ ), .Z(_05679_ ) );
INV_X1 _13400_ ( .A(_05679_ ), .ZN(_05680_ ) );
OR3_X1 _13401_ ( .A1(_05677_ ), .A2(_05678_ ), .A3(_05680_ ), .ZN(_05681_ ) );
OR2_X1 _13402_ ( .A1(\mylsu.state [0] ), .A2(\mylsu.state [4] ), .ZN(_05682_ ) );
INV_X1 _13403_ ( .A(_02346_ ), .ZN(_05683_ ) );
OAI21_X1 _13404_ ( .A(_05682_ ), .B1(_05683_ ), .B2(io_master_awready ), .ZN(_05684_ ) );
AOI21_X1 _13405_ ( .A(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .B1(_05684_ ), .B2(EXU_valid_LSU ), .ZN(_05685_ ) );
AOI21_X1 _13406_ ( .A(_02404_ ), .B1(_05681_ ), .B2(_05685_ ), .ZN(_00187_ ) );
NOR3_X1 _13407_ ( .A1(_04920_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00188_ ) );
NOR3_X1 _13408_ ( .A1(_02412_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00189_ ) );
NOR3_X1 _13409_ ( .A1(_04511_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00190_ ) );
NOR3_X1 _13410_ ( .A1(_04860_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00191_ ) );
BUF_X4 _13411_ ( .A(_04771_ ), .Z(_05686_ ) );
NOR3_X1 _13412_ ( .A1(_05686_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00192_ ) );
NOR3_X1 _13413_ ( .A1(_04417_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00193_ ) );
BUF_X4 _13414_ ( .A(_04869_ ), .Z(_05687_ ) );
NOR3_X1 _13415_ ( .A1(_05687_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00194_ ) );
AND2_X1 _13416_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_05688_ ) );
NOR2_X1 _13417_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_05689_ ) );
AND2_X1 _13418_ ( .A1(_05688_ ), .A2(_05689_ ), .ZN(_05690_ ) );
CLKBUF_X2 _13419_ ( .A(_05690_ ), .Z(_05691_ ) );
BUF_X2 _13420_ ( .A(_05691_ ), .Z(_05692_ ) );
AND3_X2 _13421_ ( .A1(_05692_ ), .A2(\IF_ID_inst [12] ), .A3(\IF_ID_inst [6] ), .ZN(_05693_ ) );
AND2_X2 _13422_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05694_ ) );
AND2_X1 _13423_ ( .A1(_05693_ ), .A2(_05694_ ), .ZN(_05695_ ) );
INV_X1 _13424_ ( .A(\IF_ID_inst [6] ), .ZN(_05696_ ) );
NOR2_X1 _13425_ ( .A1(_05696_ ), .A2(\IF_ID_inst [12] ), .ZN(_05697_ ) );
AND3_X1 _13426_ ( .A1(_05697_ ), .A2(\IF_ID_inst [13] ), .A3(_05694_ ), .ZN(_05698_ ) );
AND2_X1 _13427_ ( .A1(_05698_ ), .A2(_05692_ ), .ZN(_05699_ ) );
NOR2_X2 _13428_ ( .A1(_05695_ ), .A2(_05699_ ), .ZN(_05700_ ) );
BUF_X4 _13429_ ( .A(_05700_ ), .Z(_05701_ ) );
INV_X1 _13430_ ( .A(\IF_ID_inst [31] ), .ZN(_05702_ ) );
AND2_X2 _13431_ ( .A1(_02388_ ), .A2(_02403_ ), .ZN(_05703_ ) );
INV_X2 _13432_ ( .A(_05703_ ), .ZN(_05704_ ) );
BUF_X4 _13433_ ( .A(_05704_ ), .Z(_05705_ ) );
NOR3_X1 _13434_ ( .A1(_05701_ ), .A2(_05702_ ), .A3(_05705_ ), .ZN(_00195_ ) );
INV_X1 _13435_ ( .A(\IF_ID_inst [30] ), .ZN(_05706_ ) );
NOR3_X1 _13436_ ( .A1(_05701_ ), .A2(_05706_ ), .A3(_05705_ ), .ZN(_00196_ ) );
INV_X1 _13437_ ( .A(\IF_ID_inst [21] ), .ZN(_05707_ ) );
NOR3_X1 _13438_ ( .A1(_05701_ ), .A2(_05707_ ), .A3(_05705_ ), .ZN(_00197_ ) );
BUF_X4 _13439_ ( .A(_05704_ ), .Z(_05708_ ) );
INV_X1 _13440_ ( .A(_05700_ ), .ZN(_05709_ ) );
INV_X1 _13441_ ( .A(\IF_ID_inst [20] ), .ZN(_05710_ ) );
AOI21_X1 _13442_ ( .A(_05708_ ), .B1(_05709_ ), .B2(_05710_ ), .ZN(_00198_ ) );
INV_X1 _13443_ ( .A(\IF_ID_inst [29] ), .ZN(_05711_ ) );
AOI21_X1 _13444_ ( .A(_05708_ ), .B1(_05709_ ), .B2(_05711_ ), .ZN(_00199_ ) );
INV_X1 _13445_ ( .A(\IF_ID_inst [28] ), .ZN(_05712_ ) );
AOI21_X1 _13446_ ( .A(_05708_ ), .B1(_05709_ ), .B2(_05712_ ), .ZN(_00200_ ) );
INV_X1 _13447_ ( .A(\IF_ID_inst [27] ), .ZN(_05713_ ) );
NOR3_X1 _13448_ ( .A1(_05701_ ), .A2(_05713_ ), .A3(_05705_ ), .ZN(_00201_ ) );
INV_X1 _13449_ ( .A(\IF_ID_inst [26] ), .ZN(_05714_ ) );
AOI21_X1 _13450_ ( .A(_05708_ ), .B1(_05709_ ), .B2(_05714_ ), .ZN(_00202_ ) );
INV_X1 _13451_ ( .A(\IF_ID_inst [25] ), .ZN(_05715_ ) );
NOR3_X1 _13452_ ( .A1(_05701_ ), .A2(_05715_ ), .A3(_05705_ ), .ZN(_00203_ ) );
INV_X1 _13453_ ( .A(\IF_ID_inst [24] ), .ZN(_05716_ ) );
NOR3_X1 _13454_ ( .A1(_05701_ ), .A2(_05716_ ), .A3(_05705_ ), .ZN(_00204_ ) );
INV_X1 _13455_ ( .A(\IF_ID_inst [23] ), .ZN(_05717_ ) );
BUF_X4 _13456_ ( .A(_05704_ ), .Z(_05718_ ) );
NOR3_X1 _13457_ ( .A1(_05701_ ), .A2(_05717_ ), .A3(_05718_ ), .ZN(_00205_ ) );
INV_X1 _13458_ ( .A(\IF_ID_inst [22] ), .ZN(_05719_ ) );
NOR3_X1 _13459_ ( .A1(_05701_ ), .A2(_05719_ ), .A3(_05718_ ), .ZN(_00206_ ) );
AND3_X1 _13460_ ( .A1(_02388_ ), .A2(_02403_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00207_ ) );
AND3_X1 _13461_ ( .A1(_02388_ ), .A2(_02403_ ), .A3(\myidu.state [2] ), .ZN(_00208_ ) );
NOR2_X1 _13462_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_05720_ ) );
NOR2_X1 _13463_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05721_ ) );
AND4_X1 _13464_ ( .A1(\IF_ID_inst [12] ), .A2(_05720_ ), .A3(_05721_ ), .A4(_05696_ ), .ZN(_05722_ ) );
AND3_X2 _13465_ ( .A1(_05688_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_05723_ ) );
CLKBUF_X2 _13466_ ( .A(_05723_ ), .Z(_05724_ ) );
AND2_X1 _13467_ ( .A1(_05722_ ), .A2(_05724_ ), .ZN(_05725_ ) );
INV_X1 _13468_ ( .A(\IF_ID_inst [7] ), .ZN(_05726_ ) );
AND4_X1 _13469_ ( .A1(\IF_ID_inst [6] ), .A2(_05691_ ), .A3(_05726_ ), .A4(_05694_ ), .ZN(_05727_ ) );
OR3_X1 _13470_ ( .A1(\IF_ID_inst [11] ), .A2(\IF_ID_inst [10] ), .A3(\IF_ID_inst [9] ), .ZN(_05728_ ) );
NOR2_X1 _13471_ ( .A1(_05728_ ), .A2(\IF_ID_inst [8] ), .ZN(_05729_ ) );
NOR4_X1 _13472_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_05730_ ) );
AND3_X1 _13473_ ( .A1(_05727_ ), .A2(_05729_ ), .A3(_05730_ ), .ZN(_05731_ ) );
NOR2_X1 _13474_ ( .A1(\IF_ID_inst [18] ), .A2(\IF_ID_inst [17] ), .ZN(_05732_ ) );
NOR2_X1 _13475_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [16] ), .ZN(_05733_ ) );
AND2_X1 _13476_ ( .A1(_05732_ ), .A2(_05733_ ), .ZN(_05734_ ) );
NOR2_X1 _13477_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_05735_ ) );
NAND4_X1 _13478_ ( .A1(_05734_ ), .A2(_05707_ ), .A3(\IF_ID_inst [20] ), .A4(_05735_ ), .ZN(_05736_ ) );
NOR3_X1 _13479_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .A3(\IF_ID_inst [24] ), .ZN(_05737_ ) );
NAND2_X1 _13480_ ( .A1(_05737_ ), .A2(_05713_ ), .ZN(_05738_ ) );
NAND4_X1 _13481_ ( .A1(_05706_ ), .A2(_05711_ ), .A3(_05712_ ), .A4(_05702_ ), .ZN(_05739_ ) );
NOR3_X1 _13482_ ( .A1(_05736_ ), .A2(_05738_ ), .A3(_05739_ ), .ZN(_05740_ ) );
AOI21_X1 _13483_ ( .A(_05725_ ), .B1(_05731_ ), .B2(_05740_ ), .ZN(_05741_ ) );
INV_X1 _13484_ ( .A(\IF_ID_inst [5] ), .ZN(_05742_ ) );
NOR2_X1 _13485_ ( .A1(_05742_ ), .A2(\IF_ID_inst [4] ), .ZN(_05743_ ) );
CLKBUF_X2 _13486_ ( .A(_05743_ ), .Z(_05744_ ) );
NOR2_X1 _13487_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_05745_ ) );
AND3_X1 _13488_ ( .A1(_05691_ ), .A2(_05744_ ), .A3(_05745_ ), .ZN(_05746_ ) );
BUF_X2 _13489_ ( .A(_05720_ ), .Z(_05747_ ) );
NAND2_X1 _13490_ ( .A1(_05746_ ), .A2(_05747_ ), .ZN(_05748_ ) );
INV_X1 _13491_ ( .A(\IF_ID_inst [12] ), .ZN(_05749_ ) );
NOR2_X1 _13492_ ( .A1(_05749_ ), .A2(\IF_ID_inst [6] ), .ZN(_05750_ ) );
AND3_X1 _13493_ ( .A1(_05750_ ), .A2(_05688_ ), .A3(_05689_ ), .ZN(_05751_ ) );
NAND3_X1 _13494_ ( .A1(_05751_ ), .A2(_05747_ ), .A3(_05744_ ), .ZN(_05752_ ) );
AND2_X1 _13495_ ( .A1(_05748_ ), .A2(_05752_ ), .ZN(_05753_ ) );
INV_X1 _13496_ ( .A(\IF_ID_inst [13] ), .ZN(_05754_ ) );
NOR2_X1 _13497_ ( .A1(_05754_ ), .A2(\IF_ID_inst [14] ), .ZN(_05755_ ) );
AND2_X1 _13498_ ( .A1(_05746_ ), .A2(_05755_ ), .ZN(_05756_ ) );
INV_X1 _13499_ ( .A(_05756_ ), .ZN(_05757_ ) );
AND3_X1 _13500_ ( .A1(_05741_ ), .A2(_05753_ ), .A3(_05757_ ), .ZN(_05758_ ) );
CLKBUF_X2 _13501_ ( .A(_05703_ ), .Z(_05759_ ) );
INV_X1 _13502_ ( .A(\IF_ID_inst [15] ), .ZN(_05760_ ) );
AND4_X1 _13503_ ( .A1(_05749_ ), .A2(_05726_ ), .A3(_05760_ ), .A4(\IF_ID_inst [6] ), .ZN(_05761_ ) );
AND3_X1 _13504_ ( .A1(_05761_ ), .A2(_05694_ ), .A3(_05720_ ), .ZN(_05762_ ) );
NAND3_X1 _13505_ ( .A1(_05762_ ), .A2(_05692_ ), .A3(_05729_ ), .ZN(_05763_ ) );
INV_X1 _13506_ ( .A(_05763_ ), .ZN(_05764_ ) );
AND4_X1 _13507_ ( .A1(\IF_ID_inst [21] ), .A2(_05706_ ), .A3(_05702_ ), .A4(\IF_ID_inst [28] ), .ZN(_05765_ ) );
NAND4_X1 _13508_ ( .A1(_05765_ ), .A2(_05710_ ), .A3(\IF_ID_inst [29] ), .A4(_05735_ ), .ZN(_05766_ ) );
INV_X1 _13509_ ( .A(_05734_ ), .ZN(_05767_ ) );
NOR3_X1 _13510_ ( .A1(_05766_ ), .A2(_05738_ ), .A3(_05767_ ), .ZN(_05768_ ) );
AND3_X1 _13511_ ( .A1(_05697_ ), .A2(_05744_ ), .A3(_05747_ ), .ZN(_05769_ ) );
AOI22_X1 _13512_ ( .A1(_05764_ ), .A2(_05768_ ), .B1(_05692_ ), .B2(_05769_ ), .ZN(_05770_ ) );
AND3_X1 _13513_ ( .A1(_05693_ ), .A2(_05754_ ), .A3(_05744_ ), .ZN(_05771_ ) );
AND2_X1 _13514_ ( .A1(_05697_ ), .A2(_05744_ ), .ZN(_05772_ ) );
AND2_X1 _13515_ ( .A1(_05772_ ), .A2(_05692_ ), .ZN(_05773_ ) );
AND2_X1 _13516_ ( .A1(_05773_ ), .A2(\IF_ID_inst [14] ), .ZN(_05774_ ) );
NOR2_X1 _13517_ ( .A1(_05771_ ), .A2(_05774_ ), .ZN(_05775_ ) );
AND2_X1 _13518_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_05776_ ) );
NAND3_X1 _13519_ ( .A1(_05693_ ), .A2(_05776_ ), .A3(_05744_ ), .ZN(_05777_ ) );
AND3_X1 _13520_ ( .A1(_05770_ ), .A2(_05775_ ), .A3(_05777_ ), .ZN(_05778_ ) );
AND4_X1 _13521_ ( .A1(\IF_ID_inst [11] ), .A2(_05758_ ), .A3(_05759_ ), .A4(_05778_ ), .ZN(_00209_ ) );
AND4_X1 _13522_ ( .A1(\IF_ID_inst [10] ), .A2(_05758_ ), .A3(_05759_ ), .A4(_05778_ ), .ZN(_00210_ ) );
AND4_X1 _13523_ ( .A1(\IF_ID_inst [9] ), .A2(_05758_ ), .A3(_05759_ ), .A4(_05778_ ), .ZN(_00211_ ) );
AND4_X1 _13524_ ( .A1(\IF_ID_inst [8] ), .A2(_05758_ ), .A3(_05759_ ), .A4(_05778_ ), .ZN(_00212_ ) );
AND4_X1 _13525_ ( .A1(\IF_ID_inst [7] ), .A2(_05758_ ), .A3(_05759_ ), .A4(_05778_ ), .ZN(_00213_ ) );
INV_X1 _13526_ ( .A(_05741_ ), .ZN(_05779_ ) );
INV_X1 _13527_ ( .A(_05743_ ), .ZN(_05780_ ) );
NOR2_X1 _13528_ ( .A1(_05780_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_05781_ ) );
AND2_X1 _13529_ ( .A1(_05781_ ), .A2(_05723_ ), .ZN(_05782_ ) );
BUF_X2 _13530_ ( .A(_05782_ ), .Z(_05783_ ) );
INV_X1 _13531_ ( .A(\IF_ID_inst [2] ), .ZN(_05784_ ) );
NOR2_X1 _13532_ ( .A1(_05784_ ), .A2(\IF_ID_inst [3] ), .ZN(_05785_ ) );
AND2_X1 _13533_ ( .A1(_05785_ ), .A2(_05688_ ), .ZN(_05786_ ) );
INV_X1 _13534_ ( .A(\IF_ID_inst [4] ), .ZN(_05787_ ) );
NOR2_X1 _13535_ ( .A1(_05787_ ), .A2(\IF_ID_inst [6] ), .ZN(_05788_ ) );
AND2_X1 _13536_ ( .A1(_05786_ ), .A2(_05788_ ), .ZN(_05789_ ) );
NOR2_X2 _13537_ ( .A1(_05783_ ), .A2(_05789_ ), .ZN(_05790_ ) );
INV_X1 _13538_ ( .A(_05768_ ), .ZN(_05791_ ) );
OAI21_X1 _13539_ ( .A(_05790_ ), .B1(_05791_ ), .B2(_05763_ ), .ZN(_05792_ ) );
INV_X1 _13540_ ( .A(\IF_ID_inst [19] ), .ZN(_05793_ ) );
NOR4_X1 _13541_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05793_ ), .A4(_05718_ ), .ZN(_00214_ ) );
INV_X1 _13542_ ( .A(\IF_ID_inst [18] ), .ZN(_05794_ ) );
NOR4_X1 _13543_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05794_ ), .A4(_05718_ ), .ZN(_00215_ ) );
INV_X1 _13544_ ( .A(\IF_ID_inst [17] ), .ZN(_05795_ ) );
NOR4_X1 _13545_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05795_ ), .A4(_05718_ ), .ZN(_00216_ ) );
AND2_X1 _13546_ ( .A1(_05753_ ), .A2(_05757_ ), .ZN(_05796_ ) );
INV_X1 _13547_ ( .A(_05796_ ), .ZN(_05797_ ) );
AND2_X1 _13548_ ( .A1(_05691_ ), .A2(_05745_ ), .ZN(_05798_ ) );
NOR2_X1 _13549_ ( .A1(_05787_ ), .A2(\IF_ID_inst [5] ), .ZN(_05799_ ) );
AND2_X1 _13550_ ( .A1(_05798_ ), .A2(_05799_ ), .ZN(_05800_ ) );
INV_X1 _13551_ ( .A(_05755_ ), .ZN(_05801_ ) );
NAND2_X1 _13552_ ( .A1(_05800_ ), .A2(_05801_ ), .ZN(_05802_ ) );
AND2_X1 _13553_ ( .A1(_05751_ ), .A2(_05799_ ), .ZN(_05803_ ) );
NAND3_X1 _13554_ ( .A1(_05803_ ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [14] ), .ZN(_05804_ ) );
AND2_X1 _13555_ ( .A1(_05802_ ), .A2(_05804_ ), .ZN(_05805_ ) );
INV_X1 _13556_ ( .A(_05805_ ), .ZN(_05806_ ) );
AND2_X1 _13557_ ( .A1(_05800_ ), .A2(_05755_ ), .ZN(_05807_ ) );
NAND3_X1 _13558_ ( .A1(_05751_ ), .A2(\IF_ID_inst [13] ), .A3(_05799_ ), .ZN(_05808_ ) );
NOR2_X1 _13559_ ( .A1(_05808_ ), .A2(\IF_ID_inst [14] ), .ZN(_05809_ ) );
OR2_X1 _13560_ ( .A1(_05807_ ), .A2(_05809_ ), .ZN(_05810_ ) );
NOR2_X1 _13561_ ( .A1(_05706_ ), .A2(\IF_ID_inst [29] ), .ZN(_05811_ ) );
NOR2_X1 _13562_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_05812_ ) );
AND3_X1 _13563_ ( .A1(_05811_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_05812_ ), .ZN(_05813_ ) );
INV_X1 _13564_ ( .A(\IF_ID_inst [14] ), .ZN(_05814_ ) );
NOR2_X1 _13565_ ( .A1(_05814_ ), .A2(\IF_ID_inst [13] ), .ZN(_05815_ ) );
NOR2_X1 _13566_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_05816_ ) );
AND2_X1 _13567_ ( .A1(_05815_ ), .A2(_05816_ ), .ZN(_05817_ ) );
AND2_X1 _13568_ ( .A1(_05813_ ), .A2(_05817_ ), .ZN(_05818_ ) );
NOR3_X1 _13569_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_05819_ ) );
AND2_X1 _13570_ ( .A1(_05819_ ), .A2(_05713_ ), .ZN(_05820_ ) );
AND4_X1 _13571_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A2(_05816_ ), .A3(_05754_ ), .A4(\IF_ID_inst [14] ), .ZN(_05821_ ) );
AND2_X1 _13572_ ( .A1(_05820_ ), .A2(_05821_ ), .ZN(_05822_ ) );
OAI21_X1 _13573_ ( .A(_05803_ ), .B1(_05818_ ), .B2(_05822_ ), .ZN(_05823_ ) );
INV_X1 _13574_ ( .A(_05823_ ), .ZN(_05824_ ) );
NOR4_X1 _13575_ ( .A1(_05797_ ), .A2(_05806_ ), .A3(_05810_ ), .A4(_05824_ ), .ZN(_05825_ ) );
AND2_X1 _13576_ ( .A1(_05798_ ), .A2(_05721_ ), .ZN(_05826_ ) );
AND2_X1 _13577_ ( .A1(_05826_ ), .A2(_05755_ ), .ZN(_05827_ ) );
AOI21_X1 _13578_ ( .A(_05827_ ), .B1(_05747_ ), .B2(_05773_ ), .ZN(_05828_ ) );
NAND3_X1 _13579_ ( .A1(_05828_ ), .A2(_05700_ ), .A3(_05775_ ), .ZN(_05829_ ) );
AND2_X1 _13580_ ( .A1(_05798_ ), .A2(_05694_ ), .ZN(_05830_ ) );
AND2_X1 _13581_ ( .A1(_05720_ ), .A2(_05816_ ), .ZN(_05831_ ) );
NAND4_X1 _13582_ ( .A1(_05831_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_05811_ ), .A4(_05812_ ), .ZN(_05832_ ) );
INV_X1 _13583_ ( .A(_05820_ ), .ZN(_05833_ ) );
NAND4_X1 _13584_ ( .A1(_05816_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(\IF_ID_inst [13] ), .A4(_05814_ ), .ZN(_05834_ ) );
OAI21_X1 _13585_ ( .A(_05832_ ), .B1(_05833_ ), .B2(_05834_ ), .ZN(_05835_ ) );
AND2_X1 _13586_ ( .A1(_05830_ ), .A2(_05835_ ), .ZN(_05836_ ) );
INV_X1 _13587_ ( .A(_05836_ ), .ZN(_05837_ ) );
AND3_X1 _13588_ ( .A1(_05819_ ), .A2(_05713_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05838_ ) );
AND2_X1 _13589_ ( .A1(_05838_ ), .A2(_05831_ ), .ZN(_05839_ ) );
AND2_X1 _13590_ ( .A1(_05839_ ), .A2(_05803_ ), .ZN(_05840_ ) );
INV_X1 _13591_ ( .A(_05840_ ), .ZN(_05841_ ) );
NAND3_X1 _13592_ ( .A1(_05798_ ), .A2(_05754_ ), .A3(_05721_ ), .ZN(_05842_ ) );
AND3_X1 _13593_ ( .A1(_05721_ ), .A2(\IF_ID_inst [12] ), .A3(_05696_ ), .ZN(_05843_ ) );
AND3_X1 _13594_ ( .A1(_05843_ ), .A2(_05692_ ), .A3(_05754_ ), .ZN(_05844_ ) );
INV_X1 _13595_ ( .A(_05844_ ), .ZN(_05845_ ) );
AND2_X1 _13596_ ( .A1(_05842_ ), .A2(_05845_ ), .ZN(_05846_ ) );
NAND3_X1 _13597_ ( .A1(_05837_ ), .A2(_05841_ ), .A3(_05846_ ), .ZN(_05847_ ) );
NOR2_X1 _13598_ ( .A1(_05829_ ), .A2(_05847_ ), .ZN(_05848_ ) );
NAND2_X1 _13599_ ( .A1(_05693_ ), .A2(_05744_ ), .ZN(_05849_ ) );
NOR3_X1 _13600_ ( .A1(_05849_ ), .A2(_05754_ ), .A3(_05814_ ), .ZN(_05850_ ) );
AND2_X1 _13601_ ( .A1(_05769_ ), .A2(_05786_ ), .ZN(_05851_ ) );
OR2_X1 _13602_ ( .A1(_05850_ ), .A2(_05851_ ), .ZN(_05852_ ) );
NOR3_X1 _13603_ ( .A1(_05779_ ), .A2(_05852_ ), .A3(_05792_ ), .ZN(_05853_ ) );
NAND3_X1 _13604_ ( .A1(_05825_ ), .A2(_05848_ ), .A3(_05853_ ), .ZN(_05854_ ) );
AND3_X1 _13605_ ( .A1(_05820_ ), .A2(_05776_ ), .A3(_05816_ ), .ZN(_05855_ ) );
AND2_X1 _13606_ ( .A1(_05855_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05856_ ) );
AND3_X1 _13607_ ( .A1(_05688_ ), .A2(\IF_ID_inst [12] ), .A3(_05689_ ), .ZN(_05857_ ) );
AND3_X1 _13608_ ( .A1(_05696_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_05858_ ) );
AND2_X2 _13609_ ( .A1(_05857_ ), .A2(_05858_ ), .ZN(_05859_ ) );
AND2_X1 _13610_ ( .A1(_05856_ ), .A2(_05859_ ), .ZN(_05860_ ) );
OAI21_X1 _13611_ ( .A(_05838_ ), .B1(_05817_ ), .B2(_05831_ ), .ZN(_05861_ ) );
INV_X1 _13612_ ( .A(_05861_ ), .ZN(_05862_ ) );
OAI22_X1 _13613_ ( .A1(_05860_ ), .A2(_05830_ ), .B1(_05862_ ), .B2(_05856_ ), .ZN(_05863_ ) );
AND2_X1 _13614_ ( .A1(_05818_ ), .A2(_05859_ ), .ZN(_05864_ ) );
INV_X1 _13615_ ( .A(_05864_ ), .ZN(_05865_ ) );
OAI21_X1 _13616_ ( .A(_05861_ ), .B1(_05833_ ), .B2(_05834_ ), .ZN(_05866_ ) );
AND2_X1 _13617_ ( .A1(_05866_ ), .A2(_05859_ ), .ZN(_05867_ ) );
INV_X1 _13618_ ( .A(_05867_ ), .ZN(_05868_ ) );
AND3_X1 _13619_ ( .A1(_05863_ ), .A2(_05865_ ), .A3(_05868_ ), .ZN(_05869_ ) );
INV_X1 _13620_ ( .A(_05869_ ), .ZN(_05870_ ) );
NOR2_X1 _13621_ ( .A1(_05854_ ), .A2(_05870_ ), .ZN(_05871_ ) );
XNOR2_X1 _13622_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_05872_ ) );
XNOR2_X1 _13623_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_05873_ ) );
XNOR2_X1 _13624_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_05874_ ) );
XNOR2_X1 _13625_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_05875_ ) );
AND4_X1 _13626_ ( .A1(_05872_ ), .A2(_05873_ ), .A3(_05874_ ), .A4(_05875_ ), .ZN(_05876_ ) );
XNOR2_X1 _13627_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_05877_ ) );
XNOR2_X1 _13628_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_05878_ ) );
XNOR2_X1 _13629_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_05879_ ) );
XNOR2_X1 _13630_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_05880_ ) );
AND4_X1 _13631_ ( .A1(_05877_ ), .A2(_05878_ ), .A3(_05879_ ), .A4(_05880_ ), .ZN(_05881_ ) );
XNOR2_X1 _13632_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_05882_ ) );
XNOR2_X1 _13633_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_05883_ ) );
XNOR2_X1 _13634_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_05884_ ) );
XNOR2_X1 _13635_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_05885_ ) );
AND4_X1 _13636_ ( .A1(_05882_ ), .A2(_05883_ ), .A3(_05884_ ), .A4(_05885_ ), .ZN(_05886_ ) );
INV_X1 _13637_ ( .A(\IF_ID_pc [2] ), .ZN(_05887_ ) );
AOI22_X1 _13638_ ( .A1(\IF_ID_pc [12] ), .A2(_05139_ ), .B1(_05887_ ), .B2(\myexu.pc_jump [2] ), .ZN(_05888_ ) );
XNOR2_X1 _13639_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_05889_ ) );
XNOR2_X1 _13640_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_05890_ ) );
AOI22_X1 _13641_ ( .A1(_02098_ ), .A2(\myexu.pc_jump [12] ), .B1(_05220_ ), .B2(\IF_ID_pc [10] ), .ZN(_05891_ ) );
AND4_X1 _13642_ ( .A1(_05888_ ), .A2(_05889_ ), .A3(_05890_ ), .A4(_05891_ ), .ZN(_05892_ ) );
AND4_X1 _13643_ ( .A1(_05876_ ), .A2(_05881_ ), .A3(_05886_ ), .A4(_05892_ ), .ZN(_05893_ ) );
XNOR2_X1 _13644_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_05894_ ) );
OAI221_X1 _13645_ ( .A(_05894_ ), .B1(\IF_ID_pc [27] ), .B2(_05473_ ), .C1(_02100_ ), .C2(\myexu.pc_jump [25] ), .ZN(_05895_ ) );
AOI22_X1 _13646_ ( .A1(\IF_ID_pc [17] ), .A2(_05002_ ), .B1(_02233_ ), .B2(\myexu.pc_jump [8] ), .ZN(_05896_ ) );
OAI221_X1 _13647_ ( .A(_05896_ ), .B1(_02091_ ), .B2(\myexu.pc_jump [21] ), .C1(\IF_ID_pc [17] ), .C2(_05002_ ), .ZN(_05897_ ) );
AOI22_X1 _13648_ ( .A1(_02269_ ), .A2(\myexu.pc_jump [28] ), .B1(_05561_ ), .B2(\IF_ID_pc [24] ), .ZN(_05898_ ) );
OAI221_X1 _13649_ ( .A(_05898_ ), .B1(\IF_ID_pc [24] ), .B2(_05561_ ), .C1(_02233_ ), .C2(\myexu.pc_jump [8] ), .ZN(_05899_ ) );
AOI22_X1 _13650_ ( .A1(\IF_ID_pc [26] ), .A2(_02391_ ), .B1(_02091_ ), .B2(\myexu.pc_jump [21] ), .ZN(_05900_ ) );
OAI221_X1 _13651_ ( .A(_05900_ ), .B1(_02280_ ), .B2(\myexu.pc_jump [27] ), .C1(\IF_ID_pc [26] ), .C2(_02391_ ), .ZN(_05901_ ) );
NOR4_X1 _13652_ ( .A1(_05895_ ), .A2(_05897_ ), .A3(_05899_ ), .A4(_05901_ ), .ZN(_05902_ ) );
XNOR2_X1 _13653_ ( .A(fanout_net_8 ), .B(\myexu.pc_jump [3] ), .ZN(_05903_ ) );
XNOR2_X1 _13654_ ( .A(fanout_net_12 ), .B(\myexu.pc_jump [4] ), .ZN(_05904_ ) );
AOI22_X1 _13655_ ( .A1(\IF_ID_pc [11] ), .A2(_05168_ ), .B1(_02208_ ), .B2(\myexu.pc_jump [10] ), .ZN(_05905_ ) );
INV_X1 _13656_ ( .A(\IF_ID_pc [11] ), .ZN(_05906_ ) );
AOI22_X1 _13657_ ( .A1(_02100_ ), .A2(\myexu.pc_jump [25] ), .B1(_05906_ ), .B2(\myexu.pc_jump [11] ), .ZN(_05907_ ) );
AND4_X1 _13658_ ( .A1(_05903_ ), .A2(_05904_ ), .A3(_05905_ ), .A4(_05907_ ), .ZN(_05908_ ) );
XNOR2_X1 _13659_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_05909_ ) );
XNOR2_X1 _13660_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_05910_ ) );
XNOR2_X1 _13661_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_05911_ ) );
AOI22_X1 _13662_ ( .A1(\IF_ID_pc [28] ), .A2(_02397_ ), .B1(_05425_ ), .B2(\IF_ID_pc [2] ), .ZN(_05912_ ) );
AND4_X1 _13663_ ( .A1(_05909_ ), .A2(_05910_ ), .A3(_05911_ ), .A4(_05912_ ), .ZN(_05913_ ) );
AND4_X1 _13664_ ( .A1(_05893_ ), .A2(_05902_ ), .A3(_05908_ ), .A4(_05913_ ), .ZN(_05914_ ) );
NOR2_X1 _13665_ ( .A1(_05914_ ), .A2(_02417_ ), .ZN(_05915_ ) );
INV_X1 _13666_ ( .A(\myifu.state [1] ), .ZN(_05916_ ) );
NOR2_X1 _13667_ ( .A1(_05916_ ), .A2(\myifu.to_reset ), .ZN(_05917_ ) );
INV_X1 _13668_ ( .A(_05917_ ), .ZN(_05918_ ) );
NOR2_X1 _13669_ ( .A1(_05915_ ), .A2(_05918_ ), .ZN(_05919_ ) );
NAND2_X1 _13670_ ( .A1(_05919_ ), .A2(IDU_ready_IFU ), .ZN(_05920_ ) );
NOR2_X1 _13671_ ( .A1(_05871_ ), .A2(_05920_ ), .ZN(_05921_ ) );
NOR2_X1 _13672_ ( .A1(_05921_ ), .A2(\ID_EX_rs1 [3] ), .ZN(_05922_ ) );
OR3_X1 _13673_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05794_ ), .ZN(_05923_ ) );
BUF_X2 _13674_ ( .A(_05921_ ), .Z(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
AOI211_X1 _13675_ ( .A(_05718_ ), .B(_05922_ ), .C1(_05923_ ), .C2(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00217_ ) );
INV_X1 _13676_ ( .A(\IF_ID_inst [16] ), .ZN(_05924_ ) );
NOR4_X1 _13677_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05924_ ), .A4(_05704_ ), .ZN(_00218_ ) );
NOR2_X1 _13678_ ( .A1(_05921_ ), .A2(\ID_EX_rs1 [2] ), .ZN(_05925_ ) );
OR3_X1 _13679_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05795_ ), .ZN(_05926_ ) );
AOI211_X1 _13680_ ( .A(_05718_ ), .B(_05925_ ), .C1(_05926_ ), .C2(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00219_ ) );
NOR4_X1 _13681_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05760_ ), .A4(_05704_ ), .ZN(_00220_ ) );
OAI21_X1 _13682_ ( .A(_05703_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [1] ), .ZN(_05927_ ) );
OR3_X1 _13683_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05924_ ), .ZN(_05928_ ) );
AOI21_X1 _13684_ ( .A(_05927_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(_05928_ ), .ZN(_00221_ ) );
NOR2_X1 _13685_ ( .A1(_05807_ ), .A2(_05789_ ), .ZN(_05929_ ) );
NOR2_X1 _13686_ ( .A1(_05824_ ), .A2(_05840_ ), .ZN(_05930_ ) );
AND2_X1 _13687_ ( .A1(_05929_ ), .A2(_05930_ ), .ZN(_05931_ ) );
NOR2_X1 _13688_ ( .A1(_05783_ ), .A2(_05851_ ), .ZN(_05932_ ) );
INV_X1 _13689_ ( .A(_05932_ ), .ZN(_05933_ ) );
NOR2_X1 _13690_ ( .A1(_05827_ ), .A2(_05933_ ), .ZN(_05934_ ) );
AND3_X2 _13691_ ( .A1(_05931_ ), .A2(_05846_ ), .A3(_05934_ ), .ZN(_05935_ ) );
AND3_X1 _13692_ ( .A1(_05762_ ), .A2(_05692_ ), .A3(_05729_ ), .ZN(_05936_ ) );
NOR2_X1 _13693_ ( .A1(_05738_ ), .A2(_05739_ ), .ZN(_05937_ ) );
AND2_X1 _13694_ ( .A1(_05936_ ), .A2(_05937_ ), .ZN(_05938_ ) );
AND4_X1 _13695_ ( .A1(_05707_ ), .A2(_05734_ ), .A3(\IF_ID_inst [20] ), .A4(_05735_ ), .ZN(_05939_ ) );
NAND2_X1 _13696_ ( .A1(_05938_ ), .A2(_05939_ ), .ZN(_05940_ ) );
NAND2_X1 _13697_ ( .A1(_05940_ ), .A2(_05700_ ), .ZN(_05941_ ) );
NOR2_X1 _13698_ ( .A1(_05791_ ), .A2(_05763_ ), .ZN(_05942_ ) );
OR2_X1 _13699_ ( .A1(_05942_ ), .A2(_05725_ ), .ZN(_05943_ ) );
AND2_X1 _13700_ ( .A1(_05802_ ), .A2(_05808_ ), .ZN(_05944_ ) );
INV_X1 _13701_ ( .A(_05944_ ), .ZN(_05945_ ) );
NOR3_X1 _13702_ ( .A1(_05941_ ), .A2(_05943_ ), .A3(_05945_ ), .ZN(_05946_ ) );
AND4_X1 _13703_ ( .A1(\IF_ID_inst [24] ), .A2(_05935_ ), .A3(_05759_ ), .A4(_05946_ ), .ZN(_00222_ ) );
NOR2_X1 _13704_ ( .A1(_05921_ ), .A2(\ID_EX_rs1 [0] ), .ZN(_05947_ ) );
OR3_X1 _13705_ ( .A1(_05779_ ), .A2(_05792_ ), .A3(_05760_ ), .ZN(_05948_ ) );
AOI211_X1 _13706_ ( .A(_05718_ ), .B(_05947_ ), .C1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .C2(_05948_ ), .ZN(_00223_ ) );
AND4_X1 _13707_ ( .A1(\IF_ID_inst [23] ), .A2(_05935_ ), .A3(_05703_ ), .A4(_05946_ ), .ZN(_00224_ ) );
AND4_X1 _13708_ ( .A1(\IF_ID_inst [22] ), .A2(_05935_ ), .A3(_05703_ ), .A4(_05946_ ), .ZN(_00225_ ) );
AND2_X1 _13709_ ( .A1(_05935_ ), .A2(_05946_ ), .ZN(_05949_ ) );
AOI211_X1 _13710_ ( .A(_05920_ ), .B(_05871_ ), .C1(\IF_ID_inst [23] ), .C2(_05949_ ), .ZN(_05950_ ) );
INV_X1 _13711_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_05951_ ) );
AOI211_X1 _13712_ ( .A(_05718_ ), .B(_05950_ ), .C1(_03637_ ), .C2(_05951_ ), .ZN(_00226_ ) );
AND4_X1 _13713_ ( .A1(\IF_ID_inst [21] ), .A2(_05935_ ), .A3(_05703_ ), .A4(_05946_ ), .ZN(_00227_ ) );
NAND3_X1 _13714_ ( .A1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .A2(\IF_ID_inst [22] ), .A3(_05949_ ), .ZN(_05952_ ) );
OAI21_X1 _13715_ ( .A(\ID_EX_rs2 [2] ), .B1(_05871_ ), .B2(_05920_ ), .ZN(_05953_ ) );
AOI21_X1 _13716_ ( .A(_05708_ ), .B1(_05952_ ), .B2(_05953_ ), .ZN(_00228_ ) );
AND4_X1 _13717_ ( .A1(\IF_ID_inst [20] ), .A2(_05935_ ), .A3(_05703_ ), .A4(_05946_ ), .ZN(_00229_ ) );
NAND3_X1 _13718_ ( .A1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .A2(\IF_ID_inst [21] ), .A3(_05949_ ), .ZN(_05954_ ) );
OAI21_X1 _13719_ ( .A(\ID_EX_rs2 [1] ), .B1(_05871_ ), .B2(_05920_ ), .ZN(_05955_ ) );
AOI21_X1 _13720_ ( .A(_05708_ ), .B1(_05954_ ), .B2(_05955_ ), .ZN(_00230_ ) );
AND4_X1 _13721_ ( .A1(_02405_ ), .A2(_05722_ ), .A3(_05703_ ), .A4(_05724_ ), .ZN(_00231_ ) );
OAI21_X1 _13722_ ( .A(_05703_ ), .B1(_05921_ ), .B2(\ID_EX_rs2 [0] ), .ZN(_05956_ ) );
NAND3_X1 _13723_ ( .A1(_05935_ ), .A2(\IF_ID_inst [20] ), .A3(_05946_ ), .ZN(_05957_ ) );
AOI21_X1 _13724_ ( .A(_05956_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(_05957_ ), .ZN(_00232_ ) );
AND2_X1 _13725_ ( .A1(_03342_ ), .A2(_02406_ ), .ZN(_05958_ ) );
XNOR2_X1 _13726_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_05959_ ) );
XNOR2_X1 _13727_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_05960_ ) );
XNOR2_X1 _13728_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_05961_ ) );
NAND4_X1 _13729_ ( .A1(_05958_ ), .A2(_05959_ ), .A3(_05960_ ), .A4(_05961_ ), .ZN(_05962_ ) );
XNOR2_X1 _13730_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_05963_ ) );
XNOR2_X1 _13731_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_05964_ ) );
NAND2_X1 _13732_ ( .A1(_05963_ ), .A2(_05964_ ), .ZN(_05965_ ) );
NOR2_X1 _13733_ ( .A1(_05962_ ), .A2(_05965_ ), .ZN(_05966_ ) );
INV_X1 _13734_ ( .A(_05827_ ), .ZN(_05967_ ) );
NAND2_X1 _13735_ ( .A1(_05967_ ), .A2(_05842_ ), .ZN(_05968_ ) );
OR4_X1 _13736_ ( .A1(_05810_ ), .A2(_05968_ ), .A3(_05844_ ), .A4(_05851_ ), .ZN(_05969_ ) );
NOR2_X2 _13737_ ( .A1(_05969_ ), .A2(_05806_ ), .ZN(_05970_ ) );
AOI21_X1 _13738_ ( .A(_05966_ ), .B1(_05970_ ), .B2(_05700_ ), .ZN(_05971_ ) );
INV_X1 _13739_ ( .A(_05942_ ), .ZN(_05972_ ) );
XNOR2_X1 _13740_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_05973_ ) );
XNOR2_X1 _13741_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_05974_ ) );
XNOR2_X1 _13742_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_05975_ ) );
AND4_X1 _13743_ ( .A1(_05958_ ), .A2(_05973_ ), .A3(_05974_ ), .A4(_05975_ ), .ZN(_05976_ ) );
XNOR2_X1 _13744_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_05977_ ) );
XNOR2_X1 _13745_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_05978_ ) );
NAND3_X1 _13746_ ( .A1(_05976_ ), .A2(_05977_ ), .A3(_05978_ ), .ZN(_05979_ ) );
OAI21_X1 _13747_ ( .A(_05979_ ), .B1(_05965_ ), .B2(_05962_ ), .ZN(_05980_ ) );
AND4_X1 _13748_ ( .A1(_05972_ ), .A2(_05741_ ), .A3(_05790_ ), .A4(_05980_ ), .ZN(_05981_ ) );
NOR4_X1 _13749_ ( .A1(_05969_ ), .A2(_05709_ ), .A3(_05806_ ), .A4(_05981_ ), .ZN(_05982_ ) );
INV_X1 _13750_ ( .A(IDU_ready_IFU ), .ZN(_05983_ ) );
NOR4_X1 _13751_ ( .A1(_05971_ ), .A2(_05982_ ), .A3(_05983_ ), .A4(_05704_ ), .ZN(_00233_ ) );
NOR2_X1 _13752_ ( .A1(_05849_ ), .A2(_05814_ ), .ZN(_05984_ ) );
NOR2_X1 _13753_ ( .A1(_05774_ ), .A2(_05984_ ), .ZN(_05985_ ) );
AND3_X1 _13754_ ( .A1(_05693_ ), .A2(_05747_ ), .A3(_05744_ ), .ZN(_05986_ ) );
AOI21_X1 _13755_ ( .A(_05986_ ), .B1(_05692_ ), .B2(_05769_ ), .ZN(_05987_ ) );
NAND2_X2 _13756_ ( .A1(_05985_ ), .A2(_05987_ ), .ZN(_05988_ ) );
NOR3_X1 _13757_ ( .A1(_05943_ ), .A2(_05988_ ), .A3(_05933_ ), .ZN(_05989_ ) );
NAND4_X1 _13758_ ( .A1(_05692_ ), .A2(_05761_ ), .A3(_05694_ ), .A4(_05747_ ), .ZN(_05990_ ) );
NOR4_X1 _13759_ ( .A1(_05990_ ), .A2(\IF_ID_inst [20] ), .A3(\IF_ID_inst [8] ), .A4(_05728_ ), .ZN(_05991_ ) );
AND3_X1 _13760_ ( .A1(_05734_ ), .A2(_05707_ ), .A3(_05735_ ), .ZN(_05992_ ) );
AND2_X1 _13761_ ( .A1(_05992_ ), .A2(_05937_ ), .ZN(_05993_ ) );
NAND2_X1 _13762_ ( .A1(_05991_ ), .A2(_05993_ ), .ZN(_05994_ ) );
AND2_X1 _13763_ ( .A1(_05994_ ), .A2(_05700_ ), .ZN(_05995_ ) );
AOI21_X1 _13764_ ( .A(_05708_ ), .B1(_05989_ ), .B2(_05995_ ), .ZN(_00234_ ) );
BUF_X4 _13765_ ( .A(_05797_ ), .Z(_05996_ ) );
AND2_X1 _13766_ ( .A1(_05843_ ), .A2(_05692_ ), .ZN(_05997_ ) );
AND2_X1 _13767_ ( .A1(_05997_ ), .A2(_05747_ ), .ZN(_05998_ ) );
AND3_X1 _13768_ ( .A1(_05997_ ), .A2(_05754_ ), .A3(\IF_ID_inst [14] ), .ZN(_05999_ ) );
NOR4_X1 _13769_ ( .A1(_05996_ ), .A2(_05968_ ), .A3(_05998_ ), .A4(_05999_ ), .ZN(_06000_ ) );
AOI21_X1 _13770_ ( .A(_05708_ ), .B1(_06000_ ), .B2(_05995_ ), .ZN(_00235_ ) );
NAND2_X1 _13771_ ( .A1(_05863_ ), .A2(_05868_ ), .ZN(_06001_ ) );
AND3_X1 _13772_ ( .A1(_05938_ ), .A2(_05710_ ), .A3(_05992_ ), .ZN(_06002_ ) );
OR2_X1 _13773_ ( .A1(_05836_ ), .A2(_05864_ ), .ZN(_06003_ ) );
NOR4_X1 _13774_ ( .A1(_06001_ ), .A2(_05945_ ), .A3(_06002_ ), .A4(_06003_ ), .ZN(_06004_ ) );
AOI21_X1 _13775_ ( .A(_05708_ ), .B1(_06004_ ), .B2(_05935_ ), .ZN(_00236_ ) );
AOI221_X4 _13776_ ( .A(_05725_ ), .B1(_05803_ ), .B2(\IF_ID_inst [13] ), .C1(_05800_ ), .C2(_05801_ ), .ZN(_06005_ ) );
AOI21_X1 _13777_ ( .A(_05708_ ), .B1(_05931_ ), .B2(_06005_ ), .ZN(_00237_ ) );
AOI221_X4 _13778_ ( .A(_05756_ ), .B1(_05830_ ), .B2(_05835_ ), .C1(_05764_ ), .C2(_05768_ ), .ZN(_06006_ ) );
AOI21_X1 _13779_ ( .A(_05705_ ), .B1(_06006_ ), .B2(_05929_ ), .ZN(_00238_ ) );
AOI211_X1 _13780_ ( .A(_05984_ ), .B(_05809_ ), .C1(\IF_ID_inst [13] ), .C2(_05695_ ), .ZN(_06007_ ) );
INV_X1 _13781_ ( .A(_05789_ ), .ZN(_06008_ ) );
AOI22_X1 _13782_ ( .A1(_05826_ ), .A2(_05755_ ), .B1(_05818_ ), .B2(_05859_ ), .ZN(_06009_ ) );
AND4_X1 _13783_ ( .A1(_05757_ ), .A2(_06007_ ), .A3(_06008_ ), .A4(_06009_ ), .ZN(_06010_ ) );
NOR3_X1 _13784_ ( .A1(_05867_ ), .A2(_05824_ ), .A3(_05840_ ), .ZN(_06011_ ) );
AOI21_X1 _13785_ ( .A(_05705_ ), .B1(_06010_ ), .B2(_06011_ ), .ZN(_00239_ ) );
NAND2_X1 _13786_ ( .A1(_05800_ ), .A2(\IF_ID_inst [14] ), .ZN(_06012_ ) );
AND3_X1 _13787_ ( .A1(_05751_ ), .A2(_05747_ ), .A3(_05744_ ), .ZN(_06013_ ) );
AOI221_X4 _13788_ ( .A(_06013_ ), .B1(_05747_ ), .B2(_05997_ ), .C1(_05786_ ), .C2(_05858_ ), .ZN(_06014_ ) );
NOR2_X1 _13789_ ( .A1(_05756_ ), .A2(_05999_ ), .ZN(_06015_ ) );
AOI21_X1 _13790_ ( .A(_05699_ ), .B1(\IF_ID_inst [14] ), .B2(_05773_ ), .ZN(_06016_ ) );
AND4_X1 _13791_ ( .A1(_06012_ ), .A2(_06014_ ), .A3(_06015_ ), .A4(_06016_ ), .ZN(_06017_ ) );
AND2_X1 _13792_ ( .A1(_05838_ ), .A2(_05817_ ), .ZN(_06018_ ) );
OAI21_X1 _13793_ ( .A(_05830_ ), .B1(_05856_ ), .B2(_06018_ ), .ZN(_06019_ ) );
OAI22_X1 _13794_ ( .A1(_05818_ ), .A2(_05822_ ), .B1(_05803_ ), .B2(_05859_ ), .ZN(_06020_ ) );
AND2_X1 _13795_ ( .A1(_06019_ ), .A2(_06020_ ), .ZN(_06021_ ) );
AOI21_X1 _13796_ ( .A(_05705_ ), .B1(_06017_ ), .B2(_06021_ ), .ZN(_00240_ ) );
NAND4_X1 _13797_ ( .A1(_05940_ ), .A2(_05753_ ), .A3(_05804_ ), .A4(_05841_ ), .ZN(_06022_ ) );
AOI21_X1 _13798_ ( .A(_05699_ ), .B1(_05826_ ), .B2(_05754_ ), .ZN(_06023_ ) );
NAND3_X1 _13799_ ( .A1(_05693_ ), .A2(_05754_ ), .A3(_05694_ ), .ZN(_06024_ ) );
AOI21_X1 _13800_ ( .A(_05814_ ), .B1(_06023_ ), .B2(_06024_ ), .ZN(_06025_ ) );
NAND3_X1 _13801_ ( .A1(_05693_ ), .A2(_05747_ ), .A3(_05744_ ), .ZN(_06026_ ) );
NAND4_X1 _13802_ ( .A1(_05798_ ), .A2(_05694_ ), .A3(_05817_ ), .A4(_05838_ ), .ZN(_06027_ ) );
NAND3_X1 _13803_ ( .A1(_06015_ ), .A2(_06026_ ), .A3(_06027_ ), .ZN(_06028_ ) );
NOR4_X1 _13804_ ( .A1(_06022_ ), .A2(_06025_ ), .A3(_06028_ ), .A4(_05852_ ), .ZN(_06029_ ) );
OAI21_X1 _13805_ ( .A(_05859_ ), .B1(_05839_ ), .B2(_05818_ ), .ZN(_06030_ ) );
AND4_X1 _13806_ ( .A1(_05751_ ), .A2(_05813_ ), .A3(_05799_ ), .A4(_05817_ ), .ZN(_06031_ ) );
AOI21_X1 _13807_ ( .A(_06031_ ), .B1(_05856_ ), .B2(_05859_ ), .ZN(_06032_ ) );
OAI21_X1 _13808_ ( .A(_05776_ ), .B1(_05695_ ), .B2(_05773_ ), .ZN(_06033_ ) );
NOR2_X1 _13809_ ( .A1(_05833_ ), .A2(_05834_ ), .ZN(_06034_ ) );
AOI22_X1 _13810_ ( .A1(_05815_ ), .A2(_05800_ ), .B1(_05830_ ), .B2(_06034_ ), .ZN(_06035_ ) );
AND4_X1 _13811_ ( .A1(_06030_ ), .A2(_06032_ ), .A3(_06033_ ), .A4(_06035_ ), .ZN(_06036_ ) );
AOI21_X1 _13812_ ( .A(_05705_ ), .B1(_06029_ ), .B2(_06036_ ), .ZN(_00241_ ) );
INV_X1 _13813_ ( .A(_05914_ ), .ZN(_06037_ ) );
INV_X1 _13814_ ( .A(\myifu.to_reset ), .ZN(_06038_ ) );
BUF_X4 _13815_ ( .A(_06038_ ), .Z(_06039_ ) );
BUF_X4 _13816_ ( .A(_06039_ ), .Z(_06040_ ) );
NAND4_X1 _13817_ ( .A1(_06037_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_06040_ ), .ZN(_06041_ ) );
NAND2_X1 _13818_ ( .A1(\mtvec [0] ), .A2(\myifu.to_reset ), .ZN(_06042_ ) );
AOI21_X1 _13819_ ( .A(fanout_net_3 ), .B1(_06041_ ), .B2(_06042_ ), .ZN(_00245_ ) );
NOR2_X1 _13820_ ( .A1(_06040_ ), .A2(\mtvec [30] ), .ZN(_06043_ ) );
NOR4_X4 _13821_ ( .A1(_05702_ ), .A2(_05742_ ), .A3(\IF_ID_inst [4] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_06044_ ) );
AND2_X1 _13822_ ( .A1(_06044_ ), .A2(_05691_ ), .ZN(_06045_ ) );
BUF_X4 _13823_ ( .A(_06045_ ), .Z(_06046_ ) );
AND2_X1 _13824_ ( .A1(_06046_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_06047_ ) );
CLKBUF_X2 _13825_ ( .A(_05781_ ), .Z(_06048_ ) );
OAI211_X1 _13826_ ( .A(_06048_ ), .B(\IF_ID_inst [31] ), .C1(_05691_ ), .C2(_05724_ ), .ZN(_06049_ ) );
NOR2_X2 _13827_ ( .A1(_06047_ ), .A2(_06049_ ), .ZN(_06050_ ) );
BUF_X4 _13828_ ( .A(_06050_ ), .Z(_06051_ ) );
BUF_X4 _13829_ ( .A(_06051_ ), .Z(_06052_ ) );
XNOR2_X1 _13830_ ( .A(_06052_ ), .B(_02064_ ), .ZN(_06053_ ) );
INV_X1 _13831_ ( .A(_06053_ ), .ZN(_06054_ ) );
XNOR2_X1 _13832_ ( .A(_06051_ ), .B(_02100_ ), .ZN(_06055_ ) );
INV_X1 _13833_ ( .A(_06055_ ), .ZN(_06056_ ) );
INV_X1 _13834_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_06057_ ) );
AND3_X1 _13835_ ( .A1(_06044_ ), .A2(_06057_ ), .A3(_05691_ ), .ZN(_06058_ ) );
AOI21_X1 _13836_ ( .A(_06058_ ), .B1(_05783_ ), .B2(\IF_ID_inst [29] ), .ZN(_06059_ ) );
XNOR2_X1 _13837_ ( .A(_06059_ ), .B(\IF_ID_pc [9] ), .ZN(_06060_ ) );
INV_X1 _13838_ ( .A(_06060_ ), .ZN(_06061_ ) );
AND2_X1 _13839_ ( .A1(_05783_ ), .A2(\IF_ID_inst [26] ), .ZN(_06062_ ) );
INV_X1 _13840_ ( .A(_06062_ ), .ZN(_06063_ ) );
INV_X1 _13841_ ( .A(_06045_ ), .ZN(_06064_ ) );
OAI21_X1 _13842_ ( .A(_06063_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_06064_ ), .ZN(_06065_ ) );
NAND2_X1 _13843_ ( .A1(_06065_ ), .A2(\IF_ID_pc [6] ), .ZN(_06066_ ) );
AND2_X1 _13844_ ( .A1(_05782_ ), .A2(\IF_ID_inst [25] ), .ZN(_06067_ ) );
INV_X1 _13845_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_06068_ ) );
AND3_X1 _13846_ ( .A1(_06044_ ), .A2(_06068_ ), .A3(_05691_ ), .ZN(_06069_ ) );
NOR2_X1 _13847_ ( .A1(_06067_ ), .A2(_06069_ ), .ZN(_06070_ ) );
OR2_X1 _13848_ ( .A1(_06064_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_06071_ ) );
NAND3_X1 _13849_ ( .A1(_06048_ ), .A2(\IF_ID_inst [24] ), .A3(_05723_ ), .ZN(_06072_ ) );
NAND2_X1 _13850_ ( .A1(_06071_ ), .A2(_06072_ ), .ZN(_06073_ ) );
NAND2_X1 _13851_ ( .A1(_06073_ ), .A2(fanout_net_12 ), .ZN(_06074_ ) );
AND3_X1 _13852_ ( .A1(_05781_ ), .A2(\IF_ID_inst [23] ), .A3(_05723_ ), .ZN(_06075_ ) );
INV_X1 _13853_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_06076_ ) );
AND3_X1 _13854_ ( .A1(_06044_ ), .A2(_06076_ ), .A3(_05691_ ), .ZN(_06077_ ) );
OR2_X1 _13855_ ( .A1(_06075_ ), .A2(_06077_ ), .ZN(_06078_ ) );
INV_X1 _13856_ ( .A(_06078_ ), .ZN(_06079_ ) );
OR2_X1 _13857_ ( .A1(_06079_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06080_ ) );
NAND3_X1 _13858_ ( .A1(_05781_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .A3(_05723_ ), .ZN(_06081_ ) );
NAND3_X1 _13859_ ( .A1(_06044_ ), .A2(_05690_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_06082_ ) );
AND3_X1 _13860_ ( .A1(_06081_ ), .A2(\IF_ID_pc [2] ), .A3(_06082_ ), .ZN(_06083_ ) );
AOI21_X1 _13861_ ( .A(\IF_ID_pc [2] ), .B1(_06081_ ), .B2(_06082_ ), .ZN(_06084_ ) );
NOR2_X1 _13862_ ( .A1(_06083_ ), .A2(_06084_ ), .ZN(_06085_ ) );
NAND3_X1 _13863_ ( .A1(_05781_ ), .A2(\IF_ID_inst [21] ), .A3(_05723_ ), .ZN(_06086_ ) );
INV_X1 _13864_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_06087_ ) );
NAND3_X1 _13865_ ( .A1(_06044_ ), .A2(_05691_ ), .A3(_06087_ ), .ZN(_06088_ ) );
NAND2_X1 _13866_ ( .A1(_06086_ ), .A2(_06088_ ), .ZN(_06089_ ) );
AND2_X1 _13867_ ( .A1(_06089_ ), .A2(\IF_ID_pc [1] ), .ZN(_06090_ ) );
AND2_X1 _13868_ ( .A1(_06085_ ), .A2(_06090_ ), .ZN(_06091_ ) );
NOR2_X1 _13869_ ( .A1(_06091_ ), .A2(_06083_ ), .ZN(_06092_ ) );
XNOR2_X1 _13870_ ( .A(_06078_ ), .B(fanout_net_8 ), .ZN(_06093_ ) );
OAI211_X1 _13871_ ( .A(_06074_ ), .B(_06080_ ), .C1(_06092_ ), .C2(_06093_ ), .ZN(_06094_ ) );
INV_X1 _13872_ ( .A(fanout_net_12 ), .ZN(_06095_ ) );
NAND3_X1 _13873_ ( .A1(_06071_ ), .A2(_06095_ ), .A3(_06072_ ), .ZN(_06096_ ) );
NAND2_X1 _13874_ ( .A1(_06094_ ), .A2(_06096_ ), .ZN(_06097_ ) );
INV_X1 _13875_ ( .A(\IF_ID_pc [5] ), .ZN(_06098_ ) );
XNOR2_X1 _13876_ ( .A(_06070_ ), .B(_06098_ ), .ZN(_06099_ ) );
OAI221_X1 _13877_ ( .A(_06066_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_06070_ ), .C1(_06097_ ), .C2(_06099_ ), .ZN(_06100_ ) );
AND2_X1 _13878_ ( .A1(_05783_ ), .A2(\IF_ID_inst [27] ), .ZN(_06101_ ) );
INV_X1 _13879_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_06102_ ) );
AOI21_X1 _13880_ ( .A(_06101_ ), .B1(_06102_ ), .B2(_06046_ ), .ZN(_06103_ ) );
XNOR2_X1 _13881_ ( .A(_06103_ ), .B(\IF_ID_pc [7] ), .ZN(_06104_ ) );
OR2_X1 _13882_ ( .A1(_06065_ ), .A2(\IF_ID_pc [6] ), .ZN(_06105_ ) );
AND3_X1 _13883_ ( .A1(_06100_ ), .A2(_06104_ ), .A3(_06105_ ), .ZN(_06106_ ) );
NOR2_X1 _13884_ ( .A1(_06103_ ), .A2(_02076_ ), .ZN(_06107_ ) );
AND2_X1 _13885_ ( .A1(_05783_ ), .A2(\IF_ID_inst [28] ), .ZN(_06108_ ) );
INV_X1 _13886_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_06109_ ) );
AOI21_X1 _13887_ ( .A(_06108_ ), .B1(_06109_ ), .B2(_06046_ ), .ZN(_06110_ ) );
INV_X1 _13888_ ( .A(_06110_ ), .ZN(_06111_ ) );
OAI22_X1 _13889_ ( .A1(_06106_ ), .A2(_06107_ ), .B1(\IF_ID_pc [8] ), .B2(_06111_ ), .ZN(_06112_ ) );
OR2_X1 _13890_ ( .A1(_06110_ ), .A2(_02233_ ), .ZN(_06113_ ) );
AOI21_X2 _13891_ ( .A(_06061_ ), .B1(_06112_ ), .B2(_06113_ ), .ZN(_06114_ ) );
AND2_X1 _13892_ ( .A1(_05783_ ), .A2(\IF_ID_inst [30] ), .ZN(_06115_ ) );
INV_X1 _13893_ ( .A(_06115_ ), .ZN(_06116_ ) );
OAI21_X1 _13894_ ( .A(_06116_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_06064_ ), .ZN(_06117_ ) );
AND2_X1 _13895_ ( .A1(_06117_ ), .A2(\IF_ID_pc [10] ), .ZN(_06118_ ) );
INV_X1 _13896_ ( .A(\IF_ID_pc [9] ), .ZN(_06119_ ) );
NOR2_X1 _13897_ ( .A1(_06059_ ), .A2(_06119_ ), .ZN(_06120_ ) );
OR3_X1 _13898_ ( .A1(_06114_ ), .A2(_06118_ ), .A3(_06120_ ), .ZN(_06121_ ) );
AND2_X1 _13899_ ( .A1(_05783_ ), .A2(\IF_ID_inst [20] ), .ZN(_06122_ ) );
INV_X1 _13900_ ( .A(_06122_ ), .ZN(_06123_ ) );
OAI21_X1 _13901_ ( .A(_06123_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_06064_ ), .ZN(_06124_ ) );
XNOR2_X1 _13902_ ( .A(_06124_ ), .B(_05906_ ), .ZN(_06125_ ) );
NOR2_X1 _13903_ ( .A1(_06117_ ), .A2(\IF_ID_pc [10] ), .ZN(_06126_ ) );
INV_X1 _13904_ ( .A(_06126_ ), .ZN(_06127_ ) );
AND3_X4 _13905_ ( .A1(_06121_ ), .A2(_06125_ ), .A3(_06127_ ), .ZN(_06128_ ) );
AND3_X1 _13906_ ( .A1(_06048_ ), .A2(\IF_ID_inst [12] ), .A3(_05724_ ), .ZN(_06129_ ) );
INV_X1 _13907_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_06130_ ) );
MUX2_X1 _13908_ ( .A(_06129_ ), .B(_06130_ ), .S(_06046_ ), .Z(_06131_ ) );
AND2_X1 _13909_ ( .A1(_06131_ ), .A2(\IF_ID_pc [12] ), .ZN(_06132_ ) );
AND2_X1 _13910_ ( .A1(_06124_ ), .A2(\IF_ID_pc [11] ), .ZN(_06133_ ) );
NOR3_X1 _13911_ ( .A1(_06128_ ), .A2(_06132_ ), .A3(_06133_ ), .ZN(_06134_ ) );
NOR2_X1 _13912_ ( .A1(_06131_ ), .A2(\IF_ID_pc [12] ), .ZN(_06135_ ) );
AND3_X1 _13913_ ( .A1(_06048_ ), .A2(\IF_ID_inst [14] ), .A3(_05723_ ), .ZN(_06136_ ) );
MUX2_X1 _13914_ ( .A(_06136_ ), .B(_06130_ ), .S(_06046_ ), .Z(_06137_ ) );
XNOR2_X1 _13915_ ( .A(_06137_ ), .B(_02081_ ), .ZN(_06138_ ) );
AND3_X1 _13916_ ( .A1(_06048_ ), .A2(\IF_ID_inst [13] ), .A3(_05724_ ), .ZN(_06139_ ) );
MUX2_X1 _13917_ ( .A(_06139_ ), .B(_06130_ ), .S(_06046_ ), .Z(_06140_ ) );
XNOR2_X1 _13918_ ( .A(_06140_ ), .B(_02157_ ), .ZN(_06141_ ) );
NAND2_X1 _13919_ ( .A1(_06138_ ), .A2(_06141_ ), .ZN(_06142_ ) );
NOR3_X2 _13920_ ( .A1(_06134_ ), .A2(_06135_ ), .A3(_06142_ ), .ZN(_06143_ ) );
INV_X1 _13921_ ( .A(_05783_ ), .ZN(_06144_ ) );
OAI21_X1 _13922_ ( .A(_06064_ ), .B1(_06144_ ), .B2(_05924_ ), .ZN(_06145_ ) );
INV_X1 _13923_ ( .A(_06047_ ), .ZN(_06146_ ) );
AND3_X1 _13924_ ( .A1(_06145_ ), .A2(\IF_ID_pc [16] ), .A3(_06146_ ), .ZN(_06147_ ) );
AOI21_X1 _13925_ ( .A(\IF_ID_pc [16] ), .B1(_06145_ ), .B2(_06146_ ), .ZN(_06148_ ) );
NAND3_X1 _13926_ ( .A1(_06048_ ), .A2(\IF_ID_inst [15] ), .A3(_05724_ ), .ZN(_06149_ ) );
MUX2_X1 _13927_ ( .A(_06149_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .S(_06046_ ), .Z(_06150_ ) );
NOR3_X1 _13928_ ( .A1(_06148_ ), .A2(_02150_ ), .A3(_06150_ ), .ZN(_06151_ ) );
AND2_X1 _13929_ ( .A1(_06137_ ), .A2(\IF_ID_pc [14] ), .ZN(_06152_ ) );
AND2_X1 _13930_ ( .A1(_06140_ ), .A2(\IF_ID_pc [13] ), .ZN(_06153_ ) );
AOI21_X1 _13931_ ( .A(_06152_ ), .B1(_06138_ ), .B2(_06153_ ), .ZN(_06154_ ) );
INV_X1 _13932_ ( .A(_06154_ ), .ZN(_06155_ ) );
NOR4_X1 _13933_ ( .A1(_06143_ ), .A2(_06147_ ), .A3(_06151_ ), .A4(_06155_ ), .ZN(_06156_ ) );
NOR2_X1 _13934_ ( .A1(_06147_ ), .A2(_06148_ ), .ZN(_06157_ ) );
XNOR2_X1 _13935_ ( .A(_06150_ ), .B(\IF_ID_pc [15] ), .ZN(_06158_ ) );
AOI211_X1 _13936_ ( .A(_06147_ ), .B(_06151_ ), .C1(_06157_ ), .C2(_06158_ ), .ZN(_06159_ ) );
NOR2_X1 _13937_ ( .A1(_06156_ ), .A2(_06159_ ), .ZN(_06160_ ) );
XNOR2_X1 _13938_ ( .A(_06050_ ), .B(_02166_ ), .ZN(_06161_ ) );
XNOR2_X1 _13939_ ( .A(_06050_ ), .B(_02091_ ), .ZN(_06162_ ) );
AND2_X1 _13940_ ( .A1(_06161_ ), .A2(_06162_ ), .ZN(_06163_ ) );
XNOR2_X1 _13941_ ( .A(_06050_ ), .B(_02276_ ), .ZN(_06164_ ) );
XNOR2_X1 _13942_ ( .A(_06050_ ), .B(_02222_ ), .ZN(_06165_ ) );
AND2_X1 _13943_ ( .A1(_06164_ ), .A2(_06165_ ), .ZN(_06166_ ) );
AND2_X1 _13944_ ( .A1(_06163_ ), .A2(_06166_ ), .ZN(_06167_ ) );
AND3_X1 _13945_ ( .A1(_06048_ ), .A2(\IF_ID_inst [19] ), .A3(_05724_ ), .ZN(_06168_ ) );
MUX2_X1 _13946_ ( .A(_06168_ ), .B(_06130_ ), .S(_06046_ ), .Z(_06169_ ) );
XNOR2_X1 _13947_ ( .A(_06169_ ), .B(_02308_ ), .ZN(_06170_ ) );
XNOR2_X1 _13948_ ( .A(_06050_ ), .B(_02069_ ), .ZN(_06171_ ) );
AND2_X1 _13949_ ( .A1(_06170_ ), .A2(_06171_ ), .ZN(_06172_ ) );
AND3_X1 _13950_ ( .A1(_06048_ ), .A2(\IF_ID_inst [18] ), .A3(_05724_ ), .ZN(_06173_ ) );
MUX2_X1 _13951_ ( .A(_06173_ ), .B(_06130_ ), .S(_06046_ ), .Z(_06174_ ) );
XNOR2_X1 _13952_ ( .A(_06174_ ), .B(_02083_ ), .ZN(_06175_ ) );
AND3_X1 _13953_ ( .A1(_06048_ ), .A2(\IF_ID_inst [17] ), .A3(_05724_ ), .ZN(_06176_ ) );
MUX2_X1 _13954_ ( .A(_06176_ ), .B(_06130_ ), .S(_06046_ ), .Z(_06177_ ) );
XNOR2_X1 _13955_ ( .A(_06177_ ), .B(_02142_ ), .ZN(_06178_ ) );
AND3_X1 _13956_ ( .A1(_06172_ ), .A2(_06175_ ), .A3(_06178_ ), .ZN(_06179_ ) );
AND3_X1 _13957_ ( .A1(_06160_ ), .A2(_06167_ ), .A3(_06179_ ), .ZN(_06180_ ) );
INV_X1 _13958_ ( .A(_06180_ ), .ZN(_06181_ ) );
NOR2_X1 _13959_ ( .A1(_06174_ ), .A2(\IF_ID_pc [18] ), .ZN(_06182_ ) );
INV_X1 _13960_ ( .A(_06182_ ), .ZN(_06183_ ) );
AND2_X1 _13961_ ( .A1(_06174_ ), .A2(\IF_ID_pc [18] ), .ZN(_06184_ ) );
AND2_X1 _13962_ ( .A1(_06177_ ), .A2(\IF_ID_pc [17] ), .ZN(_06185_ ) );
OR2_X1 _13963_ ( .A1(_06184_ ), .A2(_06185_ ), .ZN(_06186_ ) );
AND4_X1 _13964_ ( .A1(_06183_ ), .A2(_06186_ ), .A3(_06171_ ), .A4(_06170_ ), .ZN(_06187_ ) );
AND2_X1 _13965_ ( .A1(_06050_ ), .A2(\IF_ID_pc [20] ), .ZN(_06188_ ) );
AND2_X1 _13966_ ( .A1(_06169_ ), .A2(\IF_ID_pc [19] ), .ZN(_06189_ ) );
NOR2_X1 _13967_ ( .A1(_06051_ ), .A2(\IF_ID_pc [20] ), .ZN(_06190_ ) );
INV_X1 _13968_ ( .A(_06190_ ), .ZN(_06191_ ) );
AOI21_X1 _13969_ ( .A(_06188_ ), .B1(_06189_ ), .B2(_06191_ ), .ZN(_06192_ ) );
INV_X1 _13970_ ( .A(_06192_ ), .ZN(_06193_ ) );
OAI21_X1 _13971_ ( .A(_06167_ ), .B1(_06187_ ), .B2(_06193_ ), .ZN(_06194_ ) );
AND2_X1 _13972_ ( .A1(_06051_ ), .A2(\IF_ID_pc [22] ), .ZN(_06195_ ) );
AND2_X1 _13973_ ( .A1(_06051_ ), .A2(\IF_ID_pc [21] ), .ZN(_06196_ ) );
OAI21_X1 _13974_ ( .A(_06166_ ), .B1(_06195_ ), .B2(_06196_ ), .ZN(_06197_ ) );
NAND2_X1 _13975_ ( .A1(_06051_ ), .A2(\IF_ID_pc [24] ), .ZN(_06198_ ) );
NAND2_X1 _13976_ ( .A1(_06051_ ), .A2(\IF_ID_pc [23] ), .ZN(_06199_ ) );
AND3_X1 _13977_ ( .A1(_06197_ ), .A2(_06198_ ), .A3(_06199_ ), .ZN(_06200_ ) );
AND2_X1 _13978_ ( .A1(_06194_ ), .A2(_06200_ ), .ZN(_06201_ ) );
AOI21_X1 _13979_ ( .A(_06056_ ), .B1(_06181_ ), .B2(_06201_ ), .ZN(_06202_ ) );
XNOR2_X1 _13980_ ( .A(_06051_ ), .B(_02269_ ), .ZN(_06203_ ) );
XNOR2_X1 _13981_ ( .A(_06051_ ), .B(_02280_ ), .ZN(_06204_ ) );
XNOR2_X1 _13982_ ( .A(_06052_ ), .B(_02200_ ), .ZN(_06205_ ) );
NAND4_X1 _13983_ ( .A1(_06202_ ), .A2(_06203_ ), .A3(_06204_ ), .A4(_06205_ ), .ZN(_06206_ ) );
OAI21_X1 _13984_ ( .A(_06051_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_06207_ ) );
INV_X1 _13985_ ( .A(_06207_ ), .ZN(_06208_ ) );
NAND3_X1 _13986_ ( .A1(_06203_ ), .A2(_06204_ ), .A3(_06208_ ), .ZN(_06209_ ) );
NAND2_X1 _13987_ ( .A1(_06052_ ), .A2(\IF_ID_pc [28] ), .ZN(_06210_ ) );
AND2_X1 _13988_ ( .A1(_06052_ ), .A2(\IF_ID_pc [27] ), .ZN(_06211_ ) );
INV_X1 _13989_ ( .A(_06211_ ), .ZN(_06212_ ) );
AND3_X1 _13990_ ( .A1(_06209_ ), .A2(_06210_ ), .A3(_06212_ ), .ZN(_06213_ ) );
AOI21_X1 _13991_ ( .A(_06054_ ), .B1(_06206_ ), .B2(_06213_ ), .ZN(_06214_ ) );
NOR3_X1 _13992_ ( .A1(_06047_ ), .A2(_02064_ ), .A3(_06049_ ), .ZN(_06215_ ) );
OR2_X1 _13993_ ( .A1(_06214_ ), .A2(_06215_ ), .ZN(_06216_ ) );
XNOR2_X1 _13994_ ( .A(_06052_ ), .B(_02264_ ), .ZN(_06217_ ) );
XNOR2_X1 _13995_ ( .A(_06216_ ), .B(_06217_ ), .ZN(_06218_ ) );
BUF_X4 _13996_ ( .A(_05915_ ), .Z(_06219_ ) );
INV_X2 _13997_ ( .A(_06219_ ), .ZN(_06220_ ) );
BUF_X4 _13998_ ( .A(_06220_ ), .Z(_06221_ ) );
MUX2_X1 _13999_ ( .A(_02395_ ), .B(_06218_ ), .S(_06221_ ), .Z(_06222_ ) );
BUF_X4 _14000_ ( .A(_06039_ ), .Z(_06223_ ) );
AOI211_X1 _14001_ ( .A(fanout_net_3 ), .B(_06043_ ), .C1(_06222_ ), .C2(_06223_ ), .ZN(_00246_ ) );
NOR2_X1 _14002_ ( .A1(_06040_ ), .A2(\mtvec [21] ), .ZN(_06224_ ) );
AOI211_X1 _14003_ ( .A(_06188_ ), .B(_06172_ ), .C1(_06191_ ), .C2(_06189_ ), .ZN(_06225_ ) );
NAND3_X1 _14004_ ( .A1(_06143_ ), .A2(_06157_ ), .A3(_06158_ ), .ZN(_06226_ ) );
INV_X1 _14005_ ( .A(_06226_ ), .ZN(_06227_ ) );
OR3_X2 _14006_ ( .A1(_06227_ ), .A2(_06147_ ), .A3(_06151_ ), .ZN(_06228_ ) );
NAND2_X1 _14007_ ( .A1(_06157_ ), .A2(_06158_ ), .ZN(_06229_ ) );
NOR2_X1 _14008_ ( .A1(_06154_ ), .A2(_06229_ ), .ZN(_06230_ ) );
OAI21_X1 _14009_ ( .A(_06178_ ), .B1(_06228_ ), .B2(_06230_ ), .ZN(_06231_ ) );
INV_X1 _14010_ ( .A(_06175_ ), .ZN(_06232_ ) );
OR2_X1 _14011_ ( .A1(_06231_ ), .A2(_06232_ ), .ZN(_06233_ ) );
NAND2_X1 _14012_ ( .A1(_06186_ ), .A2(_06183_ ), .ZN(_06234_ ) );
AOI21_X1 _14013_ ( .A(_06188_ ), .B1(_06189_ ), .B2(_06191_ ), .ZN(_06235_ ) );
AND2_X1 _14014_ ( .A1(_06234_ ), .A2(_06235_ ), .ZN(_06236_ ) );
AOI21_X1 _14015_ ( .A(_06225_ ), .B1(_06233_ ), .B2(_06236_ ), .ZN(_06237_ ) );
XNOR2_X1 _14016_ ( .A(_06237_ ), .B(_06162_ ), .ZN(_06238_ ) );
MUX2_X1 _14017_ ( .A(_05635_ ), .B(_06238_ ), .S(_06221_ ), .Z(_06239_ ) );
AOI211_X1 _14018_ ( .A(fanout_net_3 ), .B(_06224_ ), .C1(_06239_ ), .C2(_06223_ ), .ZN(_00247_ ) );
AND3_X1 _14019_ ( .A1(_06037_ ), .A2(check_quest ), .A3(\myexu.pc_jump [20] ), .ZN(_06240_ ) );
NAND2_X1 _14020_ ( .A1(_06233_ ), .A2(_06234_ ), .ZN(_06241_ ) );
AND2_X1 _14021_ ( .A1(_06241_ ), .A2(_06170_ ), .ZN(_06242_ ) );
NOR2_X1 _14022_ ( .A1(_06242_ ), .A2(_06189_ ), .ZN(_06243_ ) );
XNOR2_X1 _14023_ ( .A(_06243_ ), .B(_06171_ ), .ZN(_06244_ ) );
AOI211_X1 _14024_ ( .A(\myifu.to_reset ), .B(_06240_ ), .C1(_06244_ ), .C2(_06221_ ), .ZN(_06245_ ) );
INV_X1 _14025_ ( .A(\mtvec [20] ), .ZN(_06246_ ) );
AOI211_X1 _14026_ ( .A(fanout_net_3 ), .B(_06245_ ), .C1(_06246_ ), .C2(\myifu.to_reset ), .ZN(_00248_ ) );
BUF_X4 _14027_ ( .A(_06039_ ), .Z(_06247_ ) );
NAND3_X1 _14028_ ( .A1(_05902_ ), .A2(_05908_ ), .A3(_05913_ ), .ZN(_06248_ ) );
NAND4_X1 _14029_ ( .A1(_05876_ ), .A2(_05881_ ), .A3(_05886_ ), .A4(_05892_ ), .ZN(_06249_ ) );
OAI211_X1 _14030_ ( .A(check_quest ), .B(_04918_ ), .C1(_06248_ ), .C2(_06249_ ), .ZN(_06250_ ) );
XOR2_X1 _14031_ ( .A(_06241_ ), .B(_06170_ ), .Z(_06251_ ) );
BUF_X4 _14032_ ( .A(_06219_ ), .Z(_06252_ ) );
OAI211_X1 _14033_ ( .A(_06247_ ), .B(_06250_ ), .C1(_06251_ ), .C2(_06252_ ), .ZN(_06253_ ) );
NAND2_X1 _14034_ ( .A1(\mtvec [19] ), .A2(\myifu.to_reset ), .ZN(_06254_ ) );
AOI21_X1 _14035_ ( .A(fanout_net_3 ), .B1(_06253_ ), .B2(_06254_ ), .ZN(_00249_ ) );
AND2_X1 _14036_ ( .A1(_06160_ ), .A2(_06178_ ), .ZN(_06255_ ) );
OR3_X1 _14037_ ( .A1(_06255_ ), .A2(_06185_ ), .A3(_06232_ ), .ZN(_06256_ ) );
BUF_X4 _14038_ ( .A(_06220_ ), .Z(_06257_ ) );
OAI21_X1 _14039_ ( .A(_06232_ ), .B1(_06255_ ), .B2(_06185_ ), .ZN(_06258_ ) );
NAND3_X1 _14040_ ( .A1(_06256_ ), .A2(_06257_ ), .A3(_06258_ ), .ZN(_06259_ ) );
OAI211_X1 _14041_ ( .A(_06259_ ), .B(_06040_ ), .C1(\myexu.pc_jump [18] ), .C2(_06257_ ), .ZN(_06260_ ) );
NAND2_X1 _14042_ ( .A1(\mtvec [18] ), .A2(\myifu.to_reset ), .ZN(_06261_ ) );
AOI21_X1 _14043_ ( .A(fanout_net_3 ), .B1(_06260_ ), .B2(_06261_ ), .ZN(_00250_ ) );
NOR2_X1 _14044_ ( .A1(_06040_ ), .A2(\mtvec [17] ), .ZN(_06262_ ) );
XNOR2_X1 _14045_ ( .A(_06160_ ), .B(_06178_ ), .ZN(_06263_ ) );
MUX2_X1 _14046_ ( .A(_05002_ ), .B(_06263_ ), .S(_06221_ ), .Z(_06264_ ) );
AOI211_X1 _14047_ ( .A(fanout_net_3 ), .B(_06262_ ), .C1(_06264_ ), .C2(_06223_ ), .ZN(_00251_ ) );
OR3_X1 _14048_ ( .A1(_05914_ ), .A2(_02417_ ), .A3(\myexu.pc_jump [16] ), .ZN(_06265_ ) );
OAI21_X1 _14049_ ( .A(_06158_ ), .B1(_06143_ ), .B2(_06155_ ), .ZN(_06266_ ) );
OR2_X1 _14050_ ( .A1(_06150_ ), .A2(_02150_ ), .ZN(_06267_ ) );
AND2_X1 _14051_ ( .A1(_06266_ ), .A2(_06267_ ), .ZN(_06268_ ) );
XNOR2_X1 _14052_ ( .A(_06268_ ), .B(_06157_ ), .ZN(_06269_ ) );
OAI211_X1 _14053_ ( .A(_06247_ ), .B(_06265_ ), .C1(_06269_ ), .C2(_06252_ ), .ZN(_06270_ ) );
NAND2_X1 _14054_ ( .A1(\mtvec [16] ), .A2(\myifu.to_reset ), .ZN(_06271_ ) );
AOI21_X1 _14055_ ( .A(fanout_net_3 ), .B1(_06270_ ), .B2(_06271_ ), .ZN(_00252_ ) );
NOR2_X1 _14056_ ( .A1(_06143_ ), .A2(_06155_ ), .ZN(_06272_ ) );
XOR2_X1 _14057_ ( .A(_06272_ ), .B(_06158_ ), .Z(_06273_ ) );
NAND2_X1 _14058_ ( .A1(_06273_ ), .A2(_06257_ ), .ZN(_06274_ ) );
OAI211_X1 _14059_ ( .A(_06274_ ), .B(_06040_ ), .C1(\myexu.pc_jump [15] ), .C2(_06257_ ), .ZN(_06275_ ) );
NAND2_X1 _14060_ ( .A1(\mtvec [15] ), .A2(\myifu.to_reset ), .ZN(_06276_ ) );
AOI21_X1 _14061_ ( .A(fanout_net_3 ), .B1(_06275_ ), .B2(_06276_ ), .ZN(_00253_ ) );
OR3_X1 _14062_ ( .A1(_05914_ ), .A2(_02417_ ), .A3(\myexu.pc_jump [14] ), .ZN(_06277_ ) );
NOR2_X1 _14063_ ( .A1(_06134_ ), .A2(_06135_ ), .ZN(_06278_ ) );
AND2_X1 _14064_ ( .A1(_06278_ ), .A2(_06141_ ), .ZN(_06279_ ) );
NOR2_X1 _14065_ ( .A1(_06279_ ), .A2(_06153_ ), .ZN(_06280_ ) );
XNOR2_X1 _14066_ ( .A(_06280_ ), .B(_06138_ ), .ZN(_06281_ ) );
OAI211_X1 _14067_ ( .A(_06247_ ), .B(_06277_ ), .C1(_06281_ ), .C2(_06252_ ), .ZN(_06282_ ) );
NAND2_X1 _14068_ ( .A1(\mtvec [14] ), .A2(\myifu.to_reset ), .ZN(_06283_ ) );
AOI21_X1 _14069_ ( .A(fanout_net_3 ), .B1(_06282_ ), .B2(_06283_ ), .ZN(_00254_ ) );
XOR2_X1 _14070_ ( .A(_06278_ ), .B(_06141_ ), .Z(_06284_ ) );
MUX2_X1 _14071_ ( .A(\myexu.pc_jump [13] ), .B(_06284_ ), .S(_06220_ ), .Z(_06285_ ) );
MUX2_X1 _14072_ ( .A(\mtvec [13] ), .B(_06285_ ), .S(_06038_ ), .Z(_06286_ ) );
AND2_X1 _14073_ ( .A1(_06286_ ), .A2(_03400_ ), .ZN(_00255_ ) );
INV_X1 _14074_ ( .A(\mtvec [12] ), .ZN(_06287_ ) );
NOR2_X1 _14075_ ( .A1(_06128_ ), .A2(_06133_ ), .ZN(_06288_ ) );
XNOR2_X1 _14076_ ( .A(_06131_ ), .B(\IF_ID_pc [12] ), .ZN(_06289_ ) );
AOI21_X1 _14077_ ( .A(_06219_ ), .B1(_06288_ ), .B2(_06289_ ), .ZN(_06290_ ) );
OAI21_X1 _14078_ ( .A(_06290_ ), .B1(_06288_ ), .B2(_06289_ ), .ZN(_06291_ ) );
AOI21_X1 _14079_ ( .A(\myifu.to_reset ), .B1(_06219_ ), .B2(\myexu.pc_jump [12] ), .ZN(_06292_ ) );
AOI221_X4 _14080_ ( .A(fanout_net_3 ), .B1(_06287_ ), .B2(\myifu.to_reset ), .C1(_06291_ ), .C2(_06292_ ), .ZN(_00256_ ) );
NOR2_X1 _14081_ ( .A1(_06040_ ), .A2(\mtvec [29] ), .ZN(_06293_ ) );
AND2_X1 _14082_ ( .A1(_06206_ ), .A2(_06213_ ), .ZN(_06294_ ) );
XNOR2_X1 _14083_ ( .A(_06294_ ), .B(_06054_ ), .ZN(_06295_ ) );
MUX2_X1 _14084_ ( .A(_02396_ ), .B(_06295_ ), .S(_06221_ ), .Z(_06296_ ) );
AOI211_X1 _14085_ ( .A(fanout_net_3 ), .B(_06293_ ), .C1(_06296_ ), .C2(_06223_ ), .ZN(_00257_ ) );
AOI21_X1 _14086_ ( .A(_06125_ ), .B1(_06121_ ), .B2(_06127_ ), .ZN(_06297_ ) );
OAI21_X1 _14087_ ( .A(_06221_ ), .B1(_06128_ ), .B2(_06297_ ), .ZN(_06298_ ) );
OAI211_X1 _14088_ ( .A(_06298_ ), .B(_06040_ ), .C1(\myexu.pc_jump [11] ), .C2(_06257_ ), .ZN(_06299_ ) );
NAND2_X1 _14089_ ( .A1(\mtvec [11] ), .A2(\myifu.to_reset ), .ZN(_06300_ ) );
AOI21_X1 _14090_ ( .A(fanout_net_3 ), .B1(_06299_ ), .B2(_06300_ ), .ZN(_00258_ ) );
NOR2_X1 _14091_ ( .A1(_06039_ ), .A2(\mtvec [10] ), .ZN(_06301_ ) );
NOR2_X1 _14092_ ( .A1(_06114_ ), .A2(_06120_ ), .ZN(_06302_ ) );
XNOR2_X1 _14093_ ( .A(_06117_ ), .B(_02208_ ), .ZN(_06303_ ) );
XOR2_X1 _14094_ ( .A(_06302_ ), .B(_06303_ ), .Z(_06304_ ) );
MUX2_X1 _14095_ ( .A(_05220_ ), .B(_06304_ ), .S(_06221_ ), .Z(_06305_ ) );
AOI211_X1 _14096_ ( .A(fanout_net_3 ), .B(_06301_ ), .C1(_06305_ ), .C2(_06223_ ), .ZN(_00259_ ) );
AND3_X1 _14097_ ( .A1(_06112_ ), .A2(_06113_ ), .A3(_06061_ ), .ZN(_06306_ ) );
OAI21_X1 _14098_ ( .A(_06221_ ), .B1(_06306_ ), .B2(_06114_ ), .ZN(_06307_ ) );
OAI211_X1 _14099_ ( .A(_06307_ ), .B(_06040_ ), .C1(\myexu.pc_jump [9] ), .C2(_06257_ ), .ZN(_06308_ ) );
NAND2_X1 _14100_ ( .A1(\mtvec [9] ), .A2(\myifu.to_reset ), .ZN(_06309_ ) );
AOI21_X1 _14101_ ( .A(fanout_net_3 ), .B1(_06308_ ), .B2(_06309_ ), .ZN(_00260_ ) );
NOR2_X1 _14102_ ( .A1(_06039_ ), .A2(\mtvec [8] ), .ZN(_06310_ ) );
NOR2_X1 _14103_ ( .A1(_06106_ ), .A2(_06107_ ), .ZN(_06311_ ) );
XNOR2_X1 _14104_ ( .A(_06110_ ), .B(_02233_ ), .ZN(_06312_ ) );
XNOR2_X1 _14105_ ( .A(_06311_ ), .B(_06312_ ), .ZN(_06313_ ) );
MUX2_X1 _14106_ ( .A(_05269_ ), .B(_06313_ ), .S(_06221_ ), .Z(_06314_ ) );
AOI211_X1 _14107_ ( .A(fanout_net_3 ), .B(_06310_ ), .C1(_06314_ ), .C2(_06223_ ), .ZN(_00261_ ) );
OR3_X1 _14108_ ( .A1(_05914_ ), .A2(_02417_ ), .A3(\myexu.pc_jump [7] ), .ZN(_06315_ ) );
NAND2_X1 _14109_ ( .A1(_06100_ ), .A2(_06105_ ), .ZN(_06316_ ) );
XNOR2_X1 _14110_ ( .A(_06316_ ), .B(_06104_ ), .ZN(_06317_ ) );
OAI211_X1 _14111_ ( .A(_06247_ ), .B(_06315_ ), .C1(_06317_ ), .C2(_06252_ ), .ZN(_06318_ ) );
NAND2_X1 _14112_ ( .A1(\mtvec [7] ), .A2(\myifu.to_reset ), .ZN(_06319_ ) );
AOI21_X1 _14113_ ( .A(fanout_net_3 ), .B1(_06318_ ), .B2(_06319_ ), .ZN(_00262_ ) );
NOR2_X1 _14114_ ( .A1(_06097_ ), .A2(_06099_ ), .ZN(_06320_ ) );
NOR2_X1 _14115_ ( .A1(_06070_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06321_ ) );
XNOR2_X1 _14116_ ( .A(_06065_ ), .B(\IF_ID_pc [6] ), .ZN(_06322_ ) );
OR3_X1 _14117_ ( .A1(_06320_ ), .A2(_06321_ ), .A3(_06322_ ), .ZN(_06323_ ) );
OAI21_X1 _14118_ ( .A(_06322_ ), .B1(_06320_ ), .B2(_06321_ ), .ZN(_06324_ ) );
AOI21_X1 _14119_ ( .A(_06219_ ), .B1(_06323_ ), .B2(_06324_ ), .ZN(_06325_ ) );
AOI211_X1 _14120_ ( .A(\myifu.to_reset ), .B(_06325_ ), .C1(\myexu.pc_jump [6] ), .C2(_06252_ ), .ZN(_06326_ ) );
INV_X1 _14121_ ( .A(\mtvec [6] ), .ZN(_06327_ ) );
AOI211_X1 _14122_ ( .A(fanout_net_3 ), .B(_06326_ ), .C1(_06327_ ), .C2(\myifu.to_reset ), .ZN(_00263_ ) );
NOR2_X1 _14123_ ( .A1(_06039_ ), .A2(\mtvec [5] ), .ZN(_06328_ ) );
XNOR2_X1 _14124_ ( .A(_06097_ ), .B(_06099_ ), .ZN(_06329_ ) );
MUX2_X1 _14125_ ( .A(_05347_ ), .B(_06329_ ), .S(_06220_ ), .Z(_06330_ ) );
AOI211_X1 _14126_ ( .A(fanout_net_3 ), .B(_06328_ ), .C1(_06330_ ), .C2(_06223_ ), .ZN(_00264_ ) );
INV_X1 _14127_ ( .A(_06093_ ), .ZN(_06331_ ) );
OAI21_X1 _14128_ ( .A(_06331_ ), .B1(_06091_ ), .B2(_06083_ ), .ZN(_06332_ ) );
AND2_X1 _14129_ ( .A1(_06074_ ), .A2(_06096_ ), .ZN(_06333_ ) );
AND3_X1 _14130_ ( .A1(_06332_ ), .A2(_06080_ ), .A3(_06333_ ), .ZN(_06334_ ) );
AOI21_X1 _14131_ ( .A(_06333_ ), .B1(_06332_ ), .B2(_06080_ ), .ZN(_06335_ ) );
OR3_X1 _14132_ ( .A1(_06334_ ), .A2(_06335_ ), .A3(_06219_ ), .ZN(_06336_ ) );
OAI211_X1 _14133_ ( .A(_06336_ ), .B(_06038_ ), .C1(\myexu.pc_jump [4] ), .C2(_06220_ ), .ZN(_06337_ ) );
NAND2_X1 _14134_ ( .A1(\mtvec [4] ), .A2(\myifu.to_reset ), .ZN(_06338_ ) );
AOI21_X1 _14135_ ( .A(fanout_net_3 ), .B1(_06337_ ), .B2(_06338_ ), .ZN(_00265_ ) );
AND2_X1 _14136_ ( .A1(\mtvec [3] ), .A2(\myifu.to_reset ), .ZN(_06339_ ) );
XNOR2_X1 _14137_ ( .A(_06092_ ), .B(_06331_ ), .ZN(_06340_ ) );
MUX2_X1 _14138_ ( .A(\myexu.pc_jump [3] ), .B(_06340_ ), .S(_06220_ ), .Z(_06341_ ) );
AOI21_X1 _14139_ ( .A(_06339_ ), .B1(_06341_ ), .B2(_06247_ ), .ZN(_06342_ ) );
NOR2_X1 _14140_ ( .A1(_06342_ ), .A2(fanout_net_3 ), .ZN(_00266_ ) );
AND2_X1 _14141_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
AND3_X1 _14142_ ( .A1(_06337_ ), .A2(_06338_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_06343_ ) );
CLKBUF_X2 _14143_ ( .A(_06095_ ), .Z(_06344_ ) );
CLKBUF_X2 _14144_ ( .A(_06344_ ), .Z(_06345_ ) );
BUF_X2 _14145_ ( .A(_06345_ ), .Z(_06346_ ) );
INV_X1 _14146_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_06347_ ) );
AOI211_X1 _14147_ ( .A(reset ), .B(_06343_ ), .C1(_06346_ ), .C2(_06347_ ), .ZN(_00267_ ) );
NOR2_X1 _14148_ ( .A1(_06039_ ), .A2(\mtvec [2] ), .ZN(_06348_ ) );
XNOR2_X1 _14149_ ( .A(_06085_ ), .B(_06090_ ), .ZN(_06349_ ) );
MUX2_X1 _14150_ ( .A(_06349_ ), .B(_05425_ ), .S(_06219_ ), .Z(_06350_ ) );
AOI211_X1 _14151_ ( .A(reset ), .B(_06348_ ), .C1(_06350_ ), .C2(_06223_ ), .ZN(_00268_ ) );
AOI211_X1 _14152_ ( .A(_06339_ ), .B(_06347_ ), .C1(_06341_ ), .C2(_06039_ ), .ZN(_06351_ ) );
INV_X1 _14153_ ( .A(fanout_net_8 ), .ZN(_06352_ ) );
BUF_X4 _14154_ ( .A(_06352_ ), .Z(_06353_ ) );
BUF_X4 _14155_ ( .A(_06353_ ), .Z(_06354_ ) );
BUF_X2 _14156_ ( .A(_06354_ ), .Z(_06355_ ) );
AOI211_X1 _14157_ ( .A(reset ), .B(_06351_ ), .C1(_06355_ ), .C2(_06347_ ), .ZN(_00269_ ) );
INV_X1 _14158_ ( .A(\mtvec [28] ), .ZN(_06356_ ) );
INV_X1 _14159_ ( .A(_06201_ ), .ZN(_06357_ ) );
NOR2_X1 _14160_ ( .A1(_06180_ ), .A2(_06357_ ), .ZN(_06358_ ) );
INV_X1 _14161_ ( .A(_06205_ ), .ZN(_06359_ ) );
NOR3_X1 _14162_ ( .A1(_06358_ ), .A2(_06359_ ), .A3(_06056_ ), .ZN(_06360_ ) );
OAI21_X1 _14163_ ( .A(_06204_ ), .B1(_06360_ ), .B2(_06208_ ), .ZN(_06361_ ) );
AND3_X1 _14164_ ( .A1(_06361_ ), .A2(_06203_ ), .A3(_06212_ ), .ZN(_06362_ ) );
AOI21_X1 _14165_ ( .A(_06203_ ), .B1(_06361_ ), .B2(_06212_ ), .ZN(_06363_ ) );
OAI21_X1 _14166_ ( .A(_06220_ ), .B1(_06362_ ), .B2(_06363_ ), .ZN(_06364_ ) );
AOI21_X1 _14167_ ( .A(\myifu.to_reset ), .B1(_06219_ ), .B2(\myexu.pc_jump [28] ), .ZN(_06365_ ) );
AOI221_X4 _14168_ ( .A(reset ), .B1(_06356_ ), .B2(\myifu.to_reset ), .C1(_06364_ ), .C2(_06365_ ), .ZN(_00270_ ) );
NOR2_X1 _14169_ ( .A1(_06039_ ), .A2(\mtvec [1] ), .ZN(_06366_ ) );
XNOR2_X1 _14170_ ( .A(_06089_ ), .B(\IF_ID_pc [1] ), .ZN(_06367_ ) );
MUX2_X1 _14171_ ( .A(_06367_ ), .B(_05445_ ), .S(_06219_ ), .Z(_06368_ ) );
AOI211_X1 _14172_ ( .A(reset ), .B(_06366_ ), .C1(_06368_ ), .C2(_06223_ ), .ZN(_00271_ ) );
OAI211_X1 _14173_ ( .A(check_quest ), .B(_05473_ ), .C1(_06248_ ), .C2(_06249_ ), .ZN(_06369_ ) );
NOR2_X1 _14174_ ( .A1(_06360_ ), .A2(_06208_ ), .ZN(_06370_ ) );
XNOR2_X1 _14175_ ( .A(_06370_ ), .B(_06204_ ), .ZN(_06371_ ) );
OAI211_X1 _14176_ ( .A(_06247_ ), .B(_06369_ ), .C1(_06371_ ), .C2(_06252_ ), .ZN(_06372_ ) );
NAND2_X1 _14177_ ( .A1(\mtvec [27] ), .A2(\myifu.to_reset ), .ZN(_06373_ ) );
AOI21_X1 _14178_ ( .A(reset ), .B1(_06372_ ), .B2(_06373_ ), .ZN(_00272_ ) );
NOR2_X1 _14179_ ( .A1(_06039_ ), .A2(\mtvec [26] ), .ZN(_06374_ ) );
AND2_X1 _14180_ ( .A1(_06052_ ), .A2(\IF_ID_pc [25] ), .ZN(_06375_ ) );
NOR2_X1 _14181_ ( .A1(_06202_ ), .A2(_06375_ ), .ZN(_06376_ ) );
XNOR2_X1 _14182_ ( .A(_06376_ ), .B(_06359_ ), .ZN(_06377_ ) );
MUX2_X1 _14183_ ( .A(_02391_ ), .B(_06377_ ), .S(_06220_ ), .Z(_06378_ ) );
AOI211_X1 _14184_ ( .A(reset ), .B(_06374_ ), .C1(_06378_ ), .C2(_06223_ ), .ZN(_00273_ ) );
OAI211_X1 _14185_ ( .A(check_quest ), .B(_02392_ ), .C1(_06248_ ), .C2(_06249_ ), .ZN(_06379_ ) );
XNOR2_X1 _14186_ ( .A(_06358_ ), .B(_06055_ ), .ZN(_06380_ ) );
OAI211_X1 _14187_ ( .A(_06247_ ), .B(_06379_ ), .C1(_06380_ ), .C2(_06252_ ), .ZN(_06381_ ) );
NAND2_X1 _14188_ ( .A1(\mtvec [25] ), .A2(\myifu.to_reset ), .ZN(_06382_ ) );
AOI21_X1 _14189_ ( .A(reset ), .B1(_06381_ ), .B2(_06382_ ), .ZN(_00274_ ) );
INV_X1 _14190_ ( .A(\mtvec [24] ), .ZN(_06383_ ) );
AND2_X1 _14191_ ( .A1(_06237_ ), .A2(_06162_ ), .ZN(_06384_ ) );
NOR2_X2 _14192_ ( .A1(_06384_ ), .A2(_06196_ ), .ZN(_06385_ ) );
INV_X1 _14193_ ( .A(_06052_ ), .ZN(_06386_ ) );
AOI21_X1 _14194_ ( .A(_06385_ ), .B1(_02166_ ), .B2(_06386_ ), .ZN(_06387_ ) );
OAI21_X1 _14195_ ( .A(_06165_ ), .B1(_06387_ ), .B2(_06195_ ), .ZN(_06388_ ) );
AND3_X1 _14196_ ( .A1(_06388_ ), .A2(_06164_ ), .A3(_06199_ ), .ZN(_06389_ ) );
AOI21_X1 _14197_ ( .A(_06164_ ), .B1(_06388_ ), .B2(_06199_ ), .ZN(_06390_ ) );
OAI21_X1 _14198_ ( .A(_06220_ ), .B1(_06389_ ), .B2(_06390_ ), .ZN(_06391_ ) );
AOI21_X1 _14199_ ( .A(\myifu.to_reset ), .B1(_06219_ ), .B2(\myexu.pc_jump [24] ), .ZN(_06392_ ) );
AOI221_X1 _14200_ ( .A(reset ), .B1(_06383_ ), .B2(\myifu.to_reset ), .C1(_06391_ ), .C2(_06392_ ), .ZN(_00275_ ) );
OAI211_X1 _14201_ ( .A(check_quest ), .B(_05587_ ), .C1(_06248_ ), .C2(_06249_ ), .ZN(_06393_ ) );
OR2_X1 _14202_ ( .A1(_06387_ ), .A2(_06195_ ), .ZN(_06394_ ) );
XOR2_X1 _14203_ ( .A(_06394_ ), .B(_06165_ ), .Z(_06395_ ) );
OAI211_X1 _14204_ ( .A(_06247_ ), .B(_06393_ ), .C1(_06395_ ), .C2(_06252_ ), .ZN(_06396_ ) );
NAND2_X1 _14205_ ( .A1(\mtvec [23] ), .A2(\myifu.to_reset ), .ZN(_06397_ ) );
AOI21_X1 _14206_ ( .A(reset ), .B1(_06396_ ), .B2(_06397_ ), .ZN(_00276_ ) );
AND3_X1 _14207_ ( .A1(_06037_ ), .A2(check_quest ), .A3(\myexu.pc_jump [22] ), .ZN(_06398_ ) );
XNOR2_X1 _14208_ ( .A(_06385_ ), .B(_06161_ ), .ZN(_06399_ ) );
AOI211_X1 _14209_ ( .A(\myifu.to_reset ), .B(_06398_ ), .C1(_06399_ ), .C2(_06257_ ), .ZN(_06400_ ) );
NOR2_X1 _14210_ ( .A1(_06247_ ), .A2(\mtvec [22] ), .ZN(_06401_ ) );
NOR3_X1 _14211_ ( .A1(_06400_ ), .A2(reset ), .A3(_06401_ ), .ZN(_00277_ ) );
INV_X1 _14212_ ( .A(\mtvec [31] ), .ZN(_06402_ ) );
OAI22_X1 _14213_ ( .A1(_06214_ ), .A2(_06215_ ), .B1(\IF_ID_pc [30] ), .B2(_06052_ ), .ZN(_06403_ ) );
NAND2_X1 _14214_ ( .A1(_06052_ ), .A2(\IF_ID_pc [30] ), .ZN(_06404_ ) );
NAND2_X1 _14215_ ( .A1(_06403_ ), .A2(_06404_ ), .ZN(_06405_ ) );
XNOR2_X1 _14216_ ( .A(_06052_ ), .B(\IF_ID_pc [31] ), .ZN(_06406_ ) );
AND2_X1 _14217_ ( .A1(_06405_ ), .A2(_06406_ ), .ZN(_06407_ ) );
OAI21_X1 _14218_ ( .A(_06221_ ), .B1(_06405_ ), .B2(_06406_ ), .ZN(_06408_ ) );
NOR2_X1 _14219_ ( .A1(_06407_ ), .A2(_06408_ ), .ZN(_06409_ ) );
OAI21_X1 _14220_ ( .A(_06040_ ), .B1(_06257_ ), .B2(\myexu.pc_jump [31] ), .ZN(_06410_ ) );
OAI221_X1 _14221_ ( .A(_03400_ ), .B1(_06402_ ), .B2(_06247_ ), .C1(_06409_ ), .C2(_06410_ ), .ZN(_00278_ ) );
AND3_X1 _14222_ ( .A1(_02296_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .A3(_02316_ ), .ZN(_06411_ ) );
NOR2_X1 _14223_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_06412_ ) );
NAND2_X1 _14224_ ( .A1(_06412_ ), .A2(io_master_rvalid ), .ZN(_06413_ ) );
AOI21_X1 _14225_ ( .A(_06411_ ), .B1(_02318_ ), .B2(_06413_ ), .ZN(_06414_ ) );
OR2_X1 _14226_ ( .A1(_02317_ ), .A2(io_master_rlast ), .ZN(_06415_ ) );
AND3_X1 _14227_ ( .A1(_06414_ ), .A2(_02321_ ), .A3(_06415_ ), .ZN(_06416_ ) );
INV_X1 _14228_ ( .A(\io_master_rid [3] ), .ZN(_06417_ ) );
INV_X1 _14229_ ( .A(\io_master_rid [2] ), .ZN(_06418_ ) );
INV_X1 _14230_ ( .A(\io_master_rid [1] ), .ZN(_06419_ ) );
NAND4_X1 _14231_ ( .A1(_06417_ ), .A2(_06418_ ), .A3(_06419_ ), .A4(\io_master_rid [0] ), .ZN(_06420_ ) );
AOI21_X1 _14232_ ( .A(_02293_ ), .B1(_02318_ ), .B2(_06420_ ), .ZN(_06421_ ) );
NAND2_X1 _14233_ ( .A1(_06416_ ), .A2(_06421_ ), .ZN(_06422_ ) );
INV_X1 _14234_ ( .A(\myifu.tmp_offset [2] ), .ZN(_06423_ ) );
NAND3_X1 _14235_ ( .A1(_06422_ ), .A2(_03400_ ), .A3(_06423_ ), .ZN(_06424_ ) );
INV_X1 _14236_ ( .A(_06424_ ), .ZN(_00279_ ) );
NOR3_X1 _14237_ ( .A1(reset ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00280_ ) );
AND3_X1 _14238_ ( .A1(_02388_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .A3(_05916_ ), .ZN(_06425_ ) );
INV_X1 _14239_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_06426_ ) );
MUX2_X1 _14240_ ( .A(_02388_ ), .B(_06426_ ), .S(\myifu.to_reset ), .Z(_06427_ ) );
AOI211_X1 _14241_ ( .A(reset ), .B(_06425_ ), .C1(_06427_ ), .C2(\myifu.state [1] ), .ZN(_00281_ ) );
INV_X1 _14242_ ( .A(\myec.state [0] ), .ZN(_06428_ ) );
NOR2_X1 _14243_ ( .A1(_06428_ ), .A2(\myec.state [1] ), .ZN(_06429_ ) );
INV_X1 _14244_ ( .A(\EX_LS_pc [2] ), .ZN(_06430_ ) );
NOR3_X1 _14245_ ( .A1(_02404_ ), .A2(_06429_ ), .A3(_06430_ ), .ZN(_00282_ ) );
INV_X1 _14246_ ( .A(\mylsu.state [3] ), .ZN(_06431_ ) );
BUF_X4 _14247_ ( .A(_06431_ ), .Z(_06432_ ) );
NOR3_X1 _14248_ ( .A1(_02404_ ), .A2(_06429_ ), .A3(_06432_ ), .ZN(_00283_ ) );
BUF_X4 _14249_ ( .A(_02345_ ), .Z(_06433_ ) );
AOI21_X1 _14250_ ( .A(\LS_WB_waddr_csreg [11] ), .B1(_06433_ ), .B2(\EX_LS_flag [2] ), .ZN(_06434_ ) );
OR2_X1 _14251_ ( .A1(_02385_ ), .A2(_05683_ ), .ZN(_06435_ ) );
BUF_X4 _14252_ ( .A(_06435_ ), .Z(_06436_ ) );
NOR2_X1 _14253_ ( .A1(_02252_ ), .A2(\EX_LS_flag [1] ), .ZN(_06437_ ) );
OR2_X1 _14254_ ( .A1(_06437_ ), .A2(_02326_ ), .ZN(_06438_ ) );
NOR2_X1 _14255_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_06439_ ) );
AND2_X2 _14256_ ( .A1(_06439_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_06440_ ) );
NOR2_X2 _14257_ ( .A1(_06438_ ), .A2(_06440_ ), .ZN(_06441_ ) );
NAND2_X1 _14258_ ( .A1(_06436_ ), .A2(_06441_ ), .ZN(_06442_ ) );
BUF_X4 _14259_ ( .A(_06442_ ), .Z(_06443_ ) );
BUF_X4 _14260_ ( .A(_06443_ ), .Z(_06444_ ) );
INV_X1 _14261_ ( .A(\EX_LS_dest_csreg_mem [11] ), .ZN(_06445_ ) );
BUF_X4 _14262_ ( .A(_04995_ ), .Z(_06446_ ) );
AOI211_X1 _14263_ ( .A(_06434_ ), .B(_06444_ ), .C1(_06445_ ), .C2(_06446_ ), .ZN(_00284_ ) );
NOR2_X1 _14264_ ( .A1(_02354_ ), .A2(_05683_ ), .ZN(_06447_ ) );
NOR2_X1 _14265_ ( .A1(_06447_ ), .A2(_06440_ ), .ZN(_06448_ ) );
INV_X1 _14266_ ( .A(_06448_ ), .ZN(_06449_ ) );
NAND3_X1 _14267_ ( .A1(_06433_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_06450_ ) );
BUF_X4 _14268_ ( .A(_02252_ ), .Z(_06451_ ) );
NAND2_X1 _14269_ ( .A1(_06451_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06452_ ) );
AOI211_X1 _14270_ ( .A(_05679_ ), .B(_06449_ ), .C1(_06450_ ), .C2(_06452_ ), .ZN(_00285_ ) );
NAND3_X1 _14271_ ( .A1(_06433_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_06453_ ) );
NAND2_X1 _14272_ ( .A1(_06451_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06454_ ) );
AOI211_X1 _14273_ ( .A(_05679_ ), .B(_06449_ ), .C1(_06453_ ), .C2(_06454_ ), .ZN(_00286_ ) );
NAND3_X1 _14274_ ( .A1(_06433_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_06455_ ) );
NAND2_X1 _14275_ ( .A1(_06451_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_06456_ ) );
AOI211_X1 _14276_ ( .A(_05679_ ), .B(_06449_ ), .C1(_06455_ ), .C2(_06456_ ), .ZN(_00287_ ) );
NAND3_X1 _14277_ ( .A1(_06433_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_06457_ ) );
NAND2_X1 _14278_ ( .A1(_06451_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06458_ ) );
AOI211_X1 _14279_ ( .A(_05679_ ), .B(_06449_ ), .C1(_06457_ ), .C2(_06458_ ), .ZN(_00288_ ) );
NAND3_X1 _14280_ ( .A1(_06433_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_06459_ ) );
NAND2_X1 _14281_ ( .A1(_06451_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_06460_ ) );
AOI211_X1 _14282_ ( .A(_05679_ ), .B(_06449_ ), .C1(_06459_ ), .C2(_06460_ ), .ZN(_00289_ ) );
NAND3_X1 _14283_ ( .A1(_06433_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_06461_ ) );
NAND2_X1 _14284_ ( .A1(_06451_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_06462_ ) );
AOI211_X1 _14285_ ( .A(_05679_ ), .B(_06449_ ), .C1(_06461_ ), .C2(_06462_ ), .ZN(_00290_ ) );
NAND3_X1 _14286_ ( .A1(_06433_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_flag [2] ), .ZN(_06463_ ) );
NAND2_X1 _14287_ ( .A1(_06451_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_06464_ ) );
AOI211_X1 _14288_ ( .A(_05679_ ), .B(_06449_ ), .C1(_06463_ ), .C2(_06464_ ), .ZN(_00291_ ) );
INV_X1 _14289_ ( .A(\EX_LS_flag [0] ), .ZN(_06465_ ) );
AND4_X1 _14290_ ( .A1(_04945_ ), .A2(_06465_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06466_ ) );
NOR2_X1 _14291_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_06467_ ) );
OAI211_X1 _14292_ ( .A(_06448_ ), .B(_05680_ ), .C1(_06466_ ), .C2(_06467_ ), .ZN(_00292_ ) );
INV_X1 _14293_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_06468_ ) );
AND4_X1 _14294_ ( .A1(_06468_ ), .A2(_06465_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06469_ ) );
NOR2_X1 _14295_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06470_ ) );
OAI211_X1 _14296_ ( .A(_06448_ ), .B(_05680_ ), .C1(_06469_ ), .C2(_06470_ ), .ZN(_00293_ ) );
INV_X1 _14297_ ( .A(\EX_LS_dest_csreg_mem [6] ), .ZN(_06471_ ) );
AND4_X1 _14298_ ( .A1(_06471_ ), .A2(_06465_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06472_ ) );
NOR2_X1 _14299_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06473_ ) );
OAI211_X1 _14300_ ( .A(_06448_ ), .B(_05680_ ), .C1(_06472_ ), .C2(_06473_ ), .ZN(_00294_ ) );
INV_X1 _14301_ ( .A(fanout_net_4 ), .ZN(_06474_ ) );
AND4_X1 _14302_ ( .A1(_06474_ ), .A2(_06465_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06475_ ) );
NOR2_X1 _14303_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_06476_ ) );
OAI211_X1 _14304_ ( .A(_06448_ ), .B(_05680_ ), .C1(_06475_ ), .C2(_06476_ ), .ZN(_00295_ ) );
NOR3_X1 _14305_ ( .A1(_02404_ ), .A2(_06429_ ), .A3(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06477_ ) );
NOR2_X1 _14306_ ( .A1(\mylsu.state [3] ), .A2(\mylsu.state [1] ), .ZN(_06478_ ) );
NAND2_X1 _14307_ ( .A1(_06477_ ), .A2(_06478_ ), .ZN(_06479_ ) );
BUF_X2 _14308_ ( .A(_02252_ ), .Z(_06480_ ) );
NOR2_X1 _14309_ ( .A1(_02399_ ), .A2(_02401_ ), .ZN(_06481_ ) );
AOI21_X1 _14310_ ( .A(_06480_ ), .B1(_06481_ ), .B2(_02344_ ), .ZN(_06482_ ) );
NOR3_X1 _14311_ ( .A1(_06447_ ), .A2(_06440_ ), .A3(_06482_ ), .ZN(_06483_ ) );
AOI21_X1 _14312_ ( .A(_06479_ ), .B1(_06483_ ), .B2(_02343_ ), .ZN(_00296_ ) );
INV_X1 _14313_ ( .A(_06433_ ), .ZN(_06484_ ) );
AOI21_X1 _14314_ ( .A(_02387_ ), .B1(_06484_ ), .B2(_06482_ ), .ZN(_06485_ ) );
AOI21_X1 _14315_ ( .A(_06479_ ), .B1(_06485_ ), .B2(_06448_ ), .ZN(_00297_ ) );
NAND3_X1 _14316_ ( .A1(_06481_ ), .A2(\EX_LS_flag [2] ), .A3(_02326_ ), .ZN(_06486_ ) );
NOR2_X1 _14317_ ( .A1(_06486_ ), .A2(_06479_ ), .ZN(_00298_ ) );
BUF_X4 _14318_ ( .A(_06436_ ), .Z(_06487_ ) );
AOI21_X1 _14319_ ( .A(_06479_ ), .B1(_06487_ ), .B2(_02343_ ), .ZN(_00299_ ) );
AOI21_X1 _14320_ ( .A(_06479_ ), .B1(_06448_ ), .B2(_06486_ ), .ZN(_00300_ ) );
NOR3_X1 _14321_ ( .A1(_06440_ ), .A2(_02404_ ), .A3(_06429_ ), .ZN(_06488_ ) );
NOR3_X1 _14322_ ( .A1(_05678_ ), .A2(\mylsu.state [3] ), .A3(\mylsu.state [1] ), .ZN(_06489_ ) );
NAND3_X1 _14323_ ( .A1(_02384_ ), .A2(_06488_ ), .A3(_06489_ ), .ZN(_06490_ ) );
INV_X1 _14324_ ( .A(_02342_ ), .ZN(_06491_ ) );
NOR3_X1 _14325_ ( .A1(_02401_ ), .A2(_06433_ ), .A3(_02252_ ), .ZN(_06492_ ) );
OAI21_X1 _14326_ ( .A(_06492_ ), .B1(_02399_ ), .B2(\EX_LS_flag [1] ), .ZN(_06493_ ) );
NOR2_X1 _14327_ ( .A1(_05677_ ), .A2(_06493_ ), .ZN(_06494_ ) );
OAI211_X1 _14328_ ( .A(_05679_ ), .B(_06491_ ), .C1(_06494_ ), .C2(_02325_ ), .ZN(_06495_ ) );
AND2_X1 _14329_ ( .A1(_02379_ ), .A2(_06493_ ), .ZN(_06496_ ) );
AOI21_X1 _14330_ ( .A(_06490_ ), .B1(_06495_ ), .B2(_06496_ ), .ZN(_00301_ ) );
INV_X1 _14331_ ( .A(_00283_ ), .ZN(_06497_ ) );
NOR2_X1 _14332_ ( .A1(_02404_ ), .A2(_06429_ ), .ZN(_06498_ ) );
NOR2_X1 _14333_ ( .A1(_06465_ ), .A2(\EX_LS_flag [1] ), .ZN(_06499_ ) );
OAI211_X1 _14334_ ( .A(_06498_ ), .B(_06489_ ), .C1(_06446_ ), .C2(_06499_ ), .ZN(_06500_ ) );
OAI21_X1 _14335_ ( .A(_06497_ ), .B1(_02347_ ), .B2(_06500_ ), .ZN(_00302_ ) );
INV_X1 _14336_ ( .A(\mysc.state [2] ), .ZN(_06501_ ) );
NOR2_X1 _14337_ ( .A1(_06501_ ), .A2(reset ), .ZN(_00303_ ) );
AND3_X1 _14338_ ( .A1(_01886_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00093_ ) );
AND2_X1 _14339_ ( .A1(_02357_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_06502_ ) );
CLKBUF_X2 _14340_ ( .A(_06502_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _14341_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .ZN(_06503_ ) );
BUF_X2 _14342_ ( .A(_06503_ ), .Z(_06504_ ) );
AND3_X1 _14343_ ( .A1(_02357_ ), .A2(_06504_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00242_ ) );
AND3_X1 _14344_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06346_ ), .A3(fanout_net_8 ), .ZN(_00243_ ) );
AND3_X1 _14345_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_12 ), .A3(_06355_ ), .ZN(_00244_ ) );
CLKBUF_X2 _14346_ ( .A(_02321_ ), .Z(\io_master_arburst [0] ) );
NOR3_X1 _14347_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(_05678_ ), .ZN(_06505_ ) );
BUF_X4 _14348_ ( .A(_05676_ ), .Z(_06506_ ) );
BUF_X4 _14349_ ( .A(_06506_ ), .Z(_06507_ ) );
INV_X1 _14350_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06508_ ) );
BUF_X4 _14351_ ( .A(_02274_ ), .Z(_06509_ ) );
INV_X1 _14352_ ( .A(_06509_ ), .ZN(_06510_ ) );
AOI211_X1 _14353_ ( .A(_06505_ ), .B(_06507_ ), .C1(_06508_ ), .C2(_06510_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _14354_ ( .A1(_02290_ ), .A2(fanout_net_4 ), .A3(_05678_ ), .ZN(_06511_ ) );
INV_X1 _14355_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06512_ ) );
AOI211_X1 _14356_ ( .A(_06511_ ), .B(_06507_ ), .C1(_06512_ ), .C2(_06510_ ), .ZN(\io_master_araddr [0] ) );
AND2_X2 _14357_ ( .A1(EXU_valid_LSU ), .A2(\mylsu.state [0] ), .ZN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _14358_ ( .A1(\EX_LS_dest_csreg_mem [15] ), .A2(_02326_ ), .A3(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A4(_06480_ ), .ZN(_06513_ ) );
AOI21_X1 _14359_ ( .A(_06513_ ), .B1(_06510_ ), .B2(\mylsu.araddr_tmp [15] ), .ZN(_06514_ ) );
BUF_X4 _14360_ ( .A(_02293_ ), .Z(_06515_ ) );
BUF_X4 _14361_ ( .A(_06515_ ), .Z(_06516_ ) );
OAI22_X1 _14362_ ( .A1(_06507_ ), .A2(_06514_ ), .B1(_02150_ ), .B2(_06516_ ), .ZN(\io_master_araddr [15] ) );
OAI221_X1 _14363_ ( .A(\IF_ID_pc [14] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02247_ ), .C2(_02248_ ), .ZN(_06517_ ) );
OR3_X1 _14364_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(_05678_ ), .ZN(_06518_ ) );
OAI211_X1 _14365_ ( .A(_02277_ ), .B(_06518_ ), .C1(\mylsu.araddr_tmp [14] ), .C2(_06509_ ), .ZN(_06519_ ) );
OAI21_X1 _14366_ ( .A(_06517_ ), .B1(\io_master_arburst [0] ), .B2(_06519_ ), .ZN(\io_master_araddr [14] ) );
NAND4_X1 _14367_ ( .A1(_02326_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_04950_ ), .A4(_06451_ ), .ZN(_06520_ ) );
OAI21_X1 _14368_ ( .A(_06520_ ), .B1(_06509_ ), .B2(\mylsu.araddr_tmp [5] ), .ZN(_06521_ ) );
OAI22_X1 _14369_ ( .A1(_06507_ ), .A2(_06521_ ), .B1(_06098_ ), .B2(_06516_ ), .ZN(\io_master_araddr [5] ) );
NAND4_X1 _14370_ ( .A1(_02326_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_04947_ ), .A4(_06480_ ), .ZN(_06522_ ) );
OAI21_X1 _14371_ ( .A(_06522_ ), .B1(_06509_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_06523_ ) );
OAI22_X1 _14372_ ( .A1(_06507_ ), .A2(_06523_ ), .B1(_06346_ ), .B2(_06516_ ), .ZN(\io_master_araddr [4] ) );
NOR2_X1 _14373_ ( .A1(_06509_ ), .A2(\mylsu.araddr_tmp [3] ), .ZN(_06524_ ) );
NOR3_X1 _14374_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(_05678_ ), .ZN(_06525_ ) );
NOR3_X1 _14375_ ( .A1(_02257_ ), .A2(_06524_ ), .A3(_06525_ ), .ZN(_06526_ ) );
BUF_X2 _14376_ ( .A(_02321_ ), .Z(_06527_ ) );
MUX2_X1 _14377_ ( .A(_06526_ ), .B(fanout_net_8 ), .S(_06527_ ), .Z(\io_master_araddr [3] ) );
OAI221_X1 _14378_ ( .A(\IF_ID_pc [13] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02247_ ), .C2(_02248_ ), .ZN(_06528_ ) );
OR3_X1 _14379_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(_05678_ ), .ZN(_06529_ ) );
OAI211_X1 _14380_ ( .A(_02277_ ), .B(_06529_ ), .C1(\mylsu.araddr_tmp [13] ), .C2(_06509_ ), .ZN(_06530_ ) );
OAI21_X1 _14381_ ( .A(_06528_ ), .B1(\io_master_arburst [0] ), .B2(_06530_ ), .ZN(\io_master_araddr [13] ) );
NOR2_X1 _14382_ ( .A1(_02274_ ), .A2(\mylsu.araddr_tmp [12] ), .ZN(_06531_ ) );
NOR3_X1 _14383_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(_02272_ ), .ZN(_06532_ ) );
NOR3_X1 _14384_ ( .A1(_02257_ ), .A2(_06531_ ), .A3(_06532_ ), .ZN(_06533_ ) );
MUX2_X1 _14385_ ( .A(_06533_ ), .B(\IF_ID_pc [12] ), .S(_06527_ ), .Z(\io_master_araddr [12] ) );
NOR3_X1 _14386_ ( .A1(_02290_ ), .A2(_06445_ ), .A3(_05678_ ), .ZN(_06534_ ) );
AOI21_X1 _14387_ ( .A(_06534_ ), .B1(_06510_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_06535_ ) );
OAI22_X1 _14388_ ( .A1(_06507_ ), .A2(_06535_ ), .B1(_05906_ ), .B2(_06516_ ), .ZN(\io_master_araddr [11] ) );
AND4_X1 _14389_ ( .A1(\EX_LS_dest_csreg_mem [10] ), .A2(_02326_ ), .A3(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A4(_06480_ ), .ZN(_06536_ ) );
AOI21_X1 _14390_ ( .A(_06536_ ), .B1(_06510_ ), .B2(\mylsu.araddr_tmp [10] ), .ZN(_06537_ ) );
OAI22_X1 _14391_ ( .A1(_06507_ ), .A2(_06537_ ), .B1(_02208_ ), .B2(_06516_ ), .ZN(\io_master_araddr [10] ) );
NAND4_X1 _14392_ ( .A1(_02326_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_04945_ ), .A4(_06480_ ), .ZN(_06538_ ) );
OAI21_X1 _14393_ ( .A(_06538_ ), .B1(_06509_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06539_ ) );
OAI22_X1 _14394_ ( .A1(_06507_ ), .A2(_06539_ ), .B1(_06119_ ), .B2(_06516_ ), .ZN(\io_master_araddr [9] ) );
NAND4_X1 _14395_ ( .A1(_02326_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_06468_ ), .A4(_06480_ ), .ZN(_06540_ ) );
OAI21_X1 _14396_ ( .A(_06540_ ), .B1(_06509_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_06541_ ) );
OAI22_X1 _14397_ ( .A1(_06507_ ), .A2(_06541_ ), .B1(_02233_ ), .B2(_06516_ ), .ZN(\io_master_araddr [8] ) );
NAND4_X1 _14398_ ( .A1(_02326_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_04954_ ), .A4(_06480_ ), .ZN(_06542_ ) );
OAI21_X1 _14399_ ( .A(_06542_ ), .B1(_06509_ ), .B2(\mylsu.araddr_tmp [7] ), .ZN(_06543_ ) );
OAI22_X1 _14400_ ( .A1(_06507_ ), .A2(_06543_ ), .B1(_02076_ ), .B2(_06516_ ), .ZN(\io_master_araddr [7] ) );
NOR2_X1 _14401_ ( .A1(_02274_ ), .A2(\mylsu.araddr_tmp [6] ), .ZN(_06544_ ) );
AOI211_X1 _14402_ ( .A(_02257_ ), .B(_06544_ ), .C1(_06471_ ), .C2(_06509_ ), .ZN(_06545_ ) );
MUX2_X1 _14403_ ( .A(_06545_ ), .B(\IF_ID_pc [6] ), .S(_06527_ ), .Z(\io_master_araddr [6] ) );
OR3_X1 _14404_ ( .A1(_02290_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(_02272_ ), .ZN(_06546_ ) );
OAI211_X1 _14405_ ( .A(_02277_ ), .B(_06546_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_02274_ ), .ZN(_06547_ ) );
NOR2_X1 _14406_ ( .A1(_02251_ ), .A2(_06547_ ), .ZN(_06548_ ) );
BUF_X4 _14407_ ( .A(_06548_ ), .Z(_06549_ ) );
BUF_X2 _14408_ ( .A(_06549_ ), .Z(\io_master_araddr [2] ) );
BUF_X2 _14409_ ( .A(_02270_ ), .Z(_06550_ ) );
BUF_X2 _14410_ ( .A(_06550_ ), .Z(\io_master_arid [1] ) );
NOR3_X1 _14411_ ( .A1(\io_master_arburst [0] ), .A2(_02332_ ), .A3(_02257_ ), .ZN(\io_master_arsize [2] ) );
NOR3_X1 _14412_ ( .A1(\io_master_arburst [0] ), .A2(_02331_ ), .A3(_02257_ ), .ZN(\io_master_arsize [0] ) );
INV_X1 _14413_ ( .A(\EX_LS_typ [2] ), .ZN(_06551_ ) );
OAI22_X1 _14414_ ( .A1(_02249_ ), .A2(_02250_ ), .B1(_06551_ ), .B2(_02257_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _14415_ ( .A(_02356_ ), .B(_02358_ ), .C1(_02296_ ), .C2(_02316_ ), .ZN(io_master_arvalid ) );
BUF_X2 _14416_ ( .A(_02346_ ), .Z(_06552_ ) );
AND2_X1 _14417_ ( .A1(_06552_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_06553_ ) );
BUF_X4 _14418_ ( .A(_06553_ ), .Z(_06554_ ) );
BUF_X4 _14419_ ( .A(_06554_ ), .Z(_06555_ ) );
MUX2_X1 _14420_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06555_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _14421_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06555_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _14422_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06555_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _14423_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06555_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _14424_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06555_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _14425_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06555_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _14426_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06555_ ), .Z(\io_master_awaddr [17] ) );
BUF_X4 _14427_ ( .A(_06554_ ), .Z(_06556_ ) );
MUX2_X1 _14428_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06556_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _14429_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06556_ ), .Z(\io_master_awaddr [15] ) );
MUX2_X1 _14430_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06556_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _14431_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06556_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _14432_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06556_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _14433_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06556_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _14434_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06556_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _14435_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06556_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _14436_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06556_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _14437_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06556_ ), .Z(\io_master_awaddr [8] ) );
BUF_X4 _14438_ ( .A(_06554_ ), .Z(_06557_ ) );
MUX2_X1 _14439_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06557_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _14440_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06557_ ), .Z(\io_master_awaddr [6] ) );
MUX2_X1 _14441_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06557_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _14442_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06557_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _14443_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06557_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _14444_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06557_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _14445_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06557_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _14446_ ( .A(\mylsu.awaddr_tmp [1] ), .B(\EX_LS_dest_csreg_mem [1] ), .S(_06557_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _14447_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_4 ), .S(_06557_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _14448_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06557_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _14449_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06554_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _14450_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06554_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _14451_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06554_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _14452_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06554_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _14453_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06554_ ), .Z(\io_master_awaddr [22] ) );
NAND4_X1 _14454_ ( .A1(_02351_ ), .A2(\EX_LS_typ [0] ), .A3(_06451_ ), .A4(_02335_ ), .ZN(\io_master_awsize [1] ) );
NOR2_X1 _14455_ ( .A1(\io_master_awsize [1] ), .A2(_02331_ ), .ZN(\io_master_awsize [0] ) );
NAND3_X1 _14456_ ( .A1(_02343_ ), .A2(_02354_ ), .A3(_06555_ ), .ZN(_06558_ ) );
INV_X1 _14457_ ( .A(\mylsu.state [4] ), .ZN(_06559_ ) );
NAND2_X1 _14458_ ( .A1(_06558_ ), .A2(_06559_ ), .ZN(io_master_awvalid ) );
INV_X1 _14459_ ( .A(\mylsu.state [2] ), .ZN(_06560_ ) );
INV_X1 _14460_ ( .A(\mylsu.state [1] ), .ZN(_06561_ ) );
NAND4_X1 _14461_ ( .A1(_06558_ ), .A2(_06560_ ), .A3(_06559_ ), .A4(_06561_ ), .ZN(io_master_bready ) );
NOR3_X1 _14462_ ( .A1(_02256_ ), .A2(\mylsu.state [0] ), .A3(\mylsu.state [1] ), .ZN(_06562_ ) );
NAND2_X1 _14463_ ( .A1(\io_master_bid [1] ), .A2(\io_master_bid [0] ), .ZN(_06563_ ) );
OR3_X1 _14464_ ( .A1(_06563_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bid [2] ), .ZN(_06564_ ) );
NOR2_X1 _14465_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_06565_ ) );
NAND2_X1 _14466_ ( .A1(_06565_ ), .A2(io_master_bvalid ), .ZN(_06566_ ) );
NOR2_X1 _14467_ ( .A1(_06564_ ), .A2(_06566_ ), .ZN(_06567_ ) );
NOR2_X1 _14468_ ( .A1(_06567_ ), .A2(_06561_ ), .ZN(_06568_ ) );
NOR3_X1 _14469_ ( .A1(_02366_ ), .A2(_02363_ ), .A3(_05676_ ), .ZN(_06569_ ) );
NOR2_X1 _14470_ ( .A1(_06419_ ), .A2(\io_master_rid [0] ), .ZN(_06570_ ) );
NAND4_X1 _14471_ ( .A1(_06570_ ), .A2(_06417_ ), .A3(_06418_ ), .A4(io_master_rlast ), .ZN(_06571_ ) );
NOR3_X1 _14472_ ( .A1(_02321_ ), .A2(_02257_ ), .A3(_06571_ ), .ZN(_06572_ ) );
OAI21_X1 _14473_ ( .A(_06414_ ), .B1(_06569_ ), .B2(_06572_ ), .ZN(_06573_ ) );
AOI211_X1 _14474_ ( .A(_06562_ ), .B(_06568_ ), .C1(_06573_ ), .C2(\mylsu.state [3] ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _14475_ ( .A(_02370_ ), .B(_02372_ ), .C1(_02296_ ), .C2(_02316_ ), .ZN(io_master_rready ) );
MUX2_X1 _14476_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_4 ), .Z(_06574_ ) );
INV_X1 _14477_ ( .A(\EX_LS_dest_csreg_mem [1] ), .ZN(_06575_ ) );
CLKBUF_X2 _14478_ ( .A(_06575_ ), .Z(_06576_ ) );
AND2_X1 _14479_ ( .A1(_06574_ ), .A2(_06576_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _14480_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_4 ), .Z(_06577_ ) );
AND2_X1 _14481_ ( .A1(_06577_ ), .A2(_06576_ ), .ZN(\io_master_wdata [14] ) );
INV_X1 _14482_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_06578_ ) );
NOR3_X1 _14483_ ( .A1(_06578_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _14484_ ( .A1(_05366_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [4] ) );
INV_X1 _14485_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_06579_ ) );
NOR3_X1 _14486_ ( .A1(_06579_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14487_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_06580_ ) );
NOR3_X1 _14488_ ( .A1(_06580_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14489_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06581_ ) );
NOR3_X1 _14490_ ( .A1(_06581_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14491_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06582_ ) );
NOR3_X1 _14492_ ( .A1(_06582_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14493_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_4 ), .Z(_06583_ ) );
AND2_X1 _14494_ ( .A1(_06583_ ), .A2(_06576_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14495_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_4 ), .Z(_06584_ ) );
AND2_X1 _14496_ ( .A1(_06584_ ), .A2(_06576_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14497_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_4 ), .Z(_06585_ ) );
AND2_X1 _14498_ ( .A1(_06585_ ), .A2(_06576_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14499_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_4 ), .Z(_06586_ ) );
AND2_X1 _14500_ ( .A1(_06586_ ), .A2(_06576_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14501_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_4 ), .Z(_06587_ ) );
AND2_X1 _14502_ ( .A1(_06587_ ), .A2(_06576_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14503_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_4 ), .Z(_06588_ ) );
AND2_X1 _14504_ ( .A1(_06588_ ), .A2(_06576_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14505_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06589_ ) );
NOR3_X1 _14506_ ( .A1(_06589_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [7] ) );
INV_X1 _14507_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_06590_ ) );
NOR3_X1 _14508_ ( .A1(_06590_ ), .A2(fanout_net_4 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14509_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_4 ), .Z(_06591_ ) );
MUX2_X1 _14510_ ( .A(_06591_ ), .B(_06574_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14511_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_4 ), .Z(_06592_ ) );
MUX2_X1 _14512_ ( .A(_06592_ ), .B(_06577_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [30] ) );
INV_X1 _14513_ ( .A(\EX_LS_result_csreg_mem [21] ), .ZN(_06593_ ) );
MUX2_X1 _14514_ ( .A(_06593_ ), .B(_05110_ ), .S(fanout_net_4 ), .Z(_06594_ ) );
NOR2_X1 _14515_ ( .A1(_06575_ ), .A2(fanout_net_4 ), .ZN(_06595_ ) );
INV_X1 _14516_ ( .A(_06595_ ), .ZN(_06596_ ) );
OAI22_X1 _14517_ ( .A1(_06594_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06596_ ), .B2(_06578_ ), .ZN(\io_master_wdata [21] ) );
OAI21_X1 _14518_ ( .A(_06575_ ), .B1(_06474_ ), .B2(\EX_LS_result_csreg_mem [12] ), .ZN(_06597_ ) );
NOR2_X1 _14519_ ( .A1(fanout_net_4 ), .A2(\EX_LS_result_csreg_mem [20] ), .ZN(_06598_ ) );
OAI22_X1 _14520_ ( .A1(_06596_ ), .A2(_05366_ ), .B1(_06597_ ), .B2(_06598_ ), .ZN(\io_master_wdata [20] ) );
OAI21_X1 _14521_ ( .A(_06575_ ), .B1(_06474_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_06599_ ) );
NOR2_X1 _14522_ ( .A1(fanout_net_4 ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_06600_ ) );
OAI22_X1 _14523_ ( .A1(_06596_ ), .A2(_06579_ ), .B1(_06599_ ), .B2(_06600_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _14524_ ( .A(_06575_ ), .B1(_06474_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_06601_ ) );
NOR2_X1 _14525_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_06602_ ) );
OAI22_X1 _14526_ ( .A1(_06596_ ), .A2(_06580_ ), .B1(_06601_ ), .B2(_06602_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _14527_ ( .A(_06575_ ), .B1(_06474_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_06603_ ) );
NOR2_X1 _14528_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_06604_ ) );
OAI22_X1 _14529_ ( .A1(_06596_ ), .A2(_06581_ ), .B1(_06603_ ), .B2(_06604_ ), .ZN(\io_master_wdata [17] ) );
INV_X1 _14530_ ( .A(\EX_LS_result_csreg_mem [16] ), .ZN(_06605_ ) );
INV_X1 _14531_ ( .A(\EX_LS_result_csreg_mem [8] ), .ZN(_06606_ ) );
MUX2_X1 _14532_ ( .A(_06605_ ), .B(_06606_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06607_ ) );
OAI22_X1 _14533_ ( .A1(_06607_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06596_ ), .B2(_06582_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14534_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06608_ ) );
MUX2_X1 _14535_ ( .A(_06608_ ), .B(_06583_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14536_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06609_ ) );
MUX2_X1 _14537_ ( .A(_06609_ ), .B(_06584_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14538_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06610_ ) );
MUX2_X1 _14539_ ( .A(_06610_ ), .B(_06585_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14540_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06611_ ) );
MUX2_X1 _14541_ ( .A(_06611_ ), .B(_06586_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14542_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06612_ ) );
MUX2_X1 _14543_ ( .A(_06612_ ), .B(_06587_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14544_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06613_ ) );
MUX2_X1 _14545_ ( .A(_06613_ ), .B(_06588_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [24] ) );
OAI21_X1 _14546_ ( .A(_06575_ ), .B1(_06474_ ), .B2(\EX_LS_result_csreg_mem [15] ), .ZN(_06614_ ) );
NOR2_X1 _14547_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [23] ), .ZN(_06615_ ) );
OAI22_X1 _14548_ ( .A1(_06596_ ), .A2(_06589_ ), .B1(_06614_ ), .B2(_06615_ ), .ZN(\io_master_wdata [23] ) );
OAI21_X1 _14549_ ( .A(_06575_ ), .B1(_06474_ ), .B2(\EX_LS_result_csreg_mem [14] ), .ZN(_06616_ ) );
NOR2_X1 _14550_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [22] ), .ZN(_06617_ ) );
OAI22_X1 _14551_ ( .A1(_06596_ ), .A2(_06590_ ), .B1(_06616_ ), .B2(_06617_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14552_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06618_ ) );
AND2_X1 _14553_ ( .A1(_06618_ ), .A2(_06576_ ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _14554_ ( .A1(_06474_ ), .A2(_06576_ ), .A3(\EX_LS_typ [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14555_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06619_ ) );
MUX2_X1 _14556_ ( .A(_06619_ ), .B(_06618_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14557_ ( .A1(_06575_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_06620_ ) );
NAND3_X1 _14558_ ( .A1(_06474_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_typ [0] ), .ZN(_06621_ ) );
OAI211_X1 _14559_ ( .A(_06620_ ), .B(_06621_ ), .C1(_02330_ ), .C2(_06551_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _14560_ ( .A1(_06558_ ), .A2(_06560_ ), .ZN(io_master_wvalid ) );
MUX2_X1 _14561_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14562_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14563_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14564_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
NOR2_X1 _14565_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06622_ ) );
AND2_X1 _14566_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06623_ ) );
NOR2_X1 _14567_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06624_ ) );
NOR2_X1 _14568_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06625_ ) );
AND4_X1 _14569_ ( .A1(_06622_ ), .A2(_06623_ ), .A3(_06624_ ), .A4(_06625_ ), .ZN(_06626_ ) );
AND2_X1 _14570_ ( .A1(_01773_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(_06627_ ) );
INV_X1 _14571_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_06628_ ) );
NOR3_X1 _14572_ ( .A1(_06628_ ), .A2(\LS_WB_waddr_csreg [3] ), .A3(\LS_WB_waddr_csreg [1] ), .ZN(_06629_ ) );
AND4_X1 _14573_ ( .A1(\LS_WB_waddr_csreg [2] ), .A2(_06626_ ), .A3(_06627_ ), .A4(_06629_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ) );
INV_X1 _14574_ ( .A(\LS_WB_waddr_csreg [7] ), .ZN(_06630_ ) );
AND3_X1 _14575_ ( .A1(_06622_ ), .A2(_06630_ ), .A3(\LS_WB_waddr_csreg [6] ), .ZN(_06631_ ) );
INV_X1 _14576_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_06632_ ) );
NOR2_X1 _14577_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_06633_ ) );
NAND4_X1 _14578_ ( .A1(_06631_ ), .A2(_06632_ ), .A3(\LS_WB_waddr_csreg [0] ), .A4(_06633_ ), .ZN(_06634_ ) );
NAND3_X1 _14579_ ( .A1(_06627_ ), .A2(_06625_ ), .A3(_06623_ ), .ZN(_06635_ ) );
NOR2_X1 _14580_ ( .A1(_06634_ ), .A2(_06635_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ) );
AND4_X1 _14581_ ( .A1(_06625_ ), .A2(_06631_ ), .A3(_06623_ ), .A4(_06633_ ), .ZN(_06636_ ) );
AND4_X1 _14582_ ( .A1(\LS_WB_waddr_csreg [1] ), .A2(_06636_ ), .A3(_06628_ ), .A4(_06627_ ), .ZN(_06637_ ) );
OR2_X1 _14583_ ( .A1(_06637_ ), .A2(_00093_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
AND2_X1 _14584_ ( .A1(_06622_ ), .A2(_06624_ ), .ZN(_06638_ ) );
NAND4_X1 _14585_ ( .A1(_06638_ ), .A2(_06632_ ), .A3(_06628_ ), .A4(_06633_ ), .ZN(_06639_ ) );
NOR2_X1 _14586_ ( .A1(_06639_ ), .A2(_06635_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _14587_ ( .A(_02355_ ), .ZN(_06640_ ) );
NOR2_X1 _14588_ ( .A1(_06481_ ), .A2(exception_quest_IDU ), .ZN(_06641_ ) );
NOR2_X1 _14589_ ( .A1(_06640_ ), .A2(_06641_ ), .ZN(_06642_ ) );
BUF_X4 _14590_ ( .A(_06642_ ), .Z(_06643_ ) );
MUX2_X1 _14591_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14592_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14593_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14594_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14595_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14596_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14597_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14598_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14599_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14600_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_06643_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14601_ ( .A(_06642_ ), .Z(_06644_ ) );
MUX2_X1 _14602_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14603_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14604_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14605_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14606_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14607_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14608_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14609_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14610_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14611_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_06644_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14612_ ( .A(_06642_ ), .Z(_06645_ ) );
MUX2_X1 _14613_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14614_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14615_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14616_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14617_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14618_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14619_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14620_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14621_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14622_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_06645_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14623_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_06642_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14624_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_06642_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
INV_X1 _14625_ ( .A(_02388_ ), .ZN(_06646_ ) );
NOR4_X1 _14626_ ( .A1(_06640_ ), .A2(exception_quest_IDU ), .A3(_06646_ ), .A4(_06641_ ), .ZN(_06647_ ) );
XNOR2_X1 _14627_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06648_ ) );
XNOR2_X1 _14628_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06649_ ) );
XNOR2_X1 _14629_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06650_ ) );
XNOR2_X1 _14630_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06651_ ) );
NAND4_X1 _14631_ ( .A1(_06648_ ), .A2(_06649_ ), .A3(_06650_ ), .A4(_06651_ ), .ZN(_06652_ ) );
XNOR2_X1 _14632_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06653_ ) );
XNOR2_X1 _14633_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06654_ ) );
NAND2_X1 _14634_ ( .A1(_06653_ ), .A2(_06654_ ), .ZN(_06655_ ) );
XOR2_X1 _14635_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .Z(_06656_ ) );
XOR2_X1 _14636_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .Z(_06657_ ) );
NOR4_X1 _14637_ ( .A1(_06652_ ), .A2(_06655_ ), .A3(_06656_ ), .A4(_06657_ ), .ZN(_06658_ ) );
XNOR2_X1 _14638_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_06659_ ) );
XNOR2_X1 _14639_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_06660_ ) );
XNOR2_X1 _14640_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_06661_ ) );
XNOR2_X1 _14641_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_06662_ ) );
AND4_X1 _14642_ ( .A1(_06659_ ), .A2(_06660_ ), .A3(_06661_ ), .A4(_06662_ ), .ZN(_06663_ ) );
XNOR2_X1 _14643_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06664_ ) );
XNOR2_X1 _14644_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06665_ ) );
XNOR2_X1 _14645_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06666_ ) );
XNOR2_X1 _14646_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06667_ ) );
AND4_X1 _14647_ ( .A1(_06664_ ), .A2(_06665_ ), .A3(_06666_ ), .A4(_06667_ ), .ZN(_06668_ ) );
AND3_X1 _14648_ ( .A1(_06658_ ), .A2(_06663_ ), .A3(_06668_ ), .ZN(_06669_ ) );
XNOR2_X1 _14649_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06670_ ) );
XNOR2_X1 _14650_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06671_ ) );
XNOR2_X1 _14651_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06672_ ) );
XNOR2_X1 _14652_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06673_ ) );
NAND4_X1 _14653_ ( .A1(_06670_ ), .A2(_06671_ ), .A3(_06672_ ), .A4(_06673_ ), .ZN(_06674_ ) );
XNOR2_X1 _14654_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06675_ ) );
XNOR2_X1 _14655_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06676_ ) );
NAND2_X1 _14656_ ( .A1(_06675_ ), .A2(_06676_ ), .ZN(_06677_ ) );
XOR2_X1 _14657_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .Z(_06678_ ) );
XOR2_X1 _14658_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .Z(_06679_ ) );
NOR4_X1 _14659_ ( .A1(_06674_ ), .A2(_06677_ ), .A3(_06678_ ), .A4(_06679_ ), .ZN(_06680_ ) );
XNOR2_X1 _14660_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06681_ ) );
XNOR2_X1 _14661_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06682_ ) );
XNOR2_X1 _14662_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06683_ ) );
XNOR2_X1 _14663_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06684_ ) );
AND4_X1 _14664_ ( .A1(_06681_ ), .A2(_06682_ ), .A3(_06683_ ), .A4(_06684_ ), .ZN(_06685_ ) );
XNOR2_X1 _14665_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06686_ ) );
XNOR2_X1 _14666_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06687_ ) );
XNOR2_X1 _14667_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06688_ ) );
XNOR2_X1 _14668_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06689_ ) );
AND4_X1 _14669_ ( .A1(_06686_ ), .A2(_06687_ ), .A3(_06688_ ), .A4(_06689_ ), .ZN(_06690_ ) );
AND3_X1 _14670_ ( .A1(_06680_ ), .A2(_06685_ ), .A3(_06690_ ), .ZN(_06691_ ) );
NAND3_X1 _14671_ ( .A1(_06669_ ), .A2(_06691_ ), .A3(excp_written ), .ZN(_06692_ ) );
AOI21_X1 _14672_ ( .A(_06647_ ), .B1(_06646_ ), .B2(_06692_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14673_ ( .A(_03341_ ), .ZN(_06693_ ) );
BUF_X4 _14674_ ( .A(_06693_ ), .Z(_06694_ ) );
BUF_X4 _14675_ ( .A(_06694_ ), .Z(_06695_ ) );
OAI22_X1 _14676_ ( .A1(_05448_ ), .A2(_03382_ ), .B1(_03563_ ), .B2(_06695_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _14677_ ( .A(_04058_ ), .B(\ID_EX_imm [0] ), .ZN(_06696_ ) );
BUF_X4 _14678_ ( .A(_03341_ ), .Z(_06697_ ) );
BUF_X4 _14679_ ( .A(_06697_ ), .Z(_06698_ ) );
AOI22_X1 _14680_ ( .A1(_06696_ ), .A2(_03344_ ), .B1(_03547_ ), .B2(_06698_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
NOR3_X1 _14681_ ( .A1(_05223_ ), .A2(_05173_ ), .A3(_03343_ ), .ZN(_06699_ ) );
BUF_X2 _14682_ ( .A(_06693_ ), .Z(_06700_ ) );
MUX2_X1 _14683_ ( .A(\ID_EX_csr [10] ), .B(_06699_ ), .S(_06700_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
INV_X2 _14684_ ( .A(_03343_ ), .ZN(_06701_ ) );
BUF_X4 _14685_ ( .A(_06701_ ), .Z(_06702_ ) );
NAND2_X1 _14686_ ( .A1(_05249_ ), .A2(_06702_ ), .ZN(_06703_ ) );
MUX2_X1 _14687_ ( .A(\ID_EX_csr [9] ), .B(_06703_ ), .S(_06700_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
NOR4_X1 _14688_ ( .A1(_05672_ ), .A2(_04920_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [8] ), .ZN(_06704_ ) );
AOI21_X1 _14689_ ( .A(_06704_ ), .B1(_05273_ ), .B2(_03344_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
OAI22_X1 _14690_ ( .A1(_05303_ ), .A2(_03382_ ), .B1(_04956_ ), .B2(_06695_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
BUF_X4 _14691_ ( .A(_03341_ ), .Z(_06705_ ) );
BUF_X4 _14692_ ( .A(_06705_ ), .Z(_06706_ ) );
AOI22_X1 _14693_ ( .A1(_05327_ ), .A2(_03344_ ), .B1(_03553_ ), .B2(_06706_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14694_ ( .A1(_05354_ ), .A2(_03344_ ), .ZN(_06707_ ) );
OAI21_X1 _14695_ ( .A(_06707_ ), .B1(_03544_ ), .B2(_06695_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
OAI22_X1 _14696_ ( .A1(_05377_ ), .A2(_03345_ ), .B1(_04937_ ), .B2(_06695_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND3_X1 _14697_ ( .A1(_05406_ ), .A2(_03344_ ), .A3(_02809_ ), .ZN(_06708_ ) );
OAI21_X1 _14698_ ( .A(_06708_ ), .B1(_03567_ ), .B2(_06695_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _14699_ ( .A1(_05428_ ), .A2(_02807_ ), .A3(_03343_ ), .ZN(_06709_ ) );
MUX2_X1 _14700_ ( .A(\ID_EX_csr [2] ), .B(_06709_ ), .S(_06700_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
NAND4_X1 _14701_ ( .A1(_02412_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_csr [11] ), .ZN(_06710_ ) );
OAI21_X1 _14702_ ( .A(_06710_ ), .B1(_05175_ ), .B2(_03382_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X4 _14703_ ( .A(_06705_ ), .Z(_06711_ ) );
NAND4_X1 _14704_ ( .A1(_05190_ ), .A2(_05055_ ), .A3(_05056_ ), .A4(\mycsreg.CSReg[0][21] ), .ZN(_06712_ ) );
NAND2_X1 _14705_ ( .A1(_05627_ ), .A2(_06712_ ), .ZN(_06713_ ) );
NOR2_X1 _14706_ ( .A1(_05390_ ), .A2(_06713_ ), .ZN(_06714_ ) );
INV_X1 _14707_ ( .A(_05013_ ), .ZN(_06715_ ) );
BUF_X2 _14708_ ( .A(_05015_ ), .Z(_06716_ ) );
BUF_X2 _14709_ ( .A(_04838_ ), .Z(_06717_ ) );
NAND3_X1 _14710_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_06717_ ), .ZN(_06718_ ) );
NAND2_X1 _14711_ ( .A1(_04904_ ), .A2(\mtvec [21] ), .ZN(_06719_ ) );
NAND4_X1 _14712_ ( .A1(_06714_ ), .A2(_06715_ ), .A3(_06718_ ), .A4(_06719_ ), .ZN(_06720_ ) );
OR3_X1 _14713_ ( .A1(_05022_ ), .A2(\EX_LS_result_csreg_mem [21] ), .A3(_04913_ ), .ZN(_06721_ ) );
NAND2_X1 _14714_ ( .A1(_06720_ ), .A2(_06721_ ), .ZN(_06722_ ) );
AOI22_X1 _14715_ ( .A1(_06722_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02576_ ), .ZN(_06723_ ) );
NAND3_X1 _14716_ ( .A1(_02551_ ), .A2(_05305_ ), .A3(_02573_ ), .ZN(_06724_ ) );
AND2_X1 _14717_ ( .A1(_06723_ ), .A2(_06724_ ), .ZN(_06725_ ) );
NOR2_X1 _14718_ ( .A1(_04417_ ), .A2(\ID_EX_typ [2] ), .ZN(_06726_ ) );
BUF_X2 _14719_ ( .A(_06726_ ), .Z(_06727_ ) );
AND3_X1 _14720_ ( .A1(_06720_ ), .A2(_06727_ ), .A3(_06721_ ), .ZN(_06728_ ) );
OAI21_X1 _14721_ ( .A(_06711_ ), .B1(_06725_ ), .B2(_06728_ ), .ZN(_06729_ ) );
BUF_X4 _14722_ ( .A(_06697_ ), .Z(_06730_ ) );
BUF_X4 _14723_ ( .A(_06701_ ), .Z(_06731_ ) );
MUX2_X1 _14724_ ( .A(_05623_ ), .B(_03791_ ), .S(_06731_ ), .Z(_06732_ ) );
OAI21_X1 _14725_ ( .A(_06729_ ), .B1(_06730_ ), .B2(_06732_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
NOR3_X1 _14726_ ( .A1(_04901_ ), .A2(_06246_ ), .A3(_04902_ ), .ZN(_06733_ ) );
NOR2_X1 _14727_ ( .A1(_05390_ ), .A2(_06733_ ), .ZN(_06734_ ) );
NAND3_X1 _14728_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_06717_ ), .ZN(_06735_ ) );
NAND4_X1 _14729_ ( .A1(_04942_ ), .A2(_05076_ ), .A3(_05056_ ), .A4(\mycsreg.CSReg[0][20] ), .ZN(_06736_ ) );
AND2_X1 _14730_ ( .A1(_04834_ ), .A2(_06736_ ), .ZN(_06737_ ) );
NAND4_X1 _14731_ ( .A1(_06734_ ), .A2(_06735_ ), .A3(_05014_ ), .A4(_06737_ ), .ZN(_06738_ ) );
OR3_X1 _14732_ ( .A1(_05022_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_04913_ ), .ZN(_06739_ ) );
AND2_X1 _14733_ ( .A1(_06738_ ), .A2(_06739_ ), .ZN(_06740_ ) );
OAI22_X1 _14734_ ( .A1(_06740_ ), .A2(_05686_ ), .B1(_03516_ ), .B2(\ID_EX_imm [20] ), .ZN(_06741_ ) );
INV_X1 _14735_ ( .A(_02598_ ), .ZN(_06742_ ) );
AOI21_X1 _14736_ ( .A(_06741_ ), .B1(_05687_ ), .B2(_06742_ ), .ZN(_06743_ ) );
BUF_X4 _14737_ ( .A(_06726_ ), .Z(_06744_ ) );
NAND3_X1 _14738_ ( .A1(_06738_ ), .A2(_06744_ ), .A3(_06739_ ), .ZN(_06745_ ) );
INV_X1 _14739_ ( .A(_06745_ ), .ZN(_06746_ ) );
OAI21_X1 _14740_ ( .A(_06711_ ), .B1(_06743_ ), .B2(_06746_ ), .ZN(_06747_ ) );
MUX2_X1 _14741_ ( .A(_05621_ ), .B(_03769_ ), .S(_06731_ ), .Z(_06748_ ) );
OAI21_X1 _14742_ ( .A(_06747_ ), .B1(_06730_ ), .B2(_06748_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
AOI22_X1 _14743_ ( .A1(_04916_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02656_ ), .ZN(_06749_ ) );
BUF_X4 _14744_ ( .A(_03341_ ), .Z(_06750_ ) );
OAI211_X1 _14745_ ( .A(_06749_ ), .B(_06750_ ), .C1(fanout_net_5 ), .C2(_02655_ ), .ZN(_06751_ ) );
INV_X1 _14746_ ( .A(_06726_ ), .ZN(_06752_ ) );
OR3_X1 _14747_ ( .A1(_04916_ ), .A2(_06694_ ), .A3(_06752_ ), .ZN(_06753_ ) );
BUF_X4 _14748_ ( .A(_06701_ ), .Z(_06754_ ) );
MUX2_X1 _14749_ ( .A(_05666_ ), .B(_03655_ ), .S(_06754_ ), .Z(_06755_ ) );
OAI211_X1 _14750_ ( .A(_06751_ ), .B(_06753_ ), .C1(_06730_ ), .C2(_06755_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
AOI22_X1 _14751_ ( .A1(_04962_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02627_ ), .ZN(_06756_ ) );
OAI21_X1 _14752_ ( .A(_06756_ ), .B1(fanout_net_5 ), .B2(_02626_ ), .ZN(_06757_ ) );
OAI21_X1 _14753_ ( .A(_06744_ ), .B1(_04960_ ), .B2(_04961_ ), .ZN(_06758_ ) );
AOI21_X1 _14754_ ( .A(_06694_ ), .B1(_06757_ ), .B2(_06758_ ), .ZN(_06759_ ) );
AND3_X1 _14755_ ( .A1(_03342_ ), .A2(_05667_ ), .A3(\ID_EX_typ [7] ), .ZN(_06760_ ) );
AOI211_X1 _14756_ ( .A(_06705_ ), .B(_06760_ ), .C1(_03692_ ), .C2(_06702_ ), .ZN(_06761_ ) );
OR2_X1 _14757_ ( .A1(_06759_ ), .A2(_06761_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
NOR2_X1 _14758_ ( .A1(_06754_ ), .A2(\ID_EX_pc [17] ), .ZN(_06762_ ) );
AOI21_X1 _14759_ ( .A(_06762_ ), .B1(_03721_ ), .B2(_06731_ ), .ZN(_06763_ ) );
NAND4_X1 _14760_ ( .A1(_03573_ ), .A2(_03560_ ), .A3(_03574_ ), .A4(\mycsreg.CSReg[0][17] ), .ZN(_06764_ ) );
NAND2_X1 _14761_ ( .A1(_04983_ ), .A2(_06764_ ), .ZN(_06765_ ) );
NOR2_X1 _14762_ ( .A1(_05390_ ), .A2(_06765_ ), .ZN(_06766_ ) );
NAND3_X1 _14763_ ( .A1(_05015_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_04838_ ), .ZN(_06767_ ) );
NAND2_X1 _14764_ ( .A1(_04903_ ), .A2(\mtvec [17] ), .ZN(_06768_ ) );
AND4_X1 _14765_ ( .A1(_05014_ ), .A2(_06766_ ), .A3(_06767_ ), .A4(_06768_ ), .ZN(_06769_ ) );
NOR3_X1 _14766_ ( .A1(_05022_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_04913_ ), .ZN(_06770_ ) );
NOR2_X1 _14767_ ( .A1(_06769_ ), .A2(_06770_ ), .ZN(_06771_ ) );
OAI22_X1 _14768_ ( .A1(_06771_ ), .A2(_04771_ ), .B1(_02419_ ), .B2(\ID_EX_imm [17] ), .ZN(_06772_ ) );
AOI21_X1 _14769_ ( .A(_06772_ ), .B1(_05305_ ), .B2(_03695_ ), .ZN(_06773_ ) );
OR3_X1 _14770_ ( .A1(_06769_ ), .A2(_06752_ ), .A3(_06770_ ), .ZN(_06774_ ) );
INV_X1 _14771_ ( .A(_06774_ ), .ZN(_06775_ ) );
OR2_X1 _14772_ ( .A1(_06773_ ), .A2(_06775_ ), .ZN(_06776_ ) );
MUX2_X1 _14773_ ( .A(_06763_ ), .B(_06776_ ), .S(_06697_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
OAI22_X1 _14774_ ( .A1(_05026_ ), .A2(_05686_ ), .B1(_03516_ ), .B2(\ID_EX_imm [16] ), .ZN(_06777_ ) );
AOI21_X1 _14775_ ( .A(_06777_ ), .B1(_05687_ ), .B2(_04572_ ), .ZN(_06778_ ) );
INV_X1 _14776_ ( .A(_05025_ ), .ZN(_06779_ ) );
OAI211_X1 _14777_ ( .A(_06779_ ), .B(_06727_ ), .C1(_05020_ ), .C2(_05023_ ), .ZN(_06780_ ) );
INV_X1 _14778_ ( .A(_06780_ ), .ZN(_06781_ ) );
OAI21_X1 _14779_ ( .A(_06711_ ), .B1(_06778_ ), .B2(_06781_ ), .ZN(_06782_ ) );
MUX2_X1 _14780_ ( .A(_04974_ ), .B(_03746_ ), .S(_06731_ ), .Z(_06783_ ) );
OAI21_X1 _14781_ ( .A(_06782_ ), .B1(_06730_ ), .B2(_06783_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
AOI21_X1 _14782_ ( .A(fanout_net_5 ), .B1(_03074_ ), .B2(_03093_ ), .ZN(_06784_ ) );
AND2_X1 _14783_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [15] ), .ZN(_06785_ ) );
NAND3_X1 _14784_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(\EX_LS_result_csreg_mem [15] ), .ZN(_06786_ ) );
BUF_X4 _14785_ ( .A(_05278_ ), .Z(_06787_ ) );
NAND3_X1 _14786_ ( .A1(_06787_ ), .A2(\mtvec [15] ), .A3(_04987_ ), .ZN(_06788_ ) );
NAND3_X1 _14787_ ( .A1(_05278_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_05059_ ), .ZN(_06789_ ) );
NAND2_X1 _14788_ ( .A1(_06788_ ), .A2(_06789_ ), .ZN(_06790_ ) );
AND4_X1 _14789_ ( .A1(\mycsreg.CSReg[3][15] ), .A2(_06717_ ), .A3(_04897_ ), .A4(_04845_ ), .ZN(_06791_ ) );
AND4_X1 _14790_ ( .A1(\mepc [15] ), .A2(_05456_ ), .A3(_06717_ ), .A4(_04845_ ), .ZN(_06792_ ) );
NOR4_X1 _14791_ ( .A1(_06790_ ), .A2(_04893_ ), .A3(_06791_ ), .A4(_06792_ ), .ZN(_06793_ ) );
OAI21_X1 _14792_ ( .A(_06786_ ), .B1(_06793_ ), .B2(_05103_ ), .ZN(_06794_ ) );
OAI221_X1 _14793_ ( .A(_06697_ ), .B1(_06784_ ), .B2(_06785_ ), .C1(_05686_ ), .C2(_06794_ ), .ZN(_06795_ ) );
INV_X1 _14794_ ( .A(_05390_ ), .ZN(_06796_ ) );
AOI21_X1 _14795_ ( .A(_06791_ ), .B1(_04892_ ), .B2(_04897_ ), .ZN(_06797_ ) );
NAND2_X1 _14796_ ( .A1(_04904_ ), .A2(\mtvec [15] ), .ZN(_06798_ ) );
NAND4_X1 _14797_ ( .A1(_04991_ ), .A2(_04992_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][15] ), .ZN(_06799_ ) );
AND2_X1 _14798_ ( .A1(_05050_ ), .A2(_06799_ ), .ZN(_06800_ ) );
NAND4_X1 _14799_ ( .A1(_06796_ ), .A2(_06797_ ), .A3(_06798_ ), .A4(_06800_ ), .ZN(_06801_ ) );
BUF_X4 _14800_ ( .A(_03341_ ), .Z(_06802_ ) );
OR3_X1 _14801_ ( .A1(_05583_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_04914_ ), .ZN(_06803_ ) );
NAND4_X1 _14802_ ( .A1(_06801_ ), .A2(_06802_ ), .A3(_06744_ ), .A4(_06803_ ), .ZN(_06804_ ) );
MUX2_X1 _14803_ ( .A(_05037_ ), .B(_04153_ ), .S(_06731_ ), .Z(_06805_ ) );
OAI211_X1 _14804_ ( .A(_06795_ ), .B(_06804_ ), .C1(_06805_ ), .C2(_06698_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
AND2_X1 _14805_ ( .A1(_04903_ ), .A2(\mtvec [14] ), .ZN(_06806_ ) );
NOR2_X1 _14806_ ( .A1(_05390_ ), .A2(_06806_ ), .ZN(_06807_ ) );
NAND3_X1 _14807_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_06717_ ), .ZN(_06808_ ) );
NAND4_X1 _14808_ ( .A1(_04842_ ), .A2(_04833_ ), .A3(_04846_ ), .A4(\mycsreg.CSReg[0][14] ), .ZN(_06809_ ) );
AND2_X1 _14809_ ( .A1(_05077_ ), .A2(_06809_ ), .ZN(_06810_ ) );
AND4_X1 _14810_ ( .A1(_05014_ ), .A2(_06807_ ), .A3(_06808_ ), .A4(_06810_ ), .ZN(_06811_ ) );
NOR3_X1 _14811_ ( .A1(_04912_ ), .A2(\EX_LS_result_csreg_mem [14] ), .A3(_05216_ ), .ZN(_06812_ ) );
NOR2_X1 _14812_ ( .A1(_06811_ ), .A2(_06812_ ), .ZN(_06813_ ) );
OAI22_X1 _14813_ ( .A1(_06813_ ), .A2(_05686_ ), .B1(_03516_ ), .B2(\ID_EX_imm [14] ), .ZN(_06814_ ) );
AOI21_X1 _14814_ ( .A(_06814_ ), .B1(_05687_ ), .B2(_04685_ ), .ZN(_06815_ ) );
OR3_X1 _14815_ ( .A1(_06811_ ), .A2(_06752_ ), .A3(_06812_ ), .ZN(_06816_ ) );
INV_X1 _14816_ ( .A(_06816_ ), .ZN(_06817_ ) );
OAI21_X1 _14817_ ( .A(_06711_ ), .B1(_06815_ ), .B2(_06817_ ), .ZN(_06818_ ) );
MUX2_X1 _14818_ ( .A(_05035_ ), .B(_04176_ ), .S(_06731_ ), .Z(_06819_ ) );
OAI21_X1 _14819_ ( .A(_06818_ ), .B1(_06730_ ), .B2(_06819_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
INV_X1 _14820_ ( .A(_05111_ ), .ZN(_06820_ ) );
NOR2_X1 _14821_ ( .A1(_05103_ ), .A2(_05013_ ), .ZN(_06821_ ) );
INV_X1 _14822_ ( .A(_06821_ ), .ZN(_06822_ ) );
OAI211_X1 _14823_ ( .A(_06726_ ), .B(_06820_ ), .C1(_06822_ ), .C2(_05108_ ), .ZN(_06823_ ) );
INV_X1 _14824_ ( .A(_06823_ ), .ZN(_06824_ ) );
AOI22_X1 _14825_ ( .A1(_05113_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_03045_ ), .ZN(_06825_ ) );
NAND3_X1 _14826_ ( .A1(_03044_ ), .A2(_05305_ ), .A3(_03046_ ), .ZN(_06826_ ) );
AOI21_X1 _14827_ ( .A(_06824_ ), .B1(_06825_ ), .B2(_06826_ ), .ZN(_06827_ ) );
NOR2_X1 _14828_ ( .A1(_06827_ ), .A2(_06700_ ), .ZN(_06828_ ) );
NOR2_X1 _14829_ ( .A1(_06754_ ), .A2(\ID_EX_pc [13] ), .ZN(_06829_ ) );
AOI211_X1 _14830_ ( .A(_06705_ ), .B(_06829_ ), .C1(_04200_ ), .C2(_06702_ ), .ZN(_06830_ ) );
OR2_X1 _14831_ ( .A1(_06828_ ), .A2(_06830_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
NAND4_X1 _14832_ ( .A1(_04942_ ), .A2(_05076_ ), .A3(_04846_ ), .A4(\mycsreg.CSReg[0][12] ), .ZN(_06831_ ) );
NAND2_X1 _14833_ ( .A1(_05124_ ), .A2(_06831_ ), .ZN(_06832_ ) );
NOR2_X1 _14834_ ( .A1(_05390_ ), .A2(_06832_ ), .ZN(_06833_ ) );
NAND3_X1 _14835_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_06717_ ), .ZN(_06834_ ) );
OR3_X1 _14836_ ( .A1(_04901_ ), .A2(_06287_ ), .A3(_04902_ ), .ZN(_06835_ ) );
NAND4_X1 _14837_ ( .A1(_06833_ ), .A2(_05014_ ), .A3(_06834_ ), .A4(_06835_ ), .ZN(_06836_ ) );
OR3_X1 _14838_ ( .A1(_05022_ ), .A2(\EX_LS_result_csreg_mem [12] ), .A3(_04913_ ), .ZN(_06837_ ) );
AND2_X1 _14839_ ( .A1(_06836_ ), .A2(_06837_ ), .ZN(_06838_ ) );
OAI22_X1 _14840_ ( .A1(_06838_ ), .A2(_05686_ ), .B1(_03516_ ), .B2(\ID_EX_imm [12] ), .ZN(_06839_ ) );
INV_X1 _14841_ ( .A(_03070_ ), .ZN(_06840_ ) );
AOI21_X1 _14842_ ( .A(_06839_ ), .B1(_05687_ ), .B2(_06840_ ), .ZN(_06841_ ) );
NAND3_X1 _14843_ ( .A1(_06836_ ), .A2(_06727_ ), .A3(_06837_ ), .ZN(_06842_ ) );
INV_X1 _14844_ ( .A(_06842_ ), .ZN(_06843_ ) );
OAI21_X1 _14845_ ( .A(_06711_ ), .B1(_06841_ ), .B2(_06843_ ), .ZN(_06844_ ) );
MUX2_X1 _14846_ ( .A(_05095_ ), .B(_04222_ ), .S(_06754_ ), .Z(_06845_ ) );
OAI21_X1 _14847_ ( .A(_06844_ ), .B1(_06730_ ), .B2(_06845_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
NAND2_X1 _14848_ ( .A1(_04903_ ), .A2(\mtvec [30] ), .ZN(_06846_ ) );
OAI21_X1 _14849_ ( .A(_06846_ ), .B1(_05022_ ), .B2(_04913_ ), .ZN(_06847_ ) );
AND3_X1 _14850_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_05210_ ), .ZN(_06848_ ) );
NAND4_X1 _14851_ ( .A1(_04942_ ), .A2(_05076_ ), .A3(_05056_ ), .A4(\mycsreg.CSReg[0][30] ), .ZN(_06849_ ) );
NAND2_X1 _14852_ ( .A1(_03561_ ), .A2(_06849_ ), .ZN(_06850_ ) );
NOR4_X1 _14853_ ( .A1(_06847_ ), .A2(_05013_ ), .A3(_06848_ ), .A4(_06850_ ), .ZN(_06851_ ) );
NOR3_X1 _14854_ ( .A1(_04912_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_05216_ ), .ZN(_06852_ ) );
NOR2_X1 _14855_ ( .A1(_06851_ ), .A2(_06852_ ), .ZN(_06853_ ) );
OAI22_X1 _14856_ ( .A1(_06853_ ), .A2(_04771_ ), .B1(_03516_ ), .B2(\ID_EX_imm [30] ), .ZN(_06854_ ) );
AOI21_X1 _14857_ ( .A(_06854_ ), .B1(_03310_ ), .B2(_04785_ ), .ZN(_06855_ ) );
OR3_X1 _14858_ ( .A1(_06851_ ), .A2(_06752_ ), .A3(_06852_ ), .ZN(_06856_ ) );
INV_X1 _14859_ ( .A(_06856_ ), .ZN(_06857_ ) );
OAI21_X1 _14860_ ( .A(_06711_ ), .B1(_06855_ ), .B2(_06857_ ), .ZN(_06858_ ) );
MUX2_X1 _14861_ ( .A(_03599_ ), .B(_03938_ ), .S(_06754_ ), .Z(_06859_ ) );
OAI21_X1 _14862_ ( .A(_06858_ ), .B1(_06730_ ), .B2(_06859_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _14863_ ( .A1(_04939_ ), .A2(\mtvec [11] ), .A3(_04940_ ), .ZN(_06860_ ) );
NAND3_X1 _14864_ ( .A1(_04939_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_04942_ ), .ZN(_06861_ ) );
NAND3_X1 _14865_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_05210_ ), .ZN(_06862_ ) );
NAND4_X1 _14866_ ( .A1(_04934_ ), .A2(_04838_ ), .A3(\mepc [11] ), .A4(_04844_ ), .ZN(_06863_ ) );
NAND4_X1 _14867_ ( .A1(_06860_ ), .A2(_06861_ ), .A3(_06862_ ), .A4(_06863_ ), .ZN(_06864_ ) );
NOR4_X1 _14868_ ( .A1(_05103_ ), .A2(_06864_ ), .A3(_05013_ ), .A4(_04893_ ), .ZN(_06865_ ) );
INV_X1 _14869_ ( .A(\EX_LS_result_csreg_mem [11] ), .ZN(_06866_ ) );
AND3_X1 _14870_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_06866_ ), .ZN(_06867_ ) );
NOR2_X1 _14871_ ( .A1(_06865_ ), .A2(_06867_ ), .ZN(_06868_ ) );
OAI22_X1 _14872_ ( .A1(_06868_ ), .A2(_04771_ ), .B1(_03516_ ), .B2(\ID_EX_imm [11] ), .ZN(_06869_ ) );
AOI21_X1 _14873_ ( .A(_06869_ ), .B1(_05687_ ), .B2(_04249_ ), .ZN(_06870_ ) );
NOR3_X1 _14874_ ( .A1(_06865_ ), .A2(_06752_ ), .A3(_06867_ ), .ZN(_06871_ ) );
OAI21_X1 _14875_ ( .A(_06711_ ), .B1(_06870_ ), .B2(_06871_ ), .ZN(_06872_ ) );
MUX2_X1 _14876_ ( .A(_05149_ ), .B(_04247_ ), .S(_06754_ ), .Z(_06873_ ) );
OAI21_X1 _14877_ ( .A(_06872_ ), .B1(_06730_ ), .B2(_06873_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _14878_ ( .A(fanout_net_5 ), .B1(_02992_ ), .B2(_03011_ ), .ZN(_06874_ ) );
AND2_X1 _14879_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [10] ), .ZN(_06875_ ) );
NOR2_X1 _14880_ ( .A1(_05215_ ), .A2(_05217_ ), .ZN(_06876_ ) );
OAI221_X1 _14881_ ( .A(_06697_ ), .B1(_06874_ ), .B2(_06875_ ), .C1(_06876_ ), .C2(_05686_ ), .ZN(_06877_ ) );
NAND3_X1 _14882_ ( .A1(_06876_ ), .A2(_06802_ ), .A3(_06744_ ), .ZN(_06878_ ) );
MUX2_X1 _14883_ ( .A(_05202_ ), .B(_04271_ ), .S(_06754_ ), .Z(_06879_ ) );
OAI211_X1 _14884_ ( .A(_06877_ ), .B(_06878_ ), .C1(_06730_ ), .C2(_06879_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
AND4_X1 _14885_ ( .A1(\mycsreg.CSReg[3][9] ), .A2(_03562_ ), .A3(_03565_ ), .A4(_04800_ ), .ZN(_06880_ ) );
AND4_X1 _14886_ ( .A1(\mepc [9] ), .A2(_04933_ ), .A3(_04798_ ), .A4(_04800_ ), .ZN(_06881_ ) );
AOI211_X1 _14887_ ( .A(_06880_ ), .B(_06881_ ), .C1(_04892_ ), .C2(_04897_ ), .ZN(_06882_ ) );
NAND3_X1 _14888_ ( .A1(_04939_ ), .A2(\mtvec [9] ), .A3(_04940_ ), .ZN(_06883_ ) );
NAND3_X1 _14889_ ( .A1(_04939_ ), .A2(\mycsreg.CSReg[0][9] ), .A3(_04842_ ), .ZN(_06884_ ) );
AND2_X1 _14890_ ( .A1(_06883_ ), .A2(_06884_ ), .ZN(_06885_ ) );
AOI21_X1 _14891_ ( .A(_05103_ ), .B1(_06882_ ), .B2(_06885_ ), .ZN(_06886_ ) );
AND3_X1 _14892_ ( .A1(_04953_ ), .A2(_04959_ ), .A3(\EX_LS_result_csreg_mem [9] ), .ZN(_06887_ ) );
NOR2_X1 _14893_ ( .A1(_06886_ ), .A2(_06887_ ), .ZN(_06888_ ) );
AOI22_X1 _14894_ ( .A1(_06888_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02964_ ), .ZN(_06889_ ) );
OAI21_X1 _14895_ ( .A(_06889_ ), .B1(fanout_net_5 ), .B2(_02963_ ), .ZN(_06890_ ) );
OAI21_X1 _14896_ ( .A(_06727_ ), .B1(_06886_ ), .B2(_06887_ ), .ZN(_06891_ ) );
AND3_X1 _14897_ ( .A1(_06890_ ), .A2(_06705_ ), .A3(_06891_ ), .ZN(_06892_ ) );
MUX2_X1 _14898_ ( .A(_05668_ ), .B(_04296_ ), .S(_06731_ ), .Z(_06893_ ) );
AOI21_X1 _14899_ ( .A(_06892_ ), .B1(_06695_ ), .B2(_06893_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _14900_ ( .A1(_05278_ ), .A2(\mtvec [8] ), .A3(_04987_ ), .ZN(_06894_ ) );
NAND3_X1 _14901_ ( .A1(_05278_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_04843_ ), .ZN(_06895_ ) );
NAND3_X1 _14902_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_04895_ ), .ZN(_06896_ ) );
NAND4_X1 _14903_ ( .A1(_04934_ ), .A2(_05210_ ), .A3(\mepc [8] ), .A4(_05052_ ), .ZN(_06897_ ) );
NAND4_X1 _14904_ ( .A1(_06894_ ), .A2(_06895_ ), .A3(_06896_ ), .A4(_06897_ ), .ZN(_06898_ ) );
NOR4_X1 _14905_ ( .A1(_05103_ ), .A2(_06898_ ), .A3(_05013_ ), .A4(_04893_ ), .ZN(_06899_ ) );
AND3_X1 _14906_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_06606_ ), .ZN(_06900_ ) );
OAI21_X1 _14907_ ( .A(\ID_EX_typ [2] ), .B1(_06899_ ), .B2(_06900_ ), .ZN(_06901_ ) );
AOI21_X1 _14908_ ( .A(fanout_net_5 ), .B1(_02918_ ), .B2(_02937_ ), .ZN(_06902_ ) );
AND2_X1 _14909_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [8] ), .ZN(_06903_ ) );
OAI21_X1 _14910_ ( .A(_06901_ ), .B1(_06902_ ), .B2(_06903_ ), .ZN(_06904_ ) );
NOR3_X1 _14911_ ( .A1(_05583_ ), .A2(\EX_LS_result_csreg_mem [8] ), .A3(_04914_ ), .ZN(_06905_ ) );
INV_X1 _14912_ ( .A(_06905_ ), .ZN(_06906_ ) );
NAND2_X1 _14913_ ( .A1(_04904_ ), .A2(\mtvec [8] ), .ZN(_06907_ ) );
NAND4_X1 _14914_ ( .A1(_05014_ ), .A2(_06896_ ), .A3(_05255_ ), .A4(_06907_ ), .ZN(_06908_ ) );
NAND4_X1 _14915_ ( .A1(_04991_ ), .A2(_04992_ ), .A3(_04993_ ), .A4(\mycsreg.CSReg[0][8] ), .ZN(_06909_ ) );
OAI21_X1 _14916_ ( .A(_06909_ ), .B1(_05583_ ), .B2(_04914_ ), .ZN(_06910_ ) );
OAI211_X1 _14917_ ( .A(_06906_ ), .B(_06727_ ), .C1(_06908_ ), .C2(_06910_ ), .ZN(_06911_ ) );
AOI21_X1 _14918_ ( .A(_06694_ ), .B1(_06904_ ), .B2(_06911_ ), .ZN(_06912_ ) );
AND3_X1 _14919_ ( .A1(_03342_ ), .A2(_05263_ ), .A3(\ID_EX_typ [7] ), .ZN(_06913_ ) );
AOI211_X1 _14920_ ( .A(_06705_ ), .B(_06913_ ), .C1(_04319_ ), .C2(_06702_ ), .ZN(_06914_ ) );
OR2_X1 _14921_ ( .A1(_06912_ ), .A2(_06914_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
AOI21_X1 _14922_ ( .A(_06752_ ), .B1(_05286_ ), .B2(_05287_ ), .ZN(_06915_ ) );
NAND3_X1 _14923_ ( .A1(_02884_ ), .A2(_02419_ ), .A3(_02885_ ), .ZN(_06916_ ) );
NAND2_X1 _14924_ ( .A1(fanout_net_5 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_06917_ ) );
AOI21_X1 _14925_ ( .A(_06915_ ), .B1(_06916_ ), .B2(_06917_ ), .ZN(_06918_ ) );
AOI211_X1 _14926_ ( .A(_06694_ ), .B(_06918_ ), .C1(\ID_EX_typ [2] ), .C2(_05288_ ), .ZN(_06919_ ) );
AND4_X1 _14927_ ( .A1(_05294_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06920_ ) );
AOI211_X1 _14928_ ( .A(_06705_ ), .B(_06920_ ), .C1(_04342_ ), .C2(_06702_ ), .ZN(_06921_ ) );
OR2_X1 _14929_ ( .A1(_06919_ ), .A2(_06921_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
AND3_X1 _14930_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_06590_ ), .ZN(_06922_ ) );
NAND3_X1 _14931_ ( .A1(_06787_ ), .A2(\mtvec [6] ), .A3(_04987_ ), .ZN(_06923_ ) );
NAND3_X1 _14932_ ( .A1(_05278_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_05059_ ), .ZN(_06924_ ) );
NAND3_X1 _14933_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_04896_ ), .ZN(_06925_ ) );
NAND4_X1 _14934_ ( .A1(_05456_ ), .A2(_06717_ ), .A3(\mepc [6] ), .A4(_04899_ ), .ZN(_06926_ ) );
AND4_X1 _14935_ ( .A1(_06923_ ), .A2(_06924_ ), .A3(_06925_ ), .A4(_06926_ ), .ZN(_06927_ ) );
AOI21_X1 _14936_ ( .A(_06922_ ), .B1(_06821_ ), .B2(_06927_ ), .ZN(_06928_ ) );
NAND3_X1 _14937_ ( .A1(_06928_ ), .A2(_06802_ ), .A3(_06744_ ), .ZN(_06929_ ) );
MUX2_X1 _14938_ ( .A(_05317_ ), .B(_04364_ ), .S(_06701_ ), .Z(_06930_ ) );
OAI221_X1 _14939_ ( .A(_06697_ ), .B1(_05687_ ), .B2(\ID_EX_imm [6] ), .C1(_06928_ ), .C2(_05686_ ), .ZN(_06931_ ) );
AND3_X1 _14940_ ( .A1(_02888_ ), .A2(_04785_ ), .A3(_02907_ ), .ZN(_06932_ ) );
OAI221_X1 _14941_ ( .A(_06929_ ), .B1(_06706_ ), .B2(_06930_ ), .C1(_06931_ ), .C2(_06932_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14942_ ( .A(\ID_EX_pc [5] ), .B(_04411_ ), .S(_06701_ ), .Z(_06933_ ) );
NAND4_X1 _14943_ ( .A1(_05059_ ), .A2(_04845_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][5] ), .ZN(_06934_ ) );
OAI21_X1 _14944_ ( .A(_06934_ ), .B1(_04888_ ), .B2(_04890_ ), .ZN(_06935_ ) );
AOI22_X1 _14945_ ( .A1(_05391_ ), .A2(\mycsreg.CSReg[3][5] ), .B1(_04892_ ), .B2(_05456_ ), .ZN(_06936_ ) );
NAND2_X1 _14946_ ( .A1(_04904_ ), .A2(\mtvec [5] ), .ZN(_06937_ ) );
NAND3_X1 _14947_ ( .A1(_06936_ ), .A2(_05338_ ), .A3(_06937_ ), .ZN(_06938_ ) );
NOR2_X1 _14948_ ( .A1(_06935_ ), .A2(_06938_ ), .ZN(_06939_ ) );
NOR3_X1 _14949_ ( .A1(_04912_ ), .A2(\EX_LS_result_csreg_mem [5] ), .A3(_05216_ ), .ZN(_06940_ ) );
OAI21_X1 _14950_ ( .A(\ID_EX_typ [2] ), .B1(_06939_ ), .B2(_06940_ ), .ZN(_06941_ ) );
OR2_X1 _14951_ ( .A1(_02419_ ), .A2(\ID_EX_imm [5] ), .ZN(_06942_ ) );
NAND3_X1 _14952_ ( .A1(_02813_ ), .A2(_03516_ ), .A3(_02832_ ), .ZN(_06943_ ) );
NAND3_X1 _14953_ ( .A1(_06941_ ), .A2(_06942_ ), .A3(_06943_ ), .ZN(_06944_ ) );
INV_X1 _14954_ ( .A(_06940_ ), .ZN(_06945_ ) );
OAI211_X1 _14955_ ( .A(_06945_ ), .B(_06727_ ), .C1(_06938_ ), .C2(_06935_ ), .ZN(_06946_ ) );
NAND2_X1 _14956_ ( .A1(_06944_ ), .A2(_06946_ ), .ZN(_06947_ ) );
MUX2_X1 _14957_ ( .A(_06933_ ), .B(_06947_ ), .S(_06697_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
OAI21_X1 _14958_ ( .A(\ID_EX_typ [2] ), .B1(_05363_ ), .B2(_05367_ ), .ZN(_06948_ ) );
NAND3_X1 _14959_ ( .A1(_02853_ ), .A2(_05305_ ), .A3(_02854_ ), .ZN(_06949_ ) );
NAND2_X1 _14960_ ( .A1(_02856_ ), .A2(fanout_net_5 ), .ZN(_06950_ ) );
NAND3_X1 _14961_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_06950_ ), .ZN(_06951_ ) );
NAND3_X1 _14962_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_05366_ ), .ZN(_06952_ ) );
OAI211_X1 _14963_ ( .A(_06727_ ), .B(_06952_ ), .C1(_06822_ ), .C2(_05362_ ), .ZN(_06953_ ) );
AOI21_X1 _14964_ ( .A(_06694_ ), .B1(_06951_ ), .B2(_06953_ ), .ZN(_06954_ ) );
NOR2_X1 _14965_ ( .A1(_06754_ ), .A2(\ID_EX_pc [4] ), .ZN(_06955_ ) );
AOI211_X1 _14966_ ( .A(_06705_ ), .B(_06955_ ), .C1(_04389_ ), .C2(_06731_ ), .ZN(_06956_ ) );
OR2_X1 _14967_ ( .A1(_06954_ ), .A2(_06956_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14968_ ( .A(\ID_EX_pc [3] ), .B(_04106_ ), .S(_06701_ ), .Z(_06957_ ) );
NAND3_X1 _14969_ ( .A1(_02730_ ), .A2(_03516_ ), .A3(_02731_ ), .ZN(_06958_ ) );
OAI21_X1 _14970_ ( .A(\ID_EX_typ [2] ), .B1(_05398_ ), .B2(_05399_ ), .ZN(_06959_ ) );
NAND2_X1 _14971_ ( .A1(_02733_ ), .A2(fanout_net_5 ), .ZN(_06960_ ) );
NAND3_X1 _14972_ ( .A1(_06958_ ), .A2(_06959_ ), .A3(_06960_ ), .ZN(_06961_ ) );
OR3_X1 _14973_ ( .A1(_05583_ ), .A2(\EX_LS_result_csreg_mem [3] ), .A3(_05216_ ), .ZN(_06962_ ) );
NAND2_X1 _14974_ ( .A1(_04904_ ), .A2(\mtvec [3] ), .ZN(_06963_ ) );
OAI21_X1 _14975_ ( .A(_06963_ ), .B1(_05583_ ), .B2(_04914_ ), .ZN(_06964_ ) );
OAI211_X1 _14976_ ( .A(_06962_ ), .B(_06727_ ), .C1(_05396_ ), .C2(_06964_ ), .ZN(_06965_ ) );
NAND2_X1 _14977_ ( .A1(_06961_ ), .A2(_06965_ ), .ZN(_06966_ ) );
MUX2_X1 _14978_ ( .A(_06957_ ), .B(_06966_ ), .S(_06697_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
AND4_X1 _14979_ ( .A1(\mycsreg.CSReg[3][2] ), .A2(_04798_ ), .A3(_04799_ ), .A4(_04800_ ), .ZN(_06967_ ) );
AND4_X1 _14980_ ( .A1(\mepc [2] ), .A2(_04934_ ), .A3(_04798_ ), .A4(_04800_ ), .ZN(_06968_ ) );
NOR3_X1 _14981_ ( .A1(_04893_ ), .A2(_06967_ ), .A3(_06968_ ), .ZN(_06969_ ) );
NAND3_X1 _14982_ ( .A1(_04938_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_04842_ ), .ZN(_06970_ ) );
NAND3_X1 _14983_ ( .A1(_04938_ ), .A2(\mtvec [2] ), .A3(_03569_ ), .ZN(_06971_ ) );
AND2_X1 _14984_ ( .A1(_06970_ ), .A2(_06971_ ), .ZN(_06972_ ) );
AOI22_X1 _14985_ ( .A1(_06969_ ), .A2(_06972_ ), .B1(_04953_ ), .B2(_04959_ ), .ZN(_06973_ ) );
AND3_X1 _14986_ ( .A1(_04953_ ), .A2(_04959_ ), .A3(\EX_LS_result_csreg_mem [2] ), .ZN(_06974_ ) );
NOR2_X1 _14987_ ( .A1(_06973_ ), .A2(_06974_ ), .ZN(_06975_ ) );
AOI22_X1 _14988_ ( .A1(_06975_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02756_ ), .ZN(_06976_ ) );
OAI21_X1 _14989_ ( .A(_06976_ ), .B1(fanout_net_5 ), .B2(_02755_ ), .ZN(_06977_ ) );
OAI21_X1 _14990_ ( .A(_06727_ ), .B1(_06973_ ), .B2(_06974_ ), .ZN(_06978_ ) );
AND3_X1 _14991_ ( .A1(_06977_ ), .A2(_06705_ ), .A3(_06978_ ), .ZN(_06979_ ) );
MUX2_X1 _14992_ ( .A(_05669_ ), .B(_04128_ ), .S(_06731_ ), .Z(_06980_ ) );
AOI21_X1 _14993_ ( .A(_06979_ ), .B1(_06695_ ), .B2(_06980_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
NAND3_X1 _14994_ ( .A1(_05278_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_05059_ ), .ZN(_06981_ ) );
NAND3_X1 _14995_ ( .A1(_05278_ ), .A2(\mtvec [29] ), .A3(_04987_ ), .ZN(_06982_ ) );
NAND3_X1 _14996_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_06717_ ), .ZN(_06983_ ) );
NAND4_X1 _14997_ ( .A1(_05456_ ), .A2(_06717_ ), .A3(\mepc [29] ), .A4(_04845_ ), .ZN(_06984_ ) );
NAND4_X1 _14998_ ( .A1(_06981_ ), .A2(_06982_ ), .A3(_06983_ ), .A4(_06984_ ), .ZN(_06985_ ) );
NOR3_X1 _14999_ ( .A1(_05103_ ), .A2(_05013_ ), .A3(_06985_ ), .ZN(_06986_ ) );
NOR3_X1 _15000_ ( .A1(_05284_ ), .A2(_05285_ ), .A3(\EX_LS_result_csreg_mem [29] ), .ZN(_06987_ ) );
NOR2_X1 _15001_ ( .A1(_06986_ ), .A2(_06987_ ), .ZN(_06988_ ) );
OR3_X1 _15002_ ( .A1(_05284_ ), .A2(_05285_ ), .A3(\EX_LS_result_csreg_mem [29] ), .ZN(_06989_ ) );
OAI211_X1 _15003_ ( .A(_06726_ ), .B(_06989_ ), .C1(_06822_ ), .C2(_06985_ ), .ZN(_06990_ ) );
OAI21_X1 _15004_ ( .A(_06990_ ), .B1(_05687_ ), .B2(_03277_ ), .ZN(_06991_ ) );
AOI21_X1 _15005_ ( .A(fanout_net_5 ), .B1(_03256_ ), .B2(_03275_ ), .ZN(_06992_ ) );
OAI221_X1 _15006_ ( .A(_06711_ ), .B1(_05686_ ), .B2(_06988_ ), .C1(_06991_ ), .C2(_06992_ ), .ZN(_06993_ ) );
BUF_X4 _15007_ ( .A(_06694_ ), .Z(_06994_ ) );
NAND4_X1 _15008_ ( .A1(_03510_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06995_ ) );
OAI211_X1 _15009_ ( .A(_06994_ ), .B(_06995_ ), .C1(_03891_ ), .C2(_03343_ ), .ZN(_06996_ ) );
NAND2_X1 _15010_ ( .A1(_06993_ ), .A2(_06996_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR3_X1 _15011_ ( .A1(_04912_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_04890_ ), .ZN(_06997_ ) );
NAND3_X1 _15012_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_04984_ ), .ZN(_06998_ ) );
NAND2_X1 _15013_ ( .A1(_04904_ ), .A2(\mtvec [1] ), .ZN(_06999_ ) );
NAND4_X1 _15014_ ( .A1(_05190_ ), .A2(_04985_ ), .A3(_05127_ ), .A4(\mycsreg.CSReg[0][1] ), .ZN(_07000_ ) );
AND4_X1 _15015_ ( .A1(_06998_ ), .A2(_06999_ ), .A3(_05437_ ), .A4(_07000_ ), .ZN(_07001_ ) );
OAI21_X1 _15016_ ( .A(_07001_ ), .B1(_05583_ ), .B2(_04914_ ), .ZN(_07002_ ) );
NAND2_X1 _15017_ ( .A1(_06997_ ), .A2(_07002_ ), .ZN(_07003_ ) );
AOI22_X1 _15018_ ( .A1(_07003_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_07004_ ) );
OAI211_X1 _15019_ ( .A(_07004_ ), .B(_06750_ ), .C1(_02779_ ), .C2(fanout_net_5 ), .ZN(_07005_ ) );
NAND4_X1 _15020_ ( .A1(_06997_ ), .A2(_06802_ ), .A3(_06744_ ), .A4(_07002_ ), .ZN(_07006_ ) );
MUX2_X1 _15021_ ( .A(_05670_ ), .B(_04056_ ), .S(_06754_ ), .Z(_07007_ ) );
OAI211_X1 _15022_ ( .A(_07005_ ), .B(_07006_ ), .C1(_06730_ ), .C2(_07007_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
OR3_X1 _15023_ ( .A1(_04888_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_04890_ ), .ZN(_07008_ ) );
NAND4_X1 _15024_ ( .A1(_04843_ ), .A2(_04845_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][0] ), .ZN(_07009_ ) );
AND2_X1 _15025_ ( .A1(_05480_ ), .A2(_07009_ ), .ZN(_07010_ ) );
OAI21_X1 _15026_ ( .A(_07010_ ), .B1(_05583_ ), .B2(_04914_ ), .ZN(_07011_ ) );
NAND4_X1 _15027_ ( .A1(_04896_ ), .A2(_04897_ ), .A3(\mycsreg.CSReg[3][0] ), .A4(_04899_ ), .ZN(_07012_ ) );
INV_X1 _15028_ ( .A(\mtvec [0] ), .ZN(_07013_ ) );
OR3_X1 _15029_ ( .A1(_04901_ ), .A2(_07013_ ), .A3(_04902_ ), .ZN(_07014_ ) );
NAND3_X1 _15030_ ( .A1(_04894_ ), .A2(_07012_ ), .A3(_07014_ ), .ZN(_07015_ ) );
OAI21_X1 _15031_ ( .A(_07008_ ), .B1(_07011_ ), .B2(_07015_ ), .ZN(_07016_ ) );
AOI22_X1 _15032_ ( .A1(_07016_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02782_ ), .ZN(_07017_ ) );
OAI211_X1 _15033_ ( .A(_07017_ ), .B(_06750_ ), .C1(\ID_EX_typ [0] ), .C2(_04058_ ), .ZN(_07018_ ) );
OR3_X1 _15034_ ( .A1(_07016_ ), .A2(_06693_ ), .A3(_06752_ ), .ZN(_07019_ ) );
AOI21_X1 _15035_ ( .A(_03343_ ), .B1(_04078_ ), .B2(_04080_ ), .ZN(_07020_ ) );
AOI21_X1 _15036_ ( .A(_07020_ ), .B1(\ID_EX_pc [0] ), .B2(_03343_ ), .ZN(_07021_ ) );
OAI211_X1 _15037_ ( .A(_07018_ ), .B(_07019_ ), .C1(_06698_ ), .C2(_07021_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
OR3_X1 _15038_ ( .A1(_05022_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_04913_ ), .ZN(_07022_ ) );
AOI22_X1 _15039_ ( .A1(_05391_ ), .A2(\mycsreg.CSReg[3][28] ), .B1(_04892_ ), .B2(_05456_ ), .ZN(_07023_ ) );
NAND4_X1 _15040_ ( .A1(_05059_ ), .A2(_04899_ ), .A3(_04847_ ), .A4(\mycsreg.CSReg[0][28] ), .ZN(_07024_ ) );
NAND3_X1 _15041_ ( .A1(_07023_ ), .A2(_05186_ ), .A3(_07024_ ), .ZN(_07025_ ) );
OR3_X1 _15042_ ( .A1(_04901_ ), .A2(_06356_ ), .A3(_04902_ ), .ZN(_07026_ ) );
OAI21_X1 _15043_ ( .A(_07026_ ), .B1(_04912_ ), .B2(_05216_ ), .ZN(_07027_ ) );
OAI21_X1 _15044_ ( .A(_07022_ ), .B1(_07025_ ), .B2(_07027_ ), .ZN(_07028_ ) );
AOI22_X1 _15045_ ( .A1(_04750_ ), .A2(_04785_ ), .B1(\ID_EX_typ [2] ), .B2(_07028_ ), .ZN(_07029_ ) );
OAI211_X1 _15046_ ( .A(_07029_ ), .B(_06750_ ), .C1(_05687_ ), .C2(\ID_EX_imm [28] ), .ZN(_07030_ ) );
OR3_X1 _15047_ ( .A1(_07028_ ), .A2(_06693_ ), .A3(_06752_ ), .ZN(_07031_ ) );
AND3_X1 _15048_ ( .A1(_03342_ ), .A2(\ID_EX_pc [28] ), .A3(\ID_EX_typ [7] ), .ZN(_07032_ ) );
AOI21_X1 _15049_ ( .A(_07032_ ), .B1(_03869_ ), .B2(_06702_ ), .ZN(_07033_ ) );
OAI211_X1 _15050_ ( .A(_07030_ ), .B(_07031_ ), .C1(_06698_ ), .C2(_07033_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
OR3_X1 _15051_ ( .A1(_05284_ ), .A2(_05285_ ), .A3(\EX_LS_result_csreg_mem [27] ), .ZN(_07034_ ) );
NAND3_X1 _15052_ ( .A1(_06787_ ), .A2(\mtvec [27] ), .A3(_04987_ ), .ZN(_07035_ ) );
NAND3_X1 _15053_ ( .A1(_06787_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_04991_ ), .ZN(_07036_ ) );
NAND3_X1 _15054_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_04896_ ), .ZN(_07037_ ) );
NAND4_X1 _15055_ ( .A1(_05456_ ), .A2(_04896_ ), .A3(\mepc [27] ), .A4(_04992_ ), .ZN(_07038_ ) );
NAND4_X1 _15056_ ( .A1(_07035_ ), .A2(_07036_ ), .A3(_07037_ ), .A4(_07038_ ), .ZN(_07039_ ) );
OAI211_X1 _15057_ ( .A(_07034_ ), .B(_06727_ ), .C1(_06822_ ), .C2(_07039_ ), .ZN(_07040_ ) );
NAND2_X1 _15058_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [27] ), .ZN(_07041_ ) );
NAND2_X1 _15059_ ( .A1(_07040_ ), .A2(_07041_ ), .ZN(_07042_ ) );
AOI21_X1 _15060_ ( .A(\ID_EX_typ [0] ), .B1(_02483_ ), .B2(_02493_ ), .ZN(_07043_ ) );
OAI221_X1 _15061_ ( .A(_06711_ ), .B1(_05686_ ), .B2(_05463_ ), .C1(_07042_ ), .C2(_07043_ ), .ZN(_07044_ ) );
NAND4_X1 _15062_ ( .A1(_04817_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_07045_ ) );
OAI211_X1 _15063_ ( .A(_06994_ ), .B(_07045_ ), .C1(_04009_ ), .C2(_03343_ ), .ZN(_07046_ ) );
NAND2_X1 _15064_ ( .A1(_07044_ ), .A2(_07046_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
OR3_X1 _15065_ ( .A1(_04888_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_04890_ ), .ZN(_07047_ ) );
NAND3_X1 _15066_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_04984_ ), .ZN(_07048_ ) );
NAND2_X1 _15067_ ( .A1(_04904_ ), .A2(\mtvec [26] ), .ZN(_07049_ ) );
NAND4_X1 _15068_ ( .A1(_05190_ ), .A2(_04985_ ), .A3(_05127_ ), .A4(\mycsreg.CSReg[0][26] ), .ZN(_07050_ ) );
AND4_X1 _15069_ ( .A1(_07048_ ), .A2(_07049_ ), .A3(_05505_ ), .A4(_07050_ ), .ZN(_07051_ ) );
OAI21_X1 _15070_ ( .A(_07051_ ), .B1(_05583_ ), .B2(_04914_ ), .ZN(_07052_ ) );
NAND2_X1 _15071_ ( .A1(_07047_ ), .A2(_07052_ ), .ZN(_07053_ ) );
AOI22_X1 _15072_ ( .A1(_07053_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_07054_ ) );
OAI211_X1 _15073_ ( .A(_07054_ ), .B(_06750_ ), .C1(\ID_EX_typ [0] ), .C2(_03221_ ), .ZN(_07055_ ) );
NAND4_X1 _15074_ ( .A1(_07047_ ), .A2(_06802_ ), .A3(_06744_ ), .A4(_07052_ ), .ZN(_07056_ ) );
AND3_X1 _15075_ ( .A1(_03342_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_07057_ ) );
AOI21_X1 _15076_ ( .A(_07057_ ), .B1(_04031_ ), .B2(_06702_ ), .ZN(_07058_ ) );
OAI211_X1 _15077_ ( .A(_07055_ ), .B(_07056_ ), .C1(_06698_ ), .C2(_07058_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
AOI22_X1 _15078_ ( .A1(_05539_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_03224_ ), .ZN(_07059_ ) );
OAI211_X1 _15079_ ( .A(_07059_ ), .B(_06750_ ), .C1(_03198_ ), .C2(\ID_EX_typ [0] ), .ZN(_07060_ ) );
NAND4_X1 _15080_ ( .A1(_05532_ ), .A2(_06750_ ), .A3(_06744_ ), .A4(_05538_ ), .ZN(_07061_ ) );
AND3_X1 _15081_ ( .A1(_03342_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_07062_ ) );
AOI21_X1 _15082_ ( .A(_07062_ ), .B1(_03984_ ), .B2(_06702_ ), .ZN(_07063_ ) );
OAI211_X1 _15083_ ( .A(_07060_ ), .B(_07061_ ), .C1(_06698_ ), .C2(_07063_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
OR3_X1 _15084_ ( .A1(_04888_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_04890_ ), .ZN(_07064_ ) );
NAND3_X1 _15085_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_06717_ ), .ZN(_07065_ ) );
OR3_X1 _15086_ ( .A1(_04901_ ), .A2(_06383_ ), .A3(_04902_ ), .ZN(_07066_ ) );
NAND4_X1 _15087_ ( .A1(_06715_ ), .A2(_04894_ ), .A3(_07065_ ), .A4(_07066_ ), .ZN(_07067_ ) );
NAND4_X1 _15088_ ( .A1(_05190_ ), .A2(_04898_ ), .A3(_04988_ ), .A4(\mycsreg.CSReg[0][24] ), .ZN(_07068_ ) );
AND2_X1 _15089_ ( .A1(_05548_ ), .A2(_07068_ ), .ZN(_07069_ ) );
OAI21_X1 _15090_ ( .A(_07069_ ), .B1(_04912_ ), .B2(_05216_ ), .ZN(_07070_ ) );
OAI21_X1 _15091_ ( .A(_07064_ ), .B1(_07067_ ), .B2(_07070_ ), .ZN(_07071_ ) );
AOI22_X1 _15092_ ( .A1(_04785_ ), .A2(_04483_ ), .B1(_07071_ ), .B2(\ID_EX_typ [2] ), .ZN(_07072_ ) );
OAI211_X1 _15093_ ( .A(_07072_ ), .B(_06750_ ), .C1(_05687_ ), .C2(\ID_EX_imm [24] ), .ZN(_07073_ ) );
OR3_X1 _15094_ ( .A1(_07071_ ), .A2(_06693_ ), .A3(_06752_ ), .ZN(_07074_ ) );
AND3_X1 _15095_ ( .A1(_03342_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_typ [7] ), .ZN(_07075_ ) );
AOI21_X1 _15096_ ( .A(_07075_ ), .B1(_03961_ ), .B2(_06702_ ), .ZN(_07076_ ) );
OAI211_X1 _15097_ ( .A(_07073_ ), .B(_07074_ ), .C1(_06698_ ), .C2(_07076_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
AOI22_X1 _15098_ ( .A1(_05585_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02544_ ), .ZN(_07077_ ) );
OAI211_X1 _15099_ ( .A(_07077_ ), .B(_06697_ ), .C1(_02548_ ), .C2(\ID_EX_typ [0] ), .ZN(_07078_ ) );
NAND4_X1 _15100_ ( .A1(_05577_ ), .A2(_06750_ ), .A3(_06744_ ), .A4(_05584_ ), .ZN(_07079_ ) );
MUX2_X1 _15101_ ( .A(_05671_ ), .B(_03816_ ), .S(_06754_ ), .Z(_07080_ ) );
OAI211_X1 _15102_ ( .A(_07078_ ), .B(_07079_ ), .C1(_06698_ ), .C2(_07080_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
INV_X1 _15103_ ( .A(_05602_ ), .ZN(_07081_ ) );
OR3_X1 _15104_ ( .A1(_05284_ ), .A2(_05285_ ), .A3(\EX_LS_result_csreg_mem [22] ), .ZN(_07082_ ) );
NAND2_X1 _15105_ ( .A1(_06821_ ), .A2(_04894_ ), .ZN(_07083_ ) );
NAND3_X1 _15106_ ( .A1(_04939_ ), .A2(\mtvec [22] ), .A3(_04940_ ), .ZN(_07084_ ) );
NAND3_X1 _15107_ ( .A1(_04939_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_04942_ ), .ZN(_07085_ ) );
NAND4_X1 _15108_ ( .A1(_04934_ ), .A2(_04838_ ), .A3(\mepc [22] ), .A4(_04833_ ), .ZN(_07086_ ) );
NAND4_X1 _15109_ ( .A1(_07084_ ), .A2(_07085_ ), .A3(_05594_ ), .A4(_07086_ ), .ZN(_07087_ ) );
OAI211_X1 _15110_ ( .A(_06726_ ), .B(_07082_ ), .C1(_07083_ ), .C2(_07087_ ), .ZN(_07088_ ) );
NAND2_X1 _15111_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [22] ), .ZN(_07089_ ) );
AND2_X1 _15112_ ( .A1(_07088_ ), .A2(_07089_ ), .ZN(_07090_ ) );
NAND2_X1 _15113_ ( .A1(_02522_ ), .A2(_02419_ ), .ZN(_07091_ ) );
AOI221_X4 _15114_ ( .A(_06693_ ), .B1(\ID_EX_typ [2] ), .B2(_07081_ ), .C1(_07090_ ), .C2(_07091_ ), .ZN(_07092_ ) );
NOR4_X1 _15115_ ( .A1(_02406_ ), .A2(_02409_ ), .A3(_02412_ ), .A4(\ID_EX_pc [22] ), .ZN(_07093_ ) );
AOI211_X1 _15116_ ( .A(_06705_ ), .B(_07093_ ), .C1(_03838_ ), .C2(_06731_ ), .ZN(_07094_ ) );
OR2_X1 _15117_ ( .A1(_07092_ ), .A2(_07094_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
OR3_X1 _15118_ ( .A1(_04888_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_04890_ ), .ZN(_07095_ ) );
NAND3_X1 _15119_ ( .A1(_05016_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_04984_ ), .ZN(_07096_ ) );
OR3_X1 _15120_ ( .A1(_04901_ ), .A2(_06402_ ), .A3(_04902_ ), .ZN(_07097_ ) );
NAND4_X1 _15121_ ( .A1(_05190_ ), .A2(_05126_ ), .A3(_05127_ ), .A4(\mycsreg.CSReg[0][31] ), .ZN(_07098_ ) );
AND4_X1 _15122_ ( .A1(_07096_ ), .A2(_07097_ ), .A3(_05650_ ), .A4(_07098_ ), .ZN(_07099_ ) );
OAI21_X1 _15123_ ( .A(_07099_ ), .B1(_05583_ ), .B2(_04914_ ), .ZN(_07100_ ) );
NAND2_X1 _15124_ ( .A1(_07095_ ), .A2(_07100_ ), .ZN(_07101_ ) );
AOI22_X1 _15125_ ( .A1(_07101_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_07102_ ) );
OAI211_X1 _15126_ ( .A(_07102_ ), .B(_06697_ ), .C1(_03337_ ), .C2(\ID_EX_typ [0] ), .ZN(_07103_ ) );
NAND4_X1 _15127_ ( .A1(_07095_ ), .A2(_06750_ ), .A3(_06744_ ), .A4(_07100_ ), .ZN(_07104_ ) );
AND3_X1 _15128_ ( .A1(_03342_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_07105_ ) );
AOI21_X1 _15129_ ( .A(_07105_ ), .B1(_03916_ ), .B2(_06702_ ), .ZN(_07106_ ) );
OAI211_X1 _15130_ ( .A(_07103_ ), .B(_07104_ ), .C1(_07106_ ), .C2(_06698_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
OAI21_X1 _15131_ ( .A(_06711_ ), .B1(_05626_ ), .B2(_05632_ ), .ZN(_07107_ ) );
NOR3_X1 _15132_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_07108_ ) );
AND2_X2 _15133_ ( .A1(fanout_net_6 ), .A2(\ID_EX_typ [2] ), .ZN(_07109_ ) );
AND2_X2 _15134_ ( .A1(_07108_ ), .A2(_07109_ ), .ZN(_07110_ ) );
INV_X1 _15135_ ( .A(_07110_ ), .ZN(_07111_ ) );
NOR3_X1 _15136_ ( .A1(_04417_ ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_07112_ ) );
AND2_X1 _15137_ ( .A1(_07112_ ), .A2(_07109_ ), .ZN(_07113_ ) );
BUF_X4 _15138_ ( .A(_07113_ ), .Z(_07114_ ) );
INV_X2 _15139_ ( .A(_07114_ ), .ZN(_07115_ ) );
OAI22_X1 _15140_ ( .A1(_05619_ ), .A2(_07111_ ), .B1(_02576_ ), .B2(_07115_ ), .ZN(_07116_ ) );
NAND2_X1 _15141_ ( .A1(_04457_ ), .A2(_03748_ ), .ZN(_07117_ ) );
AND2_X1 _15142_ ( .A1(_07117_ ), .A2(_04467_ ), .ZN(_07118_ ) );
INV_X1 _15143_ ( .A(_03770_ ), .ZN(_07119_ ) );
NOR2_X1 _15144_ ( .A1(_07118_ ), .A2(_07119_ ), .ZN(_07120_ ) );
NOR2_X1 _15145_ ( .A1(_07120_ ), .A2(_04473_ ), .ZN(_07121_ ) );
XNOR2_X1 _15146_ ( .A(_07121_ ), .B(_03794_ ), .ZN(_07122_ ) );
AND3_X1 _15147_ ( .A1(_03602_ ), .A2(\ID_EX_typ [3] ), .A3(_04771_ ), .ZN(_07123_ ) );
AND2_X1 _15148_ ( .A1(_07123_ ), .A2(_04511_ ), .ZN(_07124_ ) );
BUF_X2 _15149_ ( .A(_07124_ ), .Z(_07125_ ) );
BUF_X2 _15150_ ( .A(_07125_ ), .Z(_07126_ ) );
AOI21_X1 _15151_ ( .A(_07116_ ), .B1(_07122_ ), .B2(_07126_ ), .ZN(_07127_ ) );
AOI21_X1 _15152_ ( .A(_05495_ ), .B1(_07127_ ), .B2(_05672_ ), .ZN(_07128_ ) );
AND2_X1 _15153_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .ZN(_07129_ ) );
AND2_X2 _15154_ ( .A1(_07129_ ), .A2(\ID_EX_typ [2] ), .ZN(_07130_ ) );
BUF_X4 _15155_ ( .A(_07130_ ), .Z(_07131_ ) );
NAND2_X1 _15156_ ( .A1(_04651_ ), .A2(_04652_ ), .ZN(_07132_ ) );
AND2_X1 _15157_ ( .A1(_04647_ ), .A2(_07132_ ), .ZN(_07133_ ) );
AND2_X1 _15158_ ( .A1(_07133_ ), .A2(_04640_ ), .ZN(_07134_ ) );
AND2_X1 _15159_ ( .A1(_07134_ ), .A2(_04643_ ), .ZN(_07135_ ) );
AND2_X1 _15160_ ( .A1(_07135_ ), .A2(_04629_ ), .ZN(_07136_ ) );
XNOR2_X1 _15161_ ( .A(_07136_ ), .B(_04625_ ), .ZN(_07137_ ) );
INV_X2 _15162_ ( .A(_07137_ ), .ZN(_07138_ ) );
AND3_X1 _15163_ ( .A1(_04610_ ), .A2(_04611_ ), .A3(_04619_ ), .ZN(_07139_ ) );
AND3_X1 _15164_ ( .A1(_04556_ ), .A2(_04557_ ), .A3(_04554_ ), .ZN(_07140_ ) );
AND3_X1 _15165_ ( .A1(_04571_ ), .A2(_04566_ ), .A3(_04565_ ), .ZN(_07141_ ) );
AND2_X1 _15166_ ( .A1(_04549_ ), .A2(_04545_ ), .ZN(_07142_ ) );
AND4_X1 _15167_ ( .A1(_07139_ ), .A2(_07140_ ), .A3(_07141_ ), .A4(_07142_ ), .ZN(_07143_ ) );
AND4_X1 _15168_ ( .A1(_04590_ ), .A2(_04596_ ), .A3(_04665_ ), .A4(_04669_ ), .ZN(_07144_ ) );
AND2_X1 _15169_ ( .A1(_04601_ ), .A2(_04606_ ), .ZN(_07145_ ) );
AND2_X1 _15170_ ( .A1(_04579_ ), .A2(_04584_ ), .ZN(_07146_ ) );
AND4_X1 _15171_ ( .A1(_07143_ ), .A2(_07144_ ), .A3(_07145_ ), .A4(_07146_ ), .ZN(_07147_ ) );
OAI21_X1 _15172_ ( .A(_07147_ ), .B1(_07136_ ), .B2(_04661_ ), .ZN(_07148_ ) );
INV_X1 _15173_ ( .A(_04539_ ), .ZN(_07149_ ) );
INV_X1 _15174_ ( .A(_04535_ ), .ZN(_07150_ ) );
NOR3_X1 _15175_ ( .A1(_07148_ ), .A2(_07149_ ), .A3(_07150_ ), .ZN(_07151_ ) );
INV_X1 _15176_ ( .A(_04735_ ), .ZN(_07152_ ) );
NOR4_X1 _15177_ ( .A1(_04741_ ), .A2(_07152_ ), .A3(_04524_ ), .A4(_04529_ ), .ZN(_07153_ ) );
INV_X1 _15178_ ( .A(_04514_ ), .ZN(_07154_ ) );
AND4_X1 _15179_ ( .A1(_04716_ ), .A2(_04759_ ), .A3(_04721_ ), .A4(_07154_ ), .ZN(_07155_ ) );
AND3_X1 _15180_ ( .A1(_07151_ ), .A2(_07153_ ), .A3(_07155_ ), .ZN(_07156_ ) );
AND4_X1 _15181_ ( .A1(_04741_ ), .A2(_07152_ ), .A3(_04524_ ), .A4(_04529_ ), .ZN(_07157_ ) );
NAND4_X1 _15182_ ( .A1(_07157_ ), .A2(_04718_ ), .A3(_04720_ ), .A4(_04758_ ), .ZN(_07158_ ) );
NOR3_X1 _15183_ ( .A1(_07158_ ), .A2(_04716_ ), .A3(_07154_ ), .ZN(_07159_ ) );
AND2_X1 _15184_ ( .A1(_07139_ ), .A2(_07146_ ), .ZN(_07160_ ) );
AND4_X1 _15185_ ( .A1(_04590_ ), .A2(_07160_ ), .A3(_04596_ ), .A4(_07145_ ), .ZN(_07161_ ) );
AND4_X1 _15186_ ( .A1(_04665_ ), .A2(_04625_ ), .A3(_04669_ ), .A4(_04629_ ), .ZN(_07162_ ) );
NAND3_X1 _15187_ ( .A1(_07162_ ), .A2(_07134_ ), .A3(_04643_ ), .ZN(_07163_ ) );
NAND4_X1 _15188_ ( .A1(_04665_ ), .A2(_04623_ ), .A3(_04669_ ), .A4(_04624_ ), .ZN(_07164_ ) );
NAND2_X1 _15189_ ( .A1(_07163_ ), .A2(_07164_ ), .ZN(_07165_ ) );
AND2_X1 _15190_ ( .A1(_07161_ ), .A2(_07165_ ), .ZN(_07166_ ) );
AND2_X1 _15191_ ( .A1(_07140_ ), .A2(_07141_ ), .ZN(_07167_ ) );
AND3_X1 _15192_ ( .A1(_07166_ ), .A2(_07142_ ), .A3(_07167_ ), .ZN(_07168_ ) );
NAND3_X1 _15193_ ( .A1(_07168_ ), .A2(_04539_ ), .A3(_04535_ ), .ZN(_07169_ ) );
AOI21_X1 _15194_ ( .A(_07156_ ), .B1(_07159_ ), .B2(_07169_ ), .ZN(_07170_ ) );
OR3_X1 _15195_ ( .A1(_07148_ ), .A2(_07149_ ), .A3(_07150_ ), .ZN(_07171_ ) );
NAND3_X1 _15196_ ( .A1(_07148_ ), .A2(_07149_ ), .A3(_07150_ ), .ZN(_07172_ ) );
NAND2_X1 _15197_ ( .A1(_07171_ ), .A2(_07172_ ), .ZN(_07173_ ) );
INV_X1 _15198_ ( .A(_03337_ ), .ZN(_07174_ ) );
INV_X1 _15199_ ( .A(_04584_ ), .ZN(_07175_ ) );
NOR4_X1 _15200_ ( .A1(_04590_ ), .A2(_04596_ ), .A3(_04665_ ), .A4(_04669_ ), .ZN(_07176_ ) );
AOI22_X1 _15201_ ( .A1(_04600_ ), .A2(_04599_ ), .B1(_04604_ ), .B2(_04605_ ), .ZN(_07177_ ) );
AND4_X1 _15202_ ( .A1(_07175_ ), .A2(_07176_ ), .A3(_04680_ ), .A4(_07177_ ), .ZN(_07178_ ) );
NOR4_X1 _15203_ ( .A1(_04612_ ), .A2(_04567_ ), .A3(_04571_ ), .A4(_04619_ ), .ZN(_07179_ ) );
NOR4_X1 _15204_ ( .A1(_04558_ ), .A2(_04545_ ), .A3(_04549_ ), .A4(_04554_ ), .ZN(_07180_ ) );
AND3_X1 _15205_ ( .A1(_07178_ ), .A2(_07179_ ), .A3(_07180_ ), .ZN(_07181_ ) );
INV_X1 _15206_ ( .A(_07136_ ), .ZN(_07182_ ) );
NAND3_X1 _15207_ ( .A1(_07181_ ), .A2(_04625_ ), .A3(_07182_ ), .ZN(_07183_ ) );
AOI21_X1 _15208_ ( .A(_07174_ ), .B1(_07183_ ), .B2(_07148_ ), .ZN(_07184_ ) );
NAND2_X1 _15209_ ( .A1(_07173_ ), .A2(_07184_ ), .ZN(_07185_ ) );
NOR2_X1 _15210_ ( .A1(_07170_ ), .A2(_07185_ ), .ZN(_07186_ ) );
XNOR2_X1 _15211_ ( .A(_07135_ ), .B(_04630_ ), .ZN(_07187_ ) );
NOR2_X1 _15212_ ( .A1(_07186_ ), .A2(_07187_ ), .ZN(_07188_ ) );
OR4_X1 _15213_ ( .A1(_04567_ ), .A2(_04590_ ), .A3(_04571_ ), .A4(_04596_ ), .ZN(_07189_ ) );
OR3_X1 _15214_ ( .A1(_07189_ ), .A2(_04545_ ), .A3(_04554_ ), .ZN(_07190_ ) );
NOR3_X1 _15215_ ( .A1(_07190_ ), .A2(_04549_ ), .A3(_04558_ ), .ZN(_07191_ ) );
OR3_X1 _15216_ ( .A1(_04612_ ), .A2(_04601_ ), .A3(_04619_ ), .ZN(_07192_ ) );
OR4_X1 _15217_ ( .A1(_04584_ ), .A2(_04665_ ), .A3(_04669_ ), .A4(_04579_ ), .ZN(_07193_ ) );
NOR3_X1 _15218_ ( .A1(_07192_ ), .A2(_04606_ ), .A3(_07193_ ), .ZN(_07194_ ) );
NAND4_X1 _15219_ ( .A1(_07191_ ), .A2(_07182_ ), .A3(_04625_ ), .A4(_07194_ ), .ZN(_07195_ ) );
INV_X1 _15220_ ( .A(_07168_ ), .ZN(_07196_ ) );
NAND2_X1 _15221_ ( .A1(_07195_ ), .A2(_07196_ ), .ZN(_07197_ ) );
NAND3_X1 _15222_ ( .A1(_07197_ ), .A2(_03337_ ), .A3(_07173_ ), .ZN(_07198_ ) );
NOR2_X1 _15223_ ( .A1(_07170_ ), .A2(_07198_ ), .ZN(_07199_ ) );
BUF_X2 _15224_ ( .A(_07199_ ), .Z(_07200_ ) );
BUF_X4 _15225_ ( .A(_04647_ ), .Z(_07201_ ) );
BUF_X2 _15226_ ( .A(_07201_ ), .Z(_07202_ ) );
BUF_X4 _15227_ ( .A(_07132_ ), .Z(_07203_ ) );
BUF_X4 _15228_ ( .A(_07203_ ), .Z(_07204_ ) );
XNOR2_X1 _15229_ ( .A(_07202_ ), .B(_07204_ ), .ZN(_07205_ ) );
BUF_X4 _15230_ ( .A(_04641_ ), .Z(_07206_ ) );
NOR2_X1 _15231_ ( .A1(_07205_ ), .A2(_07206_ ), .ZN(_07207_ ) );
INV_X1 _15232_ ( .A(_07207_ ), .ZN(_07208_ ) );
BUF_X4 _15233_ ( .A(_04635_ ), .Z(_07209_ ) );
XNOR2_X1 _15234_ ( .A(_07134_ ), .B(_07209_ ), .ZN(_07210_ ) );
INV_X1 _15235_ ( .A(_07210_ ), .ZN(_07211_ ) );
BUF_X2 _15236_ ( .A(_07211_ ), .Z(_07212_ ) );
NAND3_X1 _15237_ ( .A1(_07200_ ), .A2(_07208_ ), .A3(_07212_ ), .ZN(_07213_ ) );
AOI211_X1 _15238_ ( .A(_07138_ ), .B(_07188_ ), .C1(_07187_ ), .C2(_07213_ ), .ZN(_07214_ ) );
BUF_X2 _15239_ ( .A(_04651_ ), .Z(_07215_ ) );
BUF_X2 _15240_ ( .A(_04652_ ), .Z(_07216_ ) );
AOI21_X1 _15241_ ( .A(_03987_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07217_ ) );
NOR2_X1 _15242_ ( .A1(_03253_ ), .A2(_07203_ ), .ZN(_07218_ ) );
NOR3_X1 _15243_ ( .A1(_07217_ ), .A2(_07218_ ), .A3(_07201_ ), .ZN(_07219_ ) );
INV_X2 _15244_ ( .A(_07201_ ), .ZN(_07220_ ) );
CLKBUF_X2 _15245_ ( .A(_04651_ ), .Z(_07221_ ) );
CLKBUF_X3 _15246_ ( .A(_04652_ ), .Z(_07222_ ) );
AND3_X1 _15247_ ( .A1(_03227_ ), .A2(_07221_ ), .A3(_07222_ ), .ZN(_07223_ ) );
BUF_X2 _15248_ ( .A(_04651_ ), .Z(_07224_ ) );
BUF_X2 _15249_ ( .A(_04652_ ), .Z(_07225_ ) );
AOI21_X1 _15250_ ( .A(_03198_ ), .B1(_07224_ ), .B2(_07225_ ), .ZN(_07226_ ) );
NOR3_X1 _15251_ ( .A1(_07220_ ), .A2(_07223_ ), .A3(_07226_ ), .ZN(_07227_ ) );
OAI21_X1 _15252_ ( .A(_04641_ ), .B1(_07219_ ), .B2(_07227_ ), .ZN(_07228_ ) );
BUF_X4 _15253_ ( .A(_07201_ ), .Z(_07229_ ) );
NOR2_X1 _15254_ ( .A1(_07203_ ), .A2(_02522_ ), .ZN(_07230_ ) );
AOI21_X1 _15255_ ( .A(_02575_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07231_ ) );
OAI21_X1 _15256_ ( .A(_07229_ ), .B1(_07230_ ), .B2(_07231_ ), .ZN(_07232_ ) );
BUF_X2 _15257_ ( .A(_07221_ ), .Z(_07233_ ) );
BUF_X2 _15258_ ( .A(_07222_ ), .Z(_07234_ ) );
AOI21_X1 _15259_ ( .A(_02548_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07235_ ) );
AND3_X1 _15260_ ( .A1(_04483_ ), .A2(_07221_ ), .A3(_07222_ ), .ZN(_07236_ ) );
OAI21_X1 _15261_ ( .A(_07220_ ), .B1(_07235_ ), .B2(_07236_ ), .ZN(_07237_ ) );
NAND3_X1 _15262_ ( .A1(_07232_ ), .A2(_07237_ ), .A3(_04640_ ), .ZN(_07238_ ) );
NAND2_X1 _15263_ ( .A1(_07228_ ), .A2(_07238_ ), .ZN(_07239_ ) );
AND2_X1 _15264_ ( .A1(_07132_ ), .A2(_03337_ ), .ZN(_07240_ ) );
INV_X1 _15265_ ( .A(_07240_ ), .ZN(_07241_ ) );
INV_X1 _15266_ ( .A(_07132_ ), .ZN(_07242_ ) );
AND2_X1 _15267_ ( .A1(_03310_ ), .A2(_07242_ ), .ZN(_07243_ ) );
AOI21_X1 _15268_ ( .A(_03276_ ), .B1(_07221_ ), .B2(_07222_ ), .ZN(_07244_ ) );
OR2_X1 _15269_ ( .A1(_07243_ ), .A2(_07244_ ), .ZN(_07245_ ) );
MUX2_X1 _15270_ ( .A(_07241_ ), .B(_07245_ ), .S(_07201_ ), .Z(_07246_ ) );
NOR2_X1 _15271_ ( .A1(_07246_ ), .A2(_04641_ ), .ZN(_07247_ ) );
MUX2_X1 _15272_ ( .A(_07239_ ), .B(_07247_ ), .S(_07209_ ), .Z(_07248_ ) );
BUF_X2 _15273_ ( .A(_04629_ ), .Z(_07249_ ) );
BUF_X2 _15274_ ( .A(_07249_ ), .Z(_07250_ ) );
BUF_X2 _15275_ ( .A(_07250_ ), .Z(_07251_ ) );
AND2_X1 _15276_ ( .A1(_07248_ ), .A2(_07251_ ), .ZN(_07252_ ) );
OAI21_X1 _15277_ ( .A(_07131_ ), .B1(_07214_ ), .B2(_07252_ ), .ZN(_07253_ ) );
BUF_X4 _15278_ ( .A(_04765_ ), .Z(_07254_ ) );
INV_X1 _15279_ ( .A(_07254_ ), .ZN(_07255_ ) );
AND3_X1 _15280_ ( .A1(_07203_ ), .A2(_02730_ ), .A3(_02731_ ), .ZN(_07256_ ) );
BUF_X4 _15281_ ( .A(_07201_ ), .Z(_07257_ ) );
BUF_X4 _15282_ ( .A(_07257_ ), .Z(_07258_ ) );
AND3_X1 _15283_ ( .A1(_04108_ ), .A2(_07221_ ), .A3(_07222_ ), .ZN(_07259_ ) );
OR3_X1 _15284_ ( .A1(_07256_ ), .A2(_07258_ ), .A3(_07259_ ), .ZN(_07260_ ) );
BUF_X2 _15285_ ( .A(_04640_ ), .Z(_07261_ ) );
BUF_X2 _15286_ ( .A(_07261_ ), .Z(_07262_ ) );
NOR2_X1 _15287_ ( .A1(_07204_ ), .A2(_02855_ ), .ZN(_07263_ ) );
BUF_X4 _15288_ ( .A(_07220_ ), .Z(_07264_ ) );
BUF_X4 _15289_ ( .A(_07264_ ), .Z(_07265_ ) );
BUF_X2 _15290_ ( .A(_07221_ ), .Z(_07266_ ) );
BUF_X2 _15291_ ( .A(_07222_ ), .Z(_07267_ ) );
AOI21_X1 _15292_ ( .A(_02833_ ), .B1(_07266_ ), .B2(_07267_ ), .ZN(_07268_ ) );
OR3_X1 _15293_ ( .A1(_07263_ ), .A2(_07265_ ), .A3(_07268_ ), .ZN(_07269_ ) );
NAND3_X1 _15294_ ( .A1(_07260_ ), .A2(_07262_ ), .A3(_07269_ ), .ZN(_07270_ ) );
BUF_X4 _15295_ ( .A(_04640_ ), .Z(_07271_ ) );
BUF_X4 _15296_ ( .A(_07271_ ), .Z(_07272_ ) );
BUF_X4 _15297_ ( .A(_07272_ ), .Z(_07273_ ) );
BUF_X4 _15298_ ( .A(_07220_ ), .Z(_07274_ ) );
BUF_X2 _15299_ ( .A(_07274_ ), .Z(_07275_ ) );
AOI21_X1 _15300_ ( .A(_02779_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07276_ ) );
NOR3_X1 _15301_ ( .A1(_07275_ ), .A2(_04653_ ), .A3(_07276_ ), .ZN(_07277_ ) );
OAI21_X1 _15302_ ( .A(_07270_ ), .B1(_07273_ ), .B2(_07277_ ), .ZN(_07278_ ) );
BUF_X4 _15303_ ( .A(_07209_ ), .Z(_07279_ ) );
BUF_X4 _15304_ ( .A(_07279_ ), .Z(_07280_ ) );
NOR2_X1 _15305_ ( .A1(_07278_ ), .A2(_07280_ ), .ZN(_07281_ ) );
INV_X1 _15306_ ( .A(_07281_ ), .ZN(_07282_ ) );
BUF_X4 _15307_ ( .A(_04630_ ), .Z(_07283_ ) );
BUF_X4 _15308_ ( .A(_07283_ ), .Z(_07284_ ) );
AOI21_X1 _15309_ ( .A(_07255_ ), .B1(_07282_ ), .B2(_07284_ ), .ZN(_07285_ ) );
BUF_X4 _15310_ ( .A(_07265_ ), .Z(_07286_ ) );
AND3_X1 _15311_ ( .A1(_06742_ ), .A2(_07224_ ), .A3(_07225_ ), .ZN(_07287_ ) );
NOR3_X1 _15312_ ( .A1(_07286_ ), .A2(_07287_ ), .A3(_07231_ ), .ZN(_07288_ ) );
INV_X1 _15313_ ( .A(_02626_ ), .ZN(_07289_ ) );
AND3_X1 _15314_ ( .A1(_07289_ ), .A2(_07224_ ), .A3(_07225_ ), .ZN(_07290_ ) );
AOI21_X1 _15315_ ( .A(_02655_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07291_ ) );
BUF_X2 _15316_ ( .A(_07202_ ), .Z(_07292_ ) );
NOR3_X1 _15317_ ( .A1(_07290_ ), .A2(_07291_ ), .A3(_07292_ ), .ZN(_07293_ ) );
OAI21_X1 _15318_ ( .A(_07273_ ), .B1(_07288_ ), .B2(_07293_ ), .ZN(_07294_ ) );
AND3_X1 _15319_ ( .A1(_04685_ ), .A2(_07221_ ), .A3(_07222_ ), .ZN(_07295_ ) );
AOI21_X1 _15320_ ( .A(_03094_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07296_ ) );
OAI21_X1 _15321_ ( .A(_07286_ ), .B1(_07295_ ), .B2(_07296_ ), .ZN(_07297_ ) );
AND3_X1 _15322_ ( .A1(_04572_ ), .A2(_07224_ ), .A3(_07225_ ), .ZN(_07298_ ) );
AOI21_X1 _15323_ ( .A(_02682_ ), .B1(_07224_ ), .B2(_07225_ ), .ZN(_07299_ ) );
OAI21_X1 _15324_ ( .A(_07292_ ), .B1(_07298_ ), .B2(_07299_ ), .ZN(_07300_ ) );
BUF_X2 _15325_ ( .A(_07206_ ), .Z(_07301_ ) );
NAND3_X1 _15326_ ( .A1(_07297_ ), .A2(_07300_ ), .A3(_07301_ ), .ZN(_07302_ ) );
NAND2_X1 _15327_ ( .A1(_07294_ ), .A2(_07302_ ), .ZN(_07303_ ) );
BUF_X4 _15328_ ( .A(_07258_ ), .Z(_07304_ ) );
AOI21_X1 _15329_ ( .A(_04179_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07305_ ) );
AND3_X1 _15330_ ( .A1(_06840_ ), .A2(_07233_ ), .A3(_07234_ ), .ZN(_07306_ ) );
OAI21_X1 _15331_ ( .A(_07304_ ), .B1(_07305_ ), .B2(_07306_ ), .ZN(_07307_ ) );
INV_X1 _15332_ ( .A(_03012_ ), .ZN(_07308_ ) );
AND3_X1 _15333_ ( .A1(_07308_ ), .A2(_07215_ ), .A3(_07216_ ), .ZN(_07309_ ) );
AOI21_X1 _15334_ ( .A(_04248_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07310_ ) );
OAI21_X1 _15335_ ( .A(_07286_ ), .B1(_07309_ ), .B2(_07310_ ), .ZN(_07311_ ) );
AOI21_X1 _15336_ ( .A(_07301_ ), .B1(_07307_ ), .B2(_07311_ ), .ZN(_07312_ ) );
AOI21_X1 _15337_ ( .A(_02886_ ), .B1(_07266_ ), .B2(_07267_ ), .ZN(_07313_ ) );
INV_X1 _15338_ ( .A(_02908_ ), .ZN(_07314_ ) );
AND3_X1 _15339_ ( .A1(_07314_ ), .A2(_07266_ ), .A3(_07267_ ), .ZN(_07315_ ) );
OAI21_X1 _15340_ ( .A(_07275_ ), .B1(_07313_ ), .B2(_07315_ ), .ZN(_07316_ ) );
AND3_X1 _15341_ ( .A1(_04679_ ), .A2(_07215_ ), .A3(_07216_ ), .ZN(_07317_ ) );
AOI21_X1 _15342_ ( .A(_02963_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07318_ ) );
OAI21_X1 _15343_ ( .A(_07292_ ), .B1(_07317_ ), .B2(_07318_ ), .ZN(_07319_ ) );
AOI21_X1 _15344_ ( .A(_07262_ ), .B1(_07316_ ), .B2(_07319_ ), .ZN(_07320_ ) );
NOR2_X1 _15345_ ( .A1(_07312_ ), .A2(_07320_ ), .ZN(_07321_ ) );
BUF_X4 _15346_ ( .A(_07209_ ), .Z(_07322_ ) );
BUF_X4 _15347_ ( .A(_07322_ ), .Z(_07323_ ) );
MUX2_X1 _15348_ ( .A(_07303_ ), .B(_07321_ ), .S(_07323_ ), .Z(_07324_ ) );
OAI21_X1 _15349_ ( .A(_07285_ ), .B1(_07284_ ), .B2(_07324_ ), .ZN(_07325_ ) );
BUF_X2 _15350_ ( .A(_04506_ ), .Z(_07326_ ) );
BUF_X2 _15351_ ( .A(_07326_ ), .Z(_07327_ ) );
NAND2_X1 _15352_ ( .A1(_04546_ ), .A2(_07327_ ), .ZN(_07328_ ) );
BUF_X4 _15353_ ( .A(_04772_ ), .Z(_07329_ ) );
OAI21_X1 _15354_ ( .A(_07329_ ), .B1(_04697_ ), .B2(_02575_ ), .ZN(_07330_ ) );
AND4_X1 _15355_ ( .A1(_07253_ ), .A2(_07325_ ), .A3(_07328_ ), .A4(_07330_ ), .ZN(_07331_ ) );
NOR2_X1 _15356_ ( .A1(_04584_ ), .A2(_04297_ ), .ZN(_07332_ ) );
NOR2_X1 _15357_ ( .A1(_04579_ ), .A2(_04679_ ), .ZN(_07333_ ) );
NAND2_X1 _15358_ ( .A1(_04584_ ), .A2(_04297_ ), .ZN(_07334_ ) );
AOI21_X1 _15359_ ( .A(_07332_ ), .B1(_07333_ ), .B2(_07334_ ), .ZN(_07335_ ) );
NOR4_X1 _15360_ ( .A1(_04613_ ), .A2(_04621_ ), .A3(_04614_ ), .A4(_07335_ ), .ZN(_07336_ ) );
NOR4_X1 _15361_ ( .A1(_04613_ ), .A2(_07308_ ), .A3(_04614_ ), .A4(_04619_ ), .ZN(_07337_ ) );
NOR3_X1 _15362_ ( .A1(_07336_ ), .A2(_07337_ ), .A3(_04613_ ), .ZN(_07338_ ) );
AND2_X2 _15363_ ( .A1(_04602_ ), .A2(_04607_ ), .ZN(_07339_ ) );
AND3_X1 _15364_ ( .A1(_04593_ ), .A2(_04597_ ), .A3(_07339_ ), .ZN(_07340_ ) );
INV_X1 _15365_ ( .A(_07340_ ), .ZN(_07341_ ) );
NOR2_X1 _15366_ ( .A1(_07338_ ), .A2(_07341_ ), .ZN(_07342_ ) );
INV_X1 _15367_ ( .A(_04179_ ), .ZN(_07343_ ) );
NOR2_X1 _15368_ ( .A1(_04606_ ), .A2(_07343_ ), .ZN(_07344_ ) );
AND2_X1 _15369_ ( .A1(_04606_ ), .A2(_07343_ ), .ZN(_07345_ ) );
INV_X1 _15370_ ( .A(_07345_ ), .ZN(_07346_ ) );
NOR2_X1 _15371_ ( .A1(_04601_ ), .A2(_06840_ ), .ZN(_07347_ ) );
AOI21_X1 _15372_ ( .A(_07344_ ), .B1(_07346_ ), .B2(_07347_ ), .ZN(_07348_ ) );
INV_X1 _15373_ ( .A(_04597_ ), .ZN(_07349_ ) );
NOR4_X1 _15374_ ( .A1(_07348_ ), .A2(_04591_ ), .A3(_07349_ ), .A4(_04592_ ), .ZN(_07350_ ) );
NOR4_X1 _15375_ ( .A1(_04591_ ), .A2(_04685_ ), .A3(_04592_ ), .A4(_04596_ ), .ZN(_07351_ ) );
NOR4_X1 _15376_ ( .A1(_07342_ ), .A2(_04591_ ), .A3(_07350_ ), .A4(_07351_ ), .ZN(_07352_ ) );
INV_X1 _15377_ ( .A(_07352_ ), .ZN(_07353_ ) );
INV_X1 _15378_ ( .A(_04658_ ), .ZN(_07354_ ) );
NOR2_X1 _15379_ ( .A1(_04640_ ), .A2(_04108_ ), .ZN(_07355_ ) );
INV_X1 _15380_ ( .A(_07355_ ), .ZN(_07356_ ) );
AND3_X2 _15381_ ( .A1(_04645_ ), .A2(_02779_ ), .A3(_04646_ ), .ZN(_07357_ ) );
INV_X1 _15382_ ( .A(_07357_ ), .ZN(_07358_ ) );
NAND2_X1 _15383_ ( .A1(_04647_ ), .A2(_02805_ ), .ZN(_07359_ ) );
NOR2_X1 _15384_ ( .A1(_07132_ ), .A2(_04650_ ), .ZN(_07360_ ) );
AND3_X2 _15385_ ( .A1(_07358_ ), .A2(_07359_ ), .A3(_07360_ ), .ZN(_07361_ ) );
NOR2_X4 _15386_ ( .A1(_07361_ ), .A2(_07357_ ), .ZN(_07362_ ) );
OAI221_X1 _15387_ ( .A(_07356_ ), .B1(_02810_ ), .B2(_04643_ ), .C1(_07362_ ), .C2(_04656_ ), .ZN(_07363_ ) );
AND2_X1 _15388_ ( .A1(_04666_ ), .A2(_04670_ ), .ZN(_07364_ ) );
INV_X1 _15389_ ( .A(_04632_ ), .ZN(_07365_ ) );
AND2_X1 _15390_ ( .A1(_04625_ ), .A2(_02833_ ), .ZN(_07366_ ) );
NOR2_X1 _15391_ ( .A1(_04625_ ), .A2(_02833_ ), .ZN(_07367_ ) );
NOR3_X1 _15392_ ( .A1(_07365_ ), .A2(_07366_ ), .A3(_07367_ ), .ZN(_07368_ ) );
AND4_X2 _15393_ ( .A1(_07354_ ), .A2(_07363_ ), .A3(_07364_ ), .A4(_07368_ ), .ZN(_07369_ ) );
NOR2_X1 _15394_ ( .A1(_04665_ ), .A2(_02912_ ), .ZN(_07370_ ) );
NOR2_X1 _15395_ ( .A1(_04669_ ), .A2(_07314_ ), .ZN(_07371_ ) );
INV_X1 _15396_ ( .A(_07366_ ), .ZN(_07372_ ) );
NOR2_X1 _15397_ ( .A1(_04629_ ), .A2(_02860_ ), .ZN(_07373_ ) );
INV_X1 _15398_ ( .A(_07373_ ), .ZN(_07374_ ) );
AOI21_X1 _15399_ ( .A(_07367_ ), .B1(_07372_ ), .B2(_07374_ ), .ZN(_07375_ ) );
AOI221_X1 _15400_ ( .A(_07370_ ), .B1(_04666_ ), .B2(_07371_ ), .C1(_07375_ ), .C2(_07364_ ), .ZN(_07376_ ) );
INV_X1 _15401_ ( .A(_07376_ ), .ZN(_07377_ ) );
NOR2_X2 _15402_ ( .A1(_07369_ ), .A2(_07377_ ), .ZN(_07378_ ) );
AND2_X1 _15403_ ( .A1(_04580_ ), .A2(_04585_ ), .ZN(_07379_ ) );
AND3_X1 _15404_ ( .A1(_04615_ ), .A2(_04620_ ), .A3(_07379_ ), .ZN(_07380_ ) );
NAND2_X1 _15405_ ( .A1(_07340_ ), .A2(_07380_ ), .ZN(_07381_ ) );
NOR2_X2 _15406_ ( .A1(_07378_ ), .A2(_07381_ ), .ZN(_07382_ ) );
NOR2_X2 _15407_ ( .A1(_07353_ ), .A2(_07382_ ), .ZN(_07383_ ) );
INV_X2 _15408_ ( .A(_07383_ ), .ZN(_07384_ ) );
AND2_X1 _15409_ ( .A1(_04568_ ), .A2(_04575_ ), .ZN(_07385_ ) );
AND4_X4 _15410_ ( .A1(_04703_ ), .A2(_07384_ ), .A3(_04555_ ), .A4(_07385_ ), .ZN(_07386_ ) );
INV_X1 _15411_ ( .A(_04555_ ), .ZN(_07387_ ) );
NOR2_X1 _15412_ ( .A1(_04567_ ), .A2(_03695_ ), .ZN(_07388_ ) );
AOI21_X1 _15413_ ( .A(_07388_ ), .B1(_04568_ ), .B2(_04573_ ), .ZN(_07389_ ) );
OR3_X1 _15414_ ( .A1(_04704_ ), .A2(_07387_ ), .A3(_07389_ ), .ZN(_07390_ ) );
NOR2_X1 _15415_ ( .A1(_04554_ ), .A2(_07289_ ), .ZN(_07391_ ) );
NAND3_X1 _15416_ ( .A1(_04560_ ), .A2(_04562_ ), .A3(_07391_ ), .ZN(_07392_ ) );
AND3_X1 _15417_ ( .A1(_07390_ ), .A2(_04560_ ), .A3(_07392_ ), .ZN(_07393_ ) );
INV_X1 _15418_ ( .A(_07393_ ), .ZN(_07394_ ) );
NOR2_X1 _15419_ ( .A1(_07386_ ), .A2(_07394_ ), .ZN(_07395_ ) );
INV_X1 _15420_ ( .A(_04550_ ), .ZN(_07396_ ) );
NOR2_X1 _15421_ ( .A1(_07395_ ), .A2(_07396_ ), .ZN(_07397_ ) );
NOR2_X1 _15422_ ( .A1(_04549_ ), .A2(_06742_ ), .ZN(_07398_ ) );
OR3_X1 _15423_ ( .A1(_07397_ ), .A2(_04546_ ), .A3(_07398_ ), .ZN(_07399_ ) );
OAI21_X1 _15424_ ( .A(_04546_ ), .B1(_07397_ ), .B2(_07398_ ), .ZN(_07400_ ) );
INV_X1 _15425_ ( .A(_04770_ ), .ZN(_07401_ ) );
AOI21_X1 _15426_ ( .A(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_07402_ ) );
AND2_X2 _15427_ ( .A1(_07401_ ), .A2(_07402_ ), .ZN(_07403_ ) );
BUF_X4 _15428_ ( .A(_07403_ ), .Z(_07404_ ) );
NAND3_X1 _15429_ ( .A1(_07399_ ), .A2(_07400_ ), .A3(_07404_ ), .ZN(_07405_ ) );
AND2_X2 _15430_ ( .A1(_04770_ ), .A2(\ID_EX_typ [2] ), .ZN(_07406_ ) );
BUF_X2 _15431_ ( .A(_07406_ ), .Z(_07407_ ) );
BUF_X2 _15432_ ( .A(_07407_ ), .Z(_07408_ ) );
BUF_X4 _15433_ ( .A(_04419_ ), .Z(_07409_ ) );
AOI22_X1 _15434_ ( .A1(_07252_ ), .A2(_07408_ ), .B1(_04698_ ), .B2(_07409_ ), .ZN(_07410_ ) );
NAND3_X1 _15435_ ( .A1(_07331_ ), .A2(_07405_ ), .A3(_07410_ ), .ZN(_07411_ ) );
NOR3_X1 _15436_ ( .A1(_07124_ ), .A2(_07110_ ), .A3(_07114_ ), .ZN(_07412_ ) );
NOR2_X1 _15437_ ( .A1(_03580_ ), .A2(\ID_EX_typ [2] ), .ZN(_07413_ ) );
AND3_X1 _15438_ ( .A1(_04764_ ), .A2(_07413_ ), .A3(_04511_ ), .ZN(_07414_ ) );
AOI21_X1 _15439_ ( .A(_07414_ ), .B1(\ID_EX_typ [4] ), .B2(_07123_ ), .ZN(_07415_ ) );
AND2_X1 _15440_ ( .A1(_07412_ ), .A2(_07415_ ), .ZN(_07416_ ) );
AND2_X2 _15441_ ( .A1(_02413_ ), .A2(_02406_ ), .ZN(_07417_ ) );
INV_X2 _15442_ ( .A(_07417_ ), .ZN(_07418_ ) );
NOR2_X1 _15443_ ( .A1(_07416_ ), .A2(_07418_ ), .ZN(_07419_ ) );
INV_X1 _15444_ ( .A(_07419_ ), .ZN(_07420_ ) );
BUF_X4 _15445_ ( .A(_07420_ ), .Z(_07421_ ) );
AOI21_X1 _15446_ ( .A(_07128_ ), .B1(_07411_ ), .B2(_07421_ ), .ZN(_07422_ ) );
OAI21_X1 _15447_ ( .A(_06994_ ), .B1(_05624_ ), .B2(_05663_ ), .ZN(_07423_ ) );
OAI21_X1 _15448_ ( .A(_07107_ ), .B1(_07422_ ), .B2(_07423_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
BUF_X4 _15449_ ( .A(_03341_ ), .Z(_07424_ ) );
OAI21_X1 _15450_ ( .A(_07424_ ), .B1(_04850_ ), .B2(_04851_ ), .ZN(_07425_ ) );
OAI21_X1 _15451_ ( .A(_07125_ ), .B1(_07118_ ), .B2(_07119_ ), .ZN(_07426_ ) );
AOI21_X1 _15452_ ( .A(_07426_ ), .B1(_07119_ ), .B2(_07118_ ), .ZN(_07427_ ) );
BUF_X2 _15453_ ( .A(_07110_ ), .Z(_07428_ ) );
NAND2_X1 _15454_ ( .A1(_04857_ ), .A2(_07428_ ), .ZN(_07429_ ) );
OAI21_X1 _15455_ ( .A(_07429_ ), .B1(_02599_ ), .B2(_07115_ ), .ZN(_07430_ ) );
OAI21_X1 _15456_ ( .A(_07417_ ), .B1(_07427_ ), .B2(_07430_ ), .ZN(_07431_ ) );
NAND2_X1 _15457_ ( .A1(_07431_ ), .A2(_04831_ ), .ZN(_07432_ ) );
BUF_X2 _15458_ ( .A(_07261_ ), .Z(_07433_ ) );
OAI21_X1 _15459_ ( .A(_07433_ ), .B1(_07286_ ), .B2(_07242_ ), .ZN(_07434_ ) );
NAND3_X1 _15460_ ( .A1(_07186_ ), .A2(_07434_ ), .A3(_07212_ ), .ZN(_07435_ ) );
AOI211_X1 _15461_ ( .A(_07138_ ), .B(_07188_ ), .C1(_07435_ ), .C2(_07187_ ), .ZN(_07436_ ) );
NOR2_X1 _15462_ ( .A1(_07203_ ), .A2(_02548_ ), .ZN(_07437_ ) );
AOI21_X1 _15463_ ( .A(_02522_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07438_ ) );
NOR3_X1 _15464_ ( .A1(_07437_ ), .A2(_07438_ ), .A3(_07229_ ), .ZN(_07439_ ) );
NOR2_X1 _15465_ ( .A1(_07203_ ), .A2(_02575_ ), .ZN(_07440_ ) );
AOI21_X1 _15466_ ( .A(_02598_ ), .B1(_07224_ ), .B2(_07225_ ), .ZN(_07441_ ) );
NOR3_X1 _15467_ ( .A1(_07440_ ), .A2(_07220_ ), .A3(_07441_ ), .ZN(_07442_ ) );
OAI21_X1 _15468_ ( .A(_07271_ ), .B1(_07439_ ), .B2(_07442_ ), .ZN(_07443_ ) );
BUF_X4 _15469_ ( .A(_04641_ ), .Z(_07444_ ) );
AND3_X1 _15470_ ( .A1(_04488_ ), .A2(_07215_ ), .A3(_07216_ ), .ZN(_07445_ ) );
AOI21_X1 _15471_ ( .A(_03172_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07446_ ) );
NOR3_X1 _15472_ ( .A1(_07264_ ), .A2(_07445_ ), .A3(_07446_ ), .ZN(_07447_ ) );
NOR2_X1 _15473_ ( .A1(_07203_ ), .A2(_03987_ ), .ZN(_07448_ ) );
AOI21_X1 _15474_ ( .A(_03221_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07449_ ) );
NOR3_X1 _15475_ ( .A1(_07448_ ), .A2(_07229_ ), .A3(_07449_ ), .ZN(_07450_ ) );
OAI21_X1 _15476_ ( .A(_07444_ ), .B1(_07447_ ), .B2(_07450_ ), .ZN(_07451_ ) );
NAND2_X1 _15477_ ( .A1(_07443_ ), .A2(_07451_ ), .ZN(_07452_ ) );
AND3_X1 _15478_ ( .A1(_07203_ ), .A2(_03251_ ), .A3(_03252_ ), .ZN(_07453_ ) );
AND3_X1 _15479_ ( .A1(_03282_ ), .A2(_07224_ ), .A3(_07225_ ), .ZN(_07454_ ) );
NOR2_X1 _15480_ ( .A1(_07453_ ), .A2(_07454_ ), .ZN(_07455_ ) );
INV_X1 _15481_ ( .A(_03310_ ), .ZN(_07456_ ) );
MUX2_X1 _15482_ ( .A(_03337_ ), .B(_07456_ ), .S(_07203_ ), .Z(_07457_ ) );
MUX2_X1 _15483_ ( .A(_07455_ ), .B(_07457_ ), .S(_07264_ ), .Z(_07458_ ) );
AND2_X1 _15484_ ( .A1(_07458_ ), .A2(_07261_ ), .ZN(_07459_ ) );
MUX2_X1 _15485_ ( .A(_07452_ ), .B(_07459_ ), .S(_07209_ ), .Z(_07460_ ) );
BUF_X2 _15486_ ( .A(_07249_ ), .Z(_07461_ ) );
AND2_X1 _15487_ ( .A1(_07460_ ), .A2(_07461_ ), .ZN(_07462_ ) );
OAI21_X1 _15488_ ( .A(_07130_ ), .B1(_07436_ ), .B2(_07462_ ), .ZN(_07463_ ) );
BUF_X2 _15489_ ( .A(_07250_ ), .Z(_07464_ ) );
NAND3_X1 _15490_ ( .A1(_07460_ ), .A2(_07464_ ), .A3(_07407_ ), .ZN(_07465_ ) );
NAND2_X1 _15491_ ( .A1(_07463_ ), .A2(_07465_ ), .ZN(_07466_ ) );
NOR2_X1 _15492_ ( .A1(_07204_ ), .A2(_02886_ ), .ZN(_07467_ ) );
AOI21_X1 _15493_ ( .A(_02938_ ), .B1(_07266_ ), .B2(_07267_ ), .ZN(_07468_ ) );
NOR3_X1 _15494_ ( .A1(_07467_ ), .A2(_07265_ ), .A3(_07468_ ), .ZN(_07469_ ) );
AND3_X1 _15495_ ( .A1(_04450_ ), .A2(_07221_ ), .A3(_07222_ ), .ZN(_07470_ ) );
AOI21_X1 _15496_ ( .A(_02908_ ), .B1(_07221_ ), .B2(_07222_ ), .ZN(_07471_ ) );
BUF_X2 _15497_ ( .A(_07229_ ), .Z(_07472_ ) );
NOR3_X1 _15498_ ( .A1(_07470_ ), .A2(_07471_ ), .A3(_07472_ ), .ZN(_07473_ ) );
NOR2_X1 _15499_ ( .A1(_07469_ ), .A2(_07473_ ), .ZN(_07474_ ) );
NOR2_X1 _15500_ ( .A1(_07474_ ), .A2(_07433_ ), .ZN(_07475_ ) );
BUF_X4 _15501_ ( .A(_04643_ ), .Z(_07476_ ) );
BUF_X2 _15502_ ( .A(_07476_ ), .Z(_07477_ ) );
BUF_X2 _15503_ ( .A(_07444_ ), .Z(_07478_ ) );
AND3_X1 _15504_ ( .A1(_04297_ ), .A2(_07266_ ), .A3(_07267_ ), .ZN(_07479_ ) );
AOI21_X1 _15505_ ( .A(_03012_ ), .B1(_07266_ ), .B2(_07267_ ), .ZN(_07480_ ) );
OR3_X1 _15506_ ( .A1(_07479_ ), .A2(_07480_ ), .A3(_07202_ ), .ZN(_07481_ ) );
AOI21_X1 _15507_ ( .A(_03070_ ), .B1(_07266_ ), .B2(_07267_ ), .ZN(_07482_ ) );
INV_X1 _15508_ ( .A(_07482_ ), .ZN(_07483_ ) );
OAI211_X1 _15509_ ( .A(_07483_ ), .B(_07258_ ), .C1(_04248_ ), .C2(_07204_ ), .ZN(_07484_ ) );
AOI21_X1 _15510_ ( .A(_07478_ ), .B1(_07481_ ), .B2(_07484_ ), .ZN(_07485_ ) );
OR3_X1 _15511_ ( .A1(_07475_ ), .A2(_07477_ ), .A3(_07485_ ), .ZN(_07486_ ) );
AND3_X1 _15512_ ( .A1(_04154_ ), .A2(_07266_ ), .A3(_07267_ ), .ZN(_07487_ ) );
AOI21_X1 _15513_ ( .A(_02706_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07488_ ) );
OR3_X1 _15514_ ( .A1(_07275_ ), .A2(_07487_ ), .A3(_07488_ ), .ZN(_07489_ ) );
NOR2_X1 _15515_ ( .A1(_07204_ ), .A2(_04179_ ), .ZN(_07490_ ) );
AOI21_X1 _15516_ ( .A(_03118_ ), .B1(_07266_ ), .B2(_07267_ ), .ZN(_07491_ ) );
OR3_X1 _15517_ ( .A1(_07490_ ), .A2(_07472_ ), .A3(_07491_ ), .ZN(_07492_ ) );
NAND3_X1 _15518_ ( .A1(_07489_ ), .A2(_07492_ ), .A3(_07301_ ), .ZN(_07493_ ) );
AND3_X1 _15519_ ( .A1(_03695_ ), .A2(_07224_ ), .A3(_07225_ ), .ZN(_07494_ ) );
AOI21_X1 _15520_ ( .A(_02626_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07495_ ) );
OAI21_X1 _15521_ ( .A(_07275_ ), .B1(_07494_ ), .B2(_07495_ ), .ZN(_07496_ ) );
AND3_X1 _15522_ ( .A1(_03656_ ), .A2(_07215_ ), .A3(_07216_ ), .ZN(_07497_ ) );
OAI21_X1 _15523_ ( .A(_07258_ ), .B1(_07497_ ), .B2(_07441_ ), .ZN(_07498_ ) );
NAND2_X1 _15524_ ( .A1(_07496_ ), .A2(_07498_ ), .ZN(_07499_ ) );
NAND2_X1 _15525_ ( .A1(_07499_ ), .A2(_07262_ ), .ZN(_07500_ ) );
AND2_X1 _15526_ ( .A1(_07493_ ), .A2(_07500_ ), .ZN(_07501_ ) );
OAI211_X1 _15527_ ( .A(_07486_ ), .B(_07251_ ), .C1(_07280_ ), .C2(_07501_ ), .ZN(_07502_ ) );
AOI21_X1 _15528_ ( .A(_04650_ ), .B1(_07233_ ), .B2(_07234_ ), .ZN(_07503_ ) );
AND2_X1 _15529_ ( .A1(_07503_ ), .A2(_07472_ ), .ZN(_07504_ ) );
INV_X1 _15530_ ( .A(_07504_ ), .ZN(_07505_ ) );
NOR2_X1 _15531_ ( .A1(_02732_ ), .A2(_07203_ ), .ZN(_07506_ ) );
AOI21_X1 _15532_ ( .A(_02855_ ), .B1(_07224_ ), .B2(_07225_ ), .ZN(_07507_ ) );
OAI21_X1 _15533_ ( .A(_07472_ ), .B1(_07506_ ), .B2(_07507_ ), .ZN(_07508_ ) );
AND3_X1 _15534_ ( .A1(_02805_ ), .A2(_07221_ ), .A3(_07222_ ), .ZN(_07509_ ) );
AOI21_X1 _15535_ ( .A(_02755_ ), .B1(_07224_ ), .B2(_07225_ ), .ZN(_07510_ ) );
OAI21_X1 _15536_ ( .A(_07265_ ), .B1(_07509_ ), .B2(_07510_ ), .ZN(_07511_ ) );
NAND2_X1 _15537_ ( .A1(_07508_ ), .A2(_07511_ ), .ZN(_07512_ ) );
MUX2_X1 _15538_ ( .A(_07505_ ), .B(_07512_ ), .S(_07272_ ), .Z(_07513_ ) );
BUF_X2 _15539_ ( .A(_07209_ ), .Z(_07514_ ) );
OR3_X1 _15540_ ( .A1(_07513_ ), .A2(_07250_ ), .A3(_07514_ ), .ZN(_07515_ ) );
AOI21_X1 _15541_ ( .A(_07255_ ), .B1(_07502_ ), .B2(_07515_ ), .ZN(_07516_ ) );
OR2_X1 _15542_ ( .A1(_07466_ ), .A2(_07516_ ), .ZN(_07517_ ) );
OAI21_X1 _15543_ ( .A(_07403_ ), .B1(_07395_ ), .B2(_07396_ ), .ZN(_07518_ ) );
AOI21_X1 _15544_ ( .A(_07518_ ), .B1(_07396_ ), .B2(_07395_ ), .ZN(_07519_ ) );
AND2_X1 _15545_ ( .A1(_04550_ ), .A2(_07326_ ), .ZN(_07520_ ) );
BUF_X4 _15546_ ( .A(_04420_ ), .Z(_07521_ ) );
NOR3_X1 _15547_ ( .A1(_04549_ ), .A2(_06742_ ), .A3(_07521_ ), .ZN(_07522_ ) );
INV_X1 _15548_ ( .A(_07329_ ), .ZN(_07523_ ) );
BUF_X2 _15549_ ( .A(_07523_ ), .Z(_07524_ ) );
AOI21_X1 _15550_ ( .A(_07524_ ), .B1(_04549_ ), .B2(_06742_ ), .ZN(_07525_ ) );
OR3_X1 _15551_ ( .A1(_07520_ ), .A2(_07522_ ), .A3(_07525_ ), .ZN(_07526_ ) );
OR3_X1 _15552_ ( .A1(_07517_ ), .A2(_07519_ ), .A3(_07526_ ), .ZN(_07527_ ) );
AOI21_X1 _15553_ ( .A(_07432_ ), .B1(_07527_ ), .B2(_07421_ ), .ZN(_07528_ ) );
OAI21_X1 _15554_ ( .A(_06994_ ), .B1(_04856_ ), .B2(_05663_ ), .ZN(_07529_ ) );
OAI21_X1 _15555_ ( .A(_07425_ ), .B1(_07528_ ), .B2(_07529_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OR2_X1 _15556_ ( .A1(_04916_ ), .A2(_06700_ ), .ZN(_07530_ ) );
BUF_X4 _15557_ ( .A(_07418_ ), .Z(_07531_ ) );
AND2_X1 _15558_ ( .A1(_03692_ ), .A2(_02626_ ), .ZN(_07532_ ) );
NAND2_X1 _15559_ ( .A1(_04457_ ), .A2(_03747_ ), .ZN(_07533_ ) );
AND2_X1 _15560_ ( .A1(_07533_ ), .A2(_04465_ ), .ZN(_07534_ ) );
OAI21_X1 _15561_ ( .A(_04464_ ), .B1(_07534_ ), .B2(_04462_ ), .ZN(_07535_ ) );
AOI21_X1 _15562_ ( .A(_07532_ ), .B1(_07535_ ), .B2(_03693_ ), .ZN(_07536_ ) );
XNOR2_X1 _15563_ ( .A(_07536_ ), .B(_03657_ ), .ZN(_07537_ ) );
NAND2_X1 _15564_ ( .A1(_07537_ ), .A2(_07126_ ), .ZN(_07538_ ) );
BUF_X4 _15565_ ( .A(_07114_ ), .Z(_07539_ ) );
AOI22_X1 _15566_ ( .A1(_04884_ ), .A2(_07428_ ), .B1(\ID_EX_imm [19] ), .B2(_07539_ ), .ZN(_07540_ ) );
AOI21_X1 _15567_ ( .A(_07531_ ), .B1(_07538_ ), .B2(_07540_ ), .ZN(_07541_ ) );
OR2_X1 _15568_ ( .A1(_07541_ ), .A2(_05180_ ), .ZN(_07542_ ) );
XNOR2_X1 _15569_ ( .A(_07133_ ), .B(_04640_ ), .ZN(_07543_ ) );
BUF_X2 _15570_ ( .A(_07212_ ), .Z(_07544_ ) );
NAND3_X1 _15571_ ( .A1(_07200_ ), .A2(_07543_ ), .A3(_07544_ ), .ZN(_07545_ ) );
AOI211_X1 _15572_ ( .A(_07138_ ), .B(_07188_ ), .C1(_07187_ ), .C2(_07545_ ), .ZN(_07546_ ) );
OAI21_X1 _15573_ ( .A(_07274_ ), .B1(_07230_ ), .B2(_07231_ ), .ZN(_07547_ ) );
OAI21_X1 _15574_ ( .A(_07202_ ), .B1(_07287_ ), .B2(_07291_ ), .ZN(_07548_ ) );
AOI21_X1 _15575_ ( .A(_07444_ ), .B1(_07547_ ), .B2(_07548_ ), .ZN(_07549_ ) );
OAI21_X1 _15576_ ( .A(_07257_ ), .B1(_07235_ ), .B2(_07236_ ), .ZN(_07550_ ) );
OAI21_X1 _15577_ ( .A(_07264_ ), .B1(_07223_ ), .B2(_07226_ ), .ZN(_07551_ ) );
AOI21_X1 _15578_ ( .A(_07271_ ), .B1(_07550_ ), .B2(_07551_ ), .ZN(_07552_ ) );
NOR2_X1 _15579_ ( .A1(_07549_ ), .A2(_07552_ ), .ZN(_07553_ ) );
OAI21_X1 _15580_ ( .A(_07264_ ), .B1(_07243_ ), .B2(_07244_ ), .ZN(_07554_ ) );
OAI21_X1 _15581_ ( .A(_07229_ ), .B1(_07217_ ), .B2(_07218_ ), .ZN(_07555_ ) );
NAND3_X1 _15582_ ( .A1(_07554_ ), .A2(_07271_ ), .A3(_07555_ ), .ZN(_07556_ ) );
NAND3_X1 _15583_ ( .A1(_07240_ ), .A2(_07444_ ), .A3(_07472_ ), .ZN(_07557_ ) );
NAND2_X1 _15584_ ( .A1(_07556_ ), .A2(_07557_ ), .ZN(_07558_ ) );
MUX2_X1 _15585_ ( .A(_07553_ ), .B(_07558_ ), .S(_07209_ ), .Z(_07559_ ) );
BUF_X2 _15586_ ( .A(_07461_ ), .Z(_07560_ ) );
AND2_X1 _15587_ ( .A1(_07559_ ), .A2(_07560_ ), .ZN(_07561_ ) );
OAI21_X1 _15588_ ( .A(_07131_ ), .B1(_07546_ ), .B2(_07561_ ), .ZN(_07562_ ) );
OAI21_X1 _15589_ ( .A(_07385_ ), .B1(_07353_ ), .B2(_07382_ ), .ZN(_07563_ ) );
AND2_X1 _15590_ ( .A1(_07563_ ), .A2(_07389_ ), .ZN(_07564_ ) );
OR2_X1 _15591_ ( .A1(_07564_ ), .A2(_07387_ ), .ZN(_07565_ ) );
INV_X1 _15592_ ( .A(_07391_ ), .ZN(_07566_ ) );
AND3_X1 _15593_ ( .A1(_07565_ ), .A2(_04703_ ), .A3(_07566_ ), .ZN(_07567_ ) );
AOI21_X1 _15594_ ( .A(_04703_ ), .B1(_07565_ ), .B2(_07566_ ), .ZN(_07568_ ) );
OAI21_X1 _15595_ ( .A(_07404_ ), .B1(_07567_ ), .B2(_07568_ ), .ZN(_07569_ ) );
NOR3_X1 _15596_ ( .A1(_07313_ ), .A2(_07264_ ), .A3(_07315_ ), .ZN(_07570_ ) );
NOR3_X1 _15597_ ( .A1(_07263_ ), .A2(_07257_ ), .A3(_07268_ ), .ZN(_07571_ ) );
NOR2_X1 _15598_ ( .A1(_07570_ ), .A2(_07571_ ), .ZN(_07572_ ) );
NAND2_X1 _15599_ ( .A1(_07572_ ), .A2(_07206_ ), .ZN(_07573_ ) );
NOR3_X1 _15600_ ( .A1(_07264_ ), .A2(_07309_ ), .A3(_07310_ ), .ZN(_07574_ ) );
NOR3_X1 _15601_ ( .A1(_07317_ ), .A2(_07318_ ), .A3(_07229_ ), .ZN(_07575_ ) );
OR3_X1 _15602_ ( .A1(_07574_ ), .A2(_07575_ ), .A3(_04641_ ), .ZN(_07576_ ) );
AOI21_X1 _15603_ ( .A(_07476_ ), .B1(_07573_ ), .B2(_07576_ ), .ZN(_07577_ ) );
BUF_X4 _15604_ ( .A(_07476_ ), .Z(_07578_ ) );
NOR3_X1 _15605_ ( .A1(_07274_ ), .A2(_07290_ ), .A3(_07291_ ), .ZN(_07579_ ) );
NOR3_X1 _15606_ ( .A1(_07298_ ), .A2(_07299_ ), .A3(_07257_ ), .ZN(_07580_ ) );
NOR2_X1 _15607_ ( .A1(_07579_ ), .A2(_07580_ ), .ZN(_07581_ ) );
NOR3_X1 _15608_ ( .A1(_07305_ ), .A2(_07306_ ), .A3(_07257_ ), .ZN(_07582_ ) );
NOR3_X1 _15609_ ( .A1(_07264_ ), .A2(_07295_ ), .A3(_07296_ ), .ZN(_07583_ ) );
NOR2_X1 _15610_ ( .A1(_07582_ ), .A2(_07583_ ), .ZN(_07584_ ) );
MUX2_X1 _15611_ ( .A(_07581_ ), .B(_07584_ ), .S(_07444_ ), .Z(_07585_ ) );
AOI211_X1 _15612_ ( .A(_07283_ ), .B(_07577_ ), .C1(_07578_ ), .C2(_07585_ ), .ZN(_07586_ ) );
OR3_X1 _15613_ ( .A1(_07256_ ), .A2(_07220_ ), .A3(_07259_ ), .ZN(_07587_ ) );
OR3_X1 _15614_ ( .A1(_04653_ ), .A2(_07276_ ), .A3(_07201_ ), .ZN(_07588_ ) );
AOI21_X1 _15615_ ( .A(_07206_ ), .B1(_07587_ ), .B2(_07588_ ), .ZN(_07589_ ) );
AND3_X1 _15616_ ( .A1(_07589_ ), .A2(_04630_ ), .A3(_07477_ ), .ZN(_07590_ ) );
OAI21_X1 _15617_ ( .A(_07254_ ), .B1(_07586_ ), .B2(_07590_ ), .ZN(_07591_ ) );
NAND3_X1 _15618_ ( .A1(_07559_ ), .A2(_07461_ ), .A3(_07406_ ), .ZN(_07592_ ) );
OAI211_X1 _15619_ ( .A(_07591_ ), .B(_07592_ ), .C1(_04561_ ), .C2(_07524_ ), .ZN(_07593_ ) );
AOI221_X4 _15620_ ( .A(_07593_ ), .B1(_04559_ ), .B2(_04419_ ), .C1(_04703_ ), .C2(_07327_ ), .ZN(_07594_ ) );
NAND3_X1 _15621_ ( .A1(_07562_ ), .A2(_07569_ ), .A3(_07594_ ), .ZN(_07595_ ) );
AOI21_X1 _15622_ ( .A(_07542_ ), .B1(_07595_ ), .B2(_07421_ ), .ZN(_07596_ ) );
OAI21_X1 _15623_ ( .A(_06994_ ), .B1(_04877_ ), .B2(_05663_ ), .ZN(_07597_ ) );
OAI21_X1 _15624_ ( .A(_07530_ ), .B1(_07596_ ), .B2(_07597_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
OAI21_X1 _15625_ ( .A(_07424_ ), .B1(_04960_ ), .B2(_04961_ ), .ZN(_07598_ ) );
INV_X1 _15626_ ( .A(_07124_ ), .ZN(_07599_ ) );
BUF_X2 _15627_ ( .A(_07599_ ), .Z(_07600_ ) );
AOI21_X1 _15628_ ( .A(_07600_ ), .B1(_07535_ ), .B2(_03693_ ), .ZN(_07601_ ) );
OAI21_X1 _15629_ ( .A(_07601_ ), .B1(_03693_ ), .B2(_07535_ ), .ZN(_07602_ ) );
BUF_X4 _15630_ ( .A(_07110_ ), .Z(_07603_ ) );
AOI22_X1 _15631_ ( .A1(_04930_ ), .A2(_07603_ ), .B1(\ID_EX_imm [18] ), .B2(_07539_ ), .ZN(_07604_ ) );
AOI21_X1 _15632_ ( .A(_07531_ ), .B1(_07602_ ), .B2(_07604_ ), .ZN(_07605_ ) );
OR2_X1 _15633_ ( .A1(_07605_ ), .A2(_05180_ ), .ZN(_07606_ ) );
NOR2_X1 _15634_ ( .A1(_07188_ ), .A2(_07138_ ), .ZN(_07607_ ) );
INV_X1 _15635_ ( .A(_07607_ ), .ZN(_07608_ ) );
NOR2_X1 _15636_ ( .A1(_07275_ ), .A2(_07204_ ), .ZN(_07609_ ) );
INV_X1 _15637_ ( .A(_07609_ ), .ZN(_07610_ ) );
AND3_X1 _15638_ ( .A1(_07186_ ), .A2(_07610_ ), .A3(_07543_ ), .ZN(_07611_ ) );
NAND2_X1 _15639_ ( .A1(_07611_ ), .A2(_07544_ ), .ZN(_07612_ ) );
AOI21_X1 _15640_ ( .A(_07608_ ), .B1(_07612_ ), .B2(_07187_ ), .ZN(_07613_ ) );
OAI21_X1 _15641_ ( .A(_07472_ ), .B1(_07437_ ), .B2(_07438_ ), .ZN(_07614_ ) );
OAI21_X1 _15642_ ( .A(_07274_ ), .B1(_07445_ ), .B2(_07446_ ), .ZN(_07615_ ) );
AOI21_X1 _15643_ ( .A(_07261_ ), .B1(_07614_ ), .B2(_07615_ ), .ZN(_07616_ ) );
OAI21_X1 _15644_ ( .A(_07274_ ), .B1(_07440_ ), .B2(_07441_ ), .ZN(_07617_ ) );
OAI21_X1 _15645_ ( .A(_07202_ ), .B1(_07497_ ), .B2(_07495_ ), .ZN(_07618_ ) );
AOI21_X1 _15646_ ( .A(_07444_ ), .B1(_07617_ ), .B2(_07618_ ), .ZN(_07619_ ) );
NOR2_X1 _15647_ ( .A1(_07616_ ), .A2(_07619_ ), .ZN(_07620_ ) );
NOR2_X1 _15648_ ( .A1(_07620_ ), .A2(_07322_ ), .ZN(_07621_ ) );
NOR3_X1 _15649_ ( .A1(_07453_ ), .A2(_07229_ ), .A3(_07454_ ), .ZN(_07622_ ) );
NOR3_X1 _15650_ ( .A1(_07448_ ), .A2(_07264_ ), .A3(_07449_ ), .ZN(_07623_ ) );
OR3_X1 _15651_ ( .A1(_07622_ ), .A2(_07623_ ), .A3(_04641_ ), .ZN(_07624_ ) );
AND2_X1 _15652_ ( .A1(_07457_ ), .A2(_07472_ ), .ZN(_07625_ ) );
OAI21_X1 _15653_ ( .A(_07624_ ), .B1(_07625_ ), .B2(_07272_ ), .ZN(_07626_ ) );
AOI21_X1 _15654_ ( .A(_07621_ ), .B1(_07626_ ), .B2(_07514_ ), .ZN(_07627_ ) );
AND2_X1 _15655_ ( .A1(_07627_ ), .A2(_07464_ ), .ZN(_07628_ ) );
OAI21_X1 _15656_ ( .A(_07131_ ), .B1(_07613_ ), .B2(_07628_ ), .ZN(_07629_ ) );
BUF_X2 _15657_ ( .A(_07476_ ), .Z(_07630_ ) );
NOR3_X1 _15658_ ( .A1(_07506_ ), .A2(_07201_ ), .A3(_07507_ ), .ZN(_07631_ ) );
NOR3_X1 _15659_ ( .A1(_07220_ ), .A2(_07470_ ), .A3(_07471_ ), .ZN(_07632_ ) );
OR3_X1 _15660_ ( .A1(_07631_ ), .A2(_07632_ ), .A3(_07433_ ), .ZN(_07633_ ) );
NOR3_X1 _15661_ ( .A1(_07274_ ), .A2(_07479_ ), .A3(_07480_ ), .ZN(_07634_ ) );
NOR3_X1 _15662_ ( .A1(_07467_ ), .A2(_07257_ ), .A3(_07468_ ), .ZN(_07635_ ) );
OR3_X1 _15663_ ( .A1(_07634_ ), .A2(_07635_ ), .A3(_07478_ ), .ZN(_07636_ ) );
AOI21_X1 _15664_ ( .A(_07630_ ), .B1(_07633_ ), .B2(_07636_ ), .ZN(_07637_ ) );
BUF_X2 _15665_ ( .A(_07578_ ), .Z(_07638_ ) );
NOR3_X1 _15666_ ( .A1(_07490_ ), .A2(_07274_ ), .A3(_07491_ ), .ZN(_07639_ ) );
AND3_X1 _15667_ ( .A1(_04249_ ), .A2(_07266_ ), .A3(_07267_ ), .ZN(_07640_ ) );
NOR3_X1 _15668_ ( .A1(_07640_ ), .A2(_07482_ ), .A3(_07257_ ), .ZN(_07641_ ) );
OAI21_X1 _15669_ ( .A(_07301_ ), .B1(_07639_ ), .B2(_07641_ ), .ZN(_07642_ ) );
NOR3_X1 _15670_ ( .A1(_07275_ ), .A2(_07494_ ), .A3(_07495_ ), .ZN(_07643_ ) );
NOR3_X1 _15671_ ( .A1(_07487_ ), .A2(_07488_ ), .A3(_07258_ ), .ZN(_07644_ ) );
OAI21_X1 _15672_ ( .A(_07262_ ), .B1(_07643_ ), .B2(_07644_ ), .ZN(_07645_ ) );
AND2_X1 _15673_ ( .A1(_07642_ ), .A2(_07645_ ), .ZN(_07646_ ) );
AOI211_X1 _15674_ ( .A(_07284_ ), .B(_07637_ ), .C1(_07638_ ), .C2(_07646_ ), .ZN(_07647_ ) );
OAI21_X1 _15675_ ( .A(_07201_ ), .B1(_07509_ ), .B2(_07510_ ), .ZN(_07648_ ) );
OAI21_X1 _15676_ ( .A(_07648_ ), .B1(_07229_ ), .B2(_07503_ ), .ZN(_07649_ ) );
BUF_X2 _15677_ ( .A(_07478_ ), .Z(_07650_ ) );
NOR4_X1 _15678_ ( .A1(_07649_ ), .A2(_07464_ ), .A3(_07280_ ), .A4(_07650_ ), .ZN(_07651_ ) );
OAI21_X1 _15679_ ( .A(_07254_ ), .B1(_07647_ ), .B2(_07651_ ), .ZN(_07652_ ) );
AOI22_X1 _15680_ ( .A1(_04555_ ), .A2(_07327_ ), .B1(_07391_ ), .B2(_07409_ ), .ZN(_07653_ ) );
AND3_X1 _15681_ ( .A1(_07629_ ), .A2(_07652_ ), .A3(_07653_ ), .ZN(_07654_ ) );
NAND3_X1 _15682_ ( .A1(_07563_ ), .A2(_07387_ ), .A3(_07389_ ), .ZN(_07655_ ) );
NAND3_X1 _15683_ ( .A1(_07565_ ), .A2(_07404_ ), .A3(_07655_ ), .ZN(_07656_ ) );
BUF_X2 _15684_ ( .A(_07523_ ), .Z(_07657_ ) );
AOI21_X1 _15685_ ( .A(_07657_ ), .B1(_04554_ ), .B2(_07289_ ), .ZN(_07658_ ) );
AOI21_X1 _15686_ ( .A(_07658_ ), .B1(_07628_ ), .B2(_07408_ ), .ZN(_07659_ ) );
NAND3_X1 _15687_ ( .A1(_07654_ ), .A2(_07656_ ), .A3(_07659_ ), .ZN(_07660_ ) );
AOI21_X1 _15688_ ( .A(_07606_ ), .B1(_07660_ ), .B2(_07421_ ), .ZN(_07661_ ) );
CLKBUF_X2 _15689_ ( .A(_02415_ ), .Z(_07662_ ) );
BUF_X4 _15690_ ( .A(_07662_ ), .Z(_07663_ ) );
NAND2_X1 _15691_ ( .A1(_04927_ ), .A2(_07663_ ), .ZN(_07664_ ) );
BUF_X4 _15692_ ( .A(_06694_ ), .Z(_07665_ ) );
NAND2_X1 _15693_ ( .A1(_07664_ ), .A2(_07665_ ), .ZN(_07666_ ) );
OAI21_X1 _15694_ ( .A(_07598_ ), .B1(_07661_ ), .B2(_07666_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
OAI21_X1 _15695_ ( .A(_07424_ ), .B1(_04997_ ), .B2(_04999_ ), .ZN(_07667_ ) );
XNOR2_X1 _15696_ ( .A(_07534_ ), .B(_03722_ ), .ZN(_07668_ ) );
NAND2_X1 _15697_ ( .A1(_07668_ ), .A2(_07126_ ), .ZN(_07669_ ) );
AOI22_X1 _15698_ ( .A1(_04981_ ), .A2(_07603_ ), .B1(\ID_EX_imm [17] ), .B2(_07539_ ), .ZN(_07670_ ) );
AOI21_X1 _15699_ ( .A(_07531_ ), .B1(_07669_ ), .B2(_07670_ ), .ZN(_07671_ ) );
OR2_X1 _15700_ ( .A1(_07671_ ), .A2(_05180_ ), .ZN(_07672_ ) );
AND3_X1 _15701_ ( .A1(_07186_ ), .A2(_07543_ ), .A3(_07212_ ), .ZN(_07673_ ) );
NAND2_X1 _15702_ ( .A1(_07673_ ), .A2(_07205_ ), .ZN(_07674_ ) );
AOI21_X1 _15703_ ( .A(_07608_ ), .B1(_07674_ ), .B2(_07187_ ), .ZN(_07675_ ) );
NAND3_X1 _15704_ ( .A1(_07232_ ), .A2(_07237_ ), .A3(_07206_ ), .ZN(_07676_ ) );
OAI21_X1 _15705_ ( .A(_07220_ ), .B1(_07287_ ), .B2(_07291_ ), .ZN(_07677_ ) );
OAI21_X1 _15706_ ( .A(_07229_ ), .B1(_07290_ ), .B2(_07299_ ), .ZN(_07678_ ) );
NAND3_X1 _15707_ ( .A1(_07677_ ), .A2(_07678_ ), .A3(_07261_ ), .ZN(_07679_ ) );
NAND2_X1 _15708_ ( .A1(_07676_ ), .A2(_07679_ ), .ZN(_07680_ ) );
NAND2_X1 _15709_ ( .A1(_07680_ ), .A2(_07578_ ), .ZN(_07681_ ) );
NAND2_X1 _15710_ ( .A1(_07246_ ), .A2(_07478_ ), .ZN(_07682_ ) );
OR3_X1 _15711_ ( .A1(_07219_ ), .A2(_07444_ ), .A3(_07227_ ), .ZN(_07683_ ) );
NAND2_X1 _15712_ ( .A1(_07682_ ), .A2(_07683_ ), .ZN(_07684_ ) );
OAI21_X1 _15713_ ( .A(_07681_ ), .B1(_07684_ ), .B2(_07630_ ), .ZN(_07685_ ) );
AND2_X1 _15714_ ( .A1(_07685_ ), .A2(_07251_ ), .ZN(_07686_ ) );
OAI21_X1 _15715_ ( .A(_07131_ ), .B1(_07675_ ), .B2(_07686_ ), .ZN(_07687_ ) );
BUF_X2 _15716_ ( .A(_07283_ ), .Z(_07688_ ) );
AOI21_X1 _15717_ ( .A(_07262_ ), .B1(_07260_ ), .B2(_07269_ ), .ZN(_07689_ ) );
AND3_X1 _15718_ ( .A1(_07316_ ), .A2(_07319_ ), .A3(_07433_ ), .ZN(_07690_ ) );
NOR3_X1 _15719_ ( .A1(_07689_ ), .A2(_07690_ ), .A3(_07630_ ), .ZN(_07691_ ) );
AOI21_X1 _15720_ ( .A(_07262_ ), .B1(_07307_ ), .B2(_07311_ ), .ZN(_07692_ ) );
AOI21_X1 _15721_ ( .A(_07301_ ), .B1(_07297_ ), .B2(_07300_ ), .ZN(_07693_ ) );
OR2_X1 _15722_ ( .A1(_07692_ ), .A2(_07693_ ), .ZN(_07694_ ) );
AOI211_X1 _15723_ ( .A(_07688_ ), .B(_07691_ ), .C1(_07638_ ), .C2(_07694_ ), .ZN(_07695_ ) );
BUF_X2 _15724_ ( .A(_07578_ ), .Z(_07696_ ) );
BUF_X2 _15725_ ( .A(_07262_ ), .Z(_07697_ ) );
AND4_X1 _15726_ ( .A1(_07688_ ), .A2(_07696_ ), .A3(_07697_ ), .A4(_07277_ ), .ZN(_07698_ ) );
OAI21_X1 _15727_ ( .A(_07254_ ), .B1(_07695_ ), .B2(_07698_ ), .ZN(_07699_ ) );
NAND2_X1 _15728_ ( .A1(_04568_ ), .A2(_07327_ ), .ZN(_07700_ ) );
AND2_X1 _15729_ ( .A1(_04567_ ), .A2(_03695_ ), .ZN(_07701_ ) );
OR2_X1 _15730_ ( .A1(_07701_ ), .A2(_07524_ ), .ZN(_07702_ ) );
AND4_X1 _15731_ ( .A1(_07687_ ), .A2(_07699_ ), .A3(_07700_ ), .A4(_07702_ ), .ZN(_07703_ ) );
OAI21_X1 _15732_ ( .A(_04575_ ), .B1(_07353_ ), .B2(_07382_ ), .ZN(_07704_ ) );
INV_X1 _15733_ ( .A(_04573_ ), .ZN(_07705_ ) );
AND3_X1 _15734_ ( .A1(_07704_ ), .A2(_04568_ ), .A3(_07705_ ), .ZN(_07706_ ) );
AOI21_X1 _15735_ ( .A(_04568_ ), .B1(_07704_ ), .B2(_07705_ ), .ZN(_07707_ ) );
OAI21_X1 _15736_ ( .A(_07404_ ), .B1(_07706_ ), .B2(_07707_ ), .ZN(_07708_ ) );
AOI22_X1 _15737_ ( .A1(_07686_ ), .A2(_07408_ ), .B1(_07388_ ), .B2(_07409_ ), .ZN(_07709_ ) );
NAND3_X1 _15738_ ( .A1(_07703_ ), .A2(_07708_ ), .A3(_07709_ ), .ZN(_07710_ ) );
AOI21_X1 _15739_ ( .A(_07672_ ), .B1(_07710_ ), .B2(_07421_ ), .ZN(_07711_ ) );
NAND2_X1 _15740_ ( .A1(_04976_ ), .A2(_07663_ ), .ZN(_07712_ ) );
NAND2_X1 _15741_ ( .A1(_07712_ ), .A2(_07665_ ), .ZN(_07713_ ) );
OAI21_X1 _15742_ ( .A(_07667_ ), .B1(_07711_ ), .B2(_07713_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _15743_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_06605_ ), .ZN(_07714_ ) );
NAND3_X1 _15744_ ( .A1(_06787_ ), .A2(\mtvec [16] ), .A3(_04987_ ), .ZN(_07715_ ) );
NAND3_X1 _15745_ ( .A1(_06787_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_04991_ ), .ZN(_07716_ ) );
NAND4_X1 _15746_ ( .A1(_05456_ ), .A2(_04896_ ), .A3(\mepc [16] ), .A4(_04992_ ), .ZN(_07717_ ) );
NAND4_X1 _15747_ ( .A1(_07715_ ), .A2(_07716_ ), .A3(_05017_ ), .A4(_07717_ ), .ZN(_07718_ ) );
OAI211_X1 _15748_ ( .A(_07424_ ), .B(_07714_ ), .C1(_07083_ ), .C2(_07718_ ), .ZN(_07719_ ) );
AOI21_X1 _15749_ ( .A(_07600_ ), .B1(_04457_ ), .B2(_03747_ ), .ZN(_07720_ ) );
OAI21_X1 _15750_ ( .A(_07720_ ), .B1(_03747_ ), .B2(_04457_ ), .ZN(_07721_ ) );
AOI22_X1 _15751_ ( .A1(_05011_ ), .A2(_07603_ ), .B1(\ID_EX_imm [16] ), .B2(_07539_ ), .ZN(_07722_ ) );
AOI21_X1 _15752_ ( .A(_07531_ ), .B1(_07721_ ), .B2(_07722_ ), .ZN(_07723_ ) );
OR2_X1 _15753_ ( .A1(_07723_ ), .A2(_07662_ ), .ZN(_07724_ ) );
BUF_X2 _15754_ ( .A(_07137_ ), .Z(_07725_ ) );
OAI211_X1 _15755_ ( .A(_07200_ ), .B(_07725_ ), .C1(_07688_ ), .C2(_07135_ ), .ZN(_07726_ ) );
INV_X1 _15756_ ( .A(_07726_ ), .ZN(_07727_ ) );
OR3_X1 _15757_ ( .A1(_07439_ ), .A2(_07442_ ), .A3(_04640_ ), .ZN(_07728_ ) );
OR3_X1 _15758_ ( .A1(_07264_ ), .A2(_07494_ ), .A3(_07488_ ), .ZN(_07729_ ) );
OR3_X1 _15759_ ( .A1(_07497_ ), .A2(_07495_ ), .A3(_07201_ ), .ZN(_07730_ ) );
NAND3_X1 _15760_ ( .A1(_07729_ ), .A2(_07730_ ), .A3(_07271_ ), .ZN(_07731_ ) );
AOI21_X1 _15761_ ( .A(_07209_ ), .B1(_07728_ ), .B2(_07731_ ), .ZN(_07732_ ) );
OR3_X1 _15762_ ( .A1(_07447_ ), .A2(_07450_ ), .A3(_04641_ ), .ZN(_07733_ ) );
OAI21_X1 _15763_ ( .A(_07733_ ), .B1(_07458_ ), .B2(_07261_ ), .ZN(_07734_ ) );
AOI21_X1 _15764_ ( .A(_07732_ ), .B1(_07734_ ), .B2(_07322_ ), .ZN(_07735_ ) );
AND2_X1 _15765_ ( .A1(_07735_ ), .A2(_07464_ ), .ZN(_07736_ ) );
OAI21_X1 _15766_ ( .A(_07131_ ), .B1(_07727_ ), .B2(_07736_ ), .ZN(_07737_ ) );
OR3_X1 _15767_ ( .A1(_07469_ ), .A2(_07473_ ), .A3(_07301_ ), .ZN(_07738_ ) );
NAND2_X1 _15768_ ( .A1(_07512_ ), .A2(_07650_ ), .ZN(_07739_ ) );
AOI21_X1 _15769_ ( .A(_07696_ ), .B1(_07738_ ), .B2(_07739_ ), .ZN(_07740_ ) );
AOI21_X1 _15770_ ( .A(_07301_ ), .B1(_07489_ ), .B2(_07492_ ), .ZN(_07741_ ) );
AOI21_X1 _15771_ ( .A(_07262_ ), .B1(_07481_ ), .B2(_07484_ ), .ZN(_07742_ ) );
NOR3_X1 _15772_ ( .A1(_07741_ ), .A2(_07742_ ), .A3(_07280_ ), .ZN(_07743_ ) );
OAI21_X1 _15773_ ( .A(_07464_ ), .B1(_07740_ ), .B2(_07743_ ), .ZN(_07744_ ) );
AND3_X1 _15774_ ( .A1(_07503_ ), .A2(_07262_ ), .A3(_07304_ ), .ZN(_07745_ ) );
NAND2_X1 _15775_ ( .A1(_07638_ ), .A2(_07745_ ), .ZN(_07746_ ) );
AOI21_X1 _15776_ ( .A(_07255_ ), .B1(_07746_ ), .B2(_07284_ ), .ZN(_07747_ ) );
NAND2_X1 _15777_ ( .A1(_07744_ ), .A2(_07747_ ), .ZN(_07748_ ) );
NAND3_X1 _15778_ ( .A1(_07735_ ), .A2(_07560_ ), .A3(_07408_ ), .ZN(_07749_ ) );
NAND3_X1 _15779_ ( .A1(_07737_ ), .A2(_07748_ ), .A3(_07749_ ), .ZN(_07750_ ) );
OAI21_X1 _15780_ ( .A(_07403_ ), .B1(_07384_ ), .B2(_04575_ ), .ZN(_07751_ ) );
AOI21_X1 _15781_ ( .A(_07751_ ), .B1(_04575_ ), .B2(_07384_ ), .ZN(_07752_ ) );
BUF_X4 _15782_ ( .A(_04768_ ), .Z(_07753_ ) );
NOR3_X1 _15783_ ( .A1(_04573_ ), .A2(_04574_ ), .A3(_07753_ ), .ZN(_07754_ ) );
NOR3_X1 _15784_ ( .A1(_04571_ ), .A2(_04572_ ), .A3(_07521_ ), .ZN(_07755_ ) );
AOI21_X1 _15785_ ( .A(_07524_ ), .B1(_04571_ ), .B2(_04572_ ), .ZN(_07756_ ) );
OR3_X1 _15786_ ( .A1(_07754_ ), .A2(_07755_ ), .A3(_07756_ ), .ZN(_07757_ ) );
OR3_X1 _15787_ ( .A1(_07750_ ), .A2(_07752_ ), .A3(_07757_ ), .ZN(_07758_ ) );
AOI21_X1 _15788_ ( .A(_07724_ ), .B1(_07758_ ), .B2(_07421_ ), .ZN(_07759_ ) );
NAND2_X1 _15789_ ( .A1(_05009_ ), .A2(_07663_ ), .ZN(_07760_ ) );
NAND2_X1 _15790_ ( .A1(_07760_ ), .A2(_07665_ ), .ZN(_07761_ ) );
OAI21_X1 _15791_ ( .A(_07719_ ), .B1(_07759_ ), .B2(_07761_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
NAND2_X1 _15792_ ( .A1(_06794_ ), .A2(_06706_ ), .ZN(_07762_ ) );
INV_X1 _15793_ ( .A(_04201_ ), .ZN(_07763_ ) );
INV_X1 _15794_ ( .A(_04223_ ), .ZN(_07764_ ) );
NAND2_X1 _15795_ ( .A1(_04454_ ), .A2(_04321_ ), .ZN(_07765_ ) );
AOI211_X1 _15796_ ( .A(_07763_ ), .B(_07764_ ), .C1(_07765_ ), .C2(_04434_ ), .ZN(_07766_ ) );
OAI21_X1 _15797_ ( .A(_04177_ ), .B1(_07766_ ), .B2(_04425_ ), .ZN(_07767_ ) );
INV_X1 _15798_ ( .A(_04155_ ), .ZN(_07768_ ) );
NAND2_X1 _15799_ ( .A1(_04176_ ), .A2(_03118_ ), .ZN(_07769_ ) );
AND3_X1 _15800_ ( .A1(_07767_ ), .A2(_07768_ ), .A3(_07769_ ), .ZN(_07770_ ) );
AOI21_X1 _15801_ ( .A(_07768_ ), .B1(_07767_ ), .B2(_07769_ ), .ZN(_07771_ ) );
OR3_X1 _15802_ ( .A1(_07770_ ), .A2(_07771_ ), .A3(_07599_ ), .ZN(_07772_ ) );
AOI22_X1 _15803_ ( .A1(_05044_ ), .A2(_07603_ ), .B1(\ID_EX_imm [15] ), .B2(_07539_ ), .ZN(_07773_ ) );
AOI21_X1 _15804_ ( .A(_07531_ ), .B1(_07772_ ), .B2(_07773_ ), .ZN(_07774_ ) );
OR2_X1 _15805_ ( .A1(_07774_ ), .A2(_07662_ ), .ZN(_07775_ ) );
NAND3_X1 _15806_ ( .A1(_04691_ ), .A2(_03094_ ), .A3(_04419_ ), .ZN(_07776_ ) );
OAI21_X1 _15807_ ( .A(_07776_ ), .B1(_04592_ ), .B2(_07657_ ), .ZN(_07777_ ) );
NAND3_X1 _15808_ ( .A1(_07554_ ), .A2(_04641_ ), .A3(_07555_ ), .ZN(_07778_ ) );
NAND3_X1 _15809_ ( .A1(_07550_ ), .A2(_07271_ ), .A3(_07551_ ), .ZN(_07779_ ) );
NAND2_X1 _15810_ ( .A1(_07778_ ), .A2(_07779_ ), .ZN(_07780_ ) );
NAND2_X1 _15811_ ( .A1(_07780_ ), .A2(_07279_ ), .ZN(_07781_ ) );
NOR3_X1 _15812_ ( .A1(_07265_ ), .A2(_07298_ ), .A3(_07296_ ), .ZN(_07782_ ) );
NOR3_X1 _15813_ ( .A1(_07290_ ), .A2(_07299_ ), .A3(_07202_ ), .ZN(_07783_ ) );
OAI21_X1 _15814_ ( .A(_07261_ ), .B1(_07782_ ), .B2(_07783_ ), .ZN(_07784_ ) );
NAND3_X1 _15815_ ( .A1(_07547_ ), .A2(_07548_ ), .A3(_07206_ ), .ZN(_07785_ ) );
AND2_X1 _15816_ ( .A1(_07784_ ), .A2(_07785_ ), .ZN(_07786_ ) );
OAI211_X1 _15817_ ( .A(_07781_ ), .B(_07461_ ), .C1(_07323_ ), .C2(_07786_ ), .ZN(_07787_ ) );
AND3_X1 _15818_ ( .A1(_07240_ ), .A2(_04640_ ), .A3(_07202_ ), .ZN(_07788_ ) );
NAND2_X1 _15819_ ( .A1(_07788_ ), .A2(_07476_ ), .ZN(_07789_ ) );
NAND2_X1 _15820_ ( .A1(_07789_ ), .A2(_07688_ ), .ZN(_07790_ ) );
NAND3_X1 _15821_ ( .A1(_07787_ ), .A2(_07407_ ), .A3(_07790_ ), .ZN(_07791_ ) );
AND2_X1 _15822_ ( .A1(_07587_ ), .A2(_07588_ ), .ZN(_07792_ ) );
MUX2_X1 _15823_ ( .A(_07572_ ), .B(_07792_ ), .S(_07444_ ), .Z(_07793_ ) );
NAND2_X1 _15824_ ( .A1(_07793_ ), .A2(_07279_ ), .ZN(_07794_ ) );
OAI21_X1 _15825_ ( .A(_07272_ ), .B1(_07582_ ), .B2(_07583_ ), .ZN(_07795_ ) );
OAI21_X1 _15826_ ( .A(_07478_ ), .B1(_07574_ ), .B2(_07575_ ), .ZN(_07796_ ) );
NAND3_X1 _15827_ ( .A1(_07795_ ), .A2(_07477_ ), .A3(_07796_ ), .ZN(_07797_ ) );
AND2_X1 _15828_ ( .A1(_07249_ ), .A2(_04765_ ), .ZN(_07798_ ) );
BUF_X2 _15829_ ( .A(_07798_ ), .Z(_07799_ ) );
NAND3_X1 _15830_ ( .A1(_07794_ ), .A2(_07797_ ), .A3(_07799_ ), .ZN(_07800_ ) );
AND2_X1 _15831_ ( .A1(_07186_ ), .A2(_07725_ ), .ZN(_07801_ ) );
INV_X1 _15832_ ( .A(_07187_ ), .ZN(_07802_ ) );
AOI22_X1 _15833_ ( .A1(_07801_ ), .A2(_07802_ ), .B1(_07787_ ), .B2(_07790_ ), .ZN(_07803_ ) );
INV_X1 _15834_ ( .A(_07130_ ), .ZN(_07804_ ) );
BUF_X4 _15835_ ( .A(_07804_ ), .Z(_07805_ ) );
OAI211_X1 _15836_ ( .A(_07791_ ), .B(_07800_ ), .C1(_07803_ ), .C2(_07805_ ), .ZN(_07806_ ) );
AOI211_X1 _15837_ ( .A(_07777_ ), .B(_07806_ ), .C1(_04593_ ), .C2(_07327_ ), .ZN(_07807_ ) );
INV_X1 _15838_ ( .A(_07403_ ), .ZN(_07808_ ) );
BUF_X2 _15839_ ( .A(_07808_ ), .Z(_07809_ ) );
OAI21_X1 _15840_ ( .A(_07380_ ), .B1(_07369_ ), .B2(_07377_ ), .ZN(_07810_ ) );
AND2_X1 _15841_ ( .A1(_07810_ ), .A2(_07338_ ), .ZN(_07811_ ) );
INV_X1 _15842_ ( .A(_07811_ ), .ZN(_07812_ ) );
NAND2_X1 _15843_ ( .A1(_07812_ ), .A2(_07339_ ), .ZN(_07813_ ) );
AOI21_X1 _15844_ ( .A(_07349_ ), .B1(_07813_ ), .B2(_07348_ ), .ZN(_07814_ ) );
NOR2_X1 _15845_ ( .A1(_04596_ ), .A2(_04685_ ), .ZN(_07815_ ) );
OR2_X1 _15846_ ( .A1(_07814_ ), .A2(_07815_ ), .ZN(_07816_ ) );
XNOR2_X1 _15847_ ( .A(_07816_ ), .B(_04593_ ), .ZN(_07817_ ) );
OAI21_X1 _15848_ ( .A(_07807_ ), .B1(_07809_ ), .B2(_07817_ ), .ZN(_07818_ ) );
AOI21_X1 _15849_ ( .A(_07775_ ), .B1(_07818_ ), .B2(_07421_ ), .ZN(_07819_ ) );
OAI21_X1 _15850_ ( .A(_06994_ ), .B1(_05038_ ), .B2(_05663_ ), .ZN(_07820_ ) );
OAI21_X1 _15851_ ( .A(_07762_ ), .B1(_07819_ ), .B2(_07820_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
OAI21_X1 _15852_ ( .A(_07424_ ), .B1(_05082_ ), .B2(_05083_ ), .ZN(_07821_ ) );
OR3_X1 _15853_ ( .A1(_07766_ ), .A2(_04177_ ), .A3(_04425_ ), .ZN(_07822_ ) );
NAND3_X1 _15854_ ( .A1(_07822_ ), .A2(_07126_ ), .A3(_07767_ ), .ZN(_07823_ ) );
AOI22_X1 _15855_ ( .A1(_05074_ ), .A2(_07603_ ), .B1(\ID_EX_imm [14] ), .B2(_07539_ ), .ZN(_07824_ ) );
AOI21_X1 _15856_ ( .A(_07531_ ), .B1(_07823_ ), .B2(_07824_ ), .ZN(_07825_ ) );
OR2_X1 _15857_ ( .A1(_07825_ ), .A2(_07662_ ), .ZN(_07826_ ) );
AND2_X2 _15858_ ( .A1(_07137_ ), .A2(_07802_ ), .ZN(_07827_ ) );
NAND3_X1 _15859_ ( .A1(_07273_ ), .A2(_07242_ ), .A3(_07304_ ), .ZN(_07828_ ) );
OAI211_X1 _15860_ ( .A(_07200_ ), .B(_07827_ ), .C1(_07544_ ), .C2(_07828_ ), .ZN(_07829_ ) );
OAI21_X1 _15861_ ( .A(_07265_ ), .B1(_07494_ ), .B2(_07488_ ), .ZN(_07830_ ) );
OAI21_X1 _15862_ ( .A(_07472_ ), .B1(_07487_ ), .B2(_07491_ ), .ZN(_07831_ ) );
NAND3_X1 _15863_ ( .A1(_07830_ ), .A2(_07831_ ), .A3(_07272_ ), .ZN(_07832_ ) );
NAND2_X1 _15864_ ( .A1(_07617_ ), .A2(_07618_ ), .ZN(_07833_ ) );
OAI211_X1 _15865_ ( .A(_07832_ ), .B(_07476_ ), .C1(_07833_ ), .C2(_07433_ ), .ZN(_07834_ ) );
OAI21_X1 _15866_ ( .A(_07206_ ), .B1(_07622_ ), .B2(_07623_ ), .ZN(_07835_ ) );
NAND3_X1 _15867_ ( .A1(_07614_ ), .A2(_07272_ ), .A3(_07615_ ), .ZN(_07836_ ) );
NAND2_X1 _15868_ ( .A1(_07835_ ), .A2(_07836_ ), .ZN(_07837_ ) );
OAI211_X1 _15869_ ( .A(_07834_ ), .B(_07249_ ), .C1(_07837_ ), .C2(_07578_ ), .ZN(_07838_ ) );
NAND4_X1 _15870_ ( .A1(_07625_ ), .A2(_07283_ ), .A3(_07578_ ), .A4(_07273_ ), .ZN(_07839_ ) );
AND2_X1 _15871_ ( .A1(_07838_ ), .A2(_07839_ ), .ZN(_07840_ ) );
AOI21_X1 _15872_ ( .A(_07805_ ), .B1(_07829_ ), .B2(_07840_ ), .ZN(_07841_ ) );
AND3_X1 _15873_ ( .A1(_07813_ ), .A2(_07349_ ), .A3(_07348_ ), .ZN(_07842_ ) );
NOR3_X1 _15874_ ( .A1(_07842_ ), .A2(_07814_ ), .A3(_07809_ ), .ZN(_07843_ ) );
NOR2_X1 _15875_ ( .A1(_07631_ ), .A2(_07632_ ), .ZN(_07844_ ) );
MUX2_X1 _15876_ ( .A(_07649_ ), .B(_07844_ ), .S(_04640_ ), .Z(_07845_ ) );
NAND2_X1 _15877_ ( .A1(_07845_ ), .A2(_07209_ ), .ZN(_07846_ ) );
OAI21_X1 _15878_ ( .A(_07444_ ), .B1(_07634_ ), .B2(_07635_ ), .ZN(_07847_ ) );
OAI21_X1 _15879_ ( .A(_07271_ ), .B1(_07639_ ), .B2(_07641_ ), .ZN(_07848_ ) );
NAND3_X1 _15880_ ( .A1(_07847_ ), .A2(_07848_ ), .A3(_07476_ ), .ZN(_07849_ ) );
AND3_X1 _15881_ ( .A1(_07846_ ), .A2(_07799_ ), .A3(_07849_ ), .ZN(_07850_ ) );
AOI221_X4 _15882_ ( .A(_07850_ ), .B1(_07815_ ), .B2(_04419_ ), .C1(_04597_ ), .C2(_07326_ ), .ZN(_07851_ ) );
INV_X1 _15883_ ( .A(_07406_ ), .ZN(_07852_ ) );
OR2_X1 _15884_ ( .A1(_07840_ ), .A2(_07852_ ), .ZN(_07853_ ) );
OAI21_X1 _15885_ ( .A(_07329_ ), .B1(_04686_ ), .B2(_03118_ ), .ZN(_07854_ ) );
NAND3_X1 _15886_ ( .A1(_07851_ ), .A2(_07853_ ), .A3(_07854_ ), .ZN(_07855_ ) );
OR3_X1 _15887_ ( .A1(_07841_ ), .A2(_07843_ ), .A3(_07855_ ), .ZN(_07856_ ) );
AOI21_X1 _15888_ ( .A(_07826_ ), .B1(_07856_ ), .B2(_07421_ ), .ZN(_07857_ ) );
NAND2_X1 _15889_ ( .A1(_05071_ ), .A2(_07663_ ), .ZN(_07858_ ) );
NAND2_X1 _15890_ ( .A1(_07858_ ), .A2(_07665_ ), .ZN(_07859_ ) );
OAI21_X1 _15891_ ( .A(_07821_ ), .B1(_07857_ ), .B2(_07859_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
OAI211_X1 _15892_ ( .A(_07424_ ), .B(_06820_ ), .C1(_06822_ ), .C2(_05108_ ), .ZN(_07860_ ) );
AND2_X1 _15893_ ( .A1(_07765_ ), .A2(_04434_ ), .ZN(_07861_ ) );
OR2_X1 _15894_ ( .A1(_07861_ ), .A2(_07764_ ), .ZN(_07862_ ) );
INV_X1 _15895_ ( .A(_04423_ ), .ZN(_07863_ ) );
AND3_X1 _15896_ ( .A1(_07862_ ), .A2(_07763_ ), .A3(_07863_ ), .ZN(_07864_ ) );
AOI21_X1 _15897_ ( .A(_07763_ ), .B1(_07862_ ), .B2(_07863_ ), .ZN(_07865_ ) );
NOR3_X1 _15898_ ( .A1(_07864_ ), .A2(_07865_ ), .A3(_07600_ ), .ZN(_07866_ ) );
AND2_X1 _15899_ ( .A1(_05101_ ), .A2(_07428_ ), .ZN(_07867_ ) );
AND3_X1 _15900_ ( .A1(_07112_ ), .A2(\ID_EX_imm [13] ), .A3(_07109_ ), .ZN(_07868_ ) );
NOR3_X1 _15901_ ( .A1(_07866_ ), .A2(_07867_ ), .A3(_07868_ ), .ZN(_07869_ ) );
AOI21_X1 _15902_ ( .A(_05495_ ), .B1(_07869_ ), .B2(_05672_ ), .ZN(_07870_ ) );
OR2_X1 _15903_ ( .A1(_07170_ ), .A2(_07185_ ), .ZN(_07871_ ) );
AND2_X1 _15904_ ( .A1(_07210_ ), .A2(_07207_ ), .ZN(_07872_ ) );
NOR4_X1 _15905_ ( .A1(_07871_ ), .A2(_07187_ ), .A3(_07138_ ), .A4(_07872_ ), .ZN(_07873_ ) );
NOR3_X1 _15906_ ( .A1(_07246_ ), .A2(_07322_ ), .A3(_07478_ ), .ZN(_07874_ ) );
OR2_X1 _15907_ ( .A1(_07874_ ), .A2(_07250_ ), .ZN(_07875_ ) );
AND2_X1 _15908_ ( .A1(_07677_ ), .A2(_07678_ ), .ZN(_07876_ ) );
OAI21_X1 _15909_ ( .A(_07229_ ), .B1(_07305_ ), .B2(_07295_ ), .ZN(_07877_ ) );
OAI21_X1 _15910_ ( .A(_07220_ ), .B1(_07298_ ), .B2(_07296_ ), .ZN(_07878_ ) );
NAND2_X1 _15911_ ( .A1(_07877_ ), .A2(_07878_ ), .ZN(_07879_ ) );
INV_X1 _15912_ ( .A(_07879_ ), .ZN(_07880_ ) );
MUX2_X1 _15913_ ( .A(_07876_ ), .B(_07880_ ), .S(_07271_ ), .Z(_07881_ ) );
NAND2_X1 _15914_ ( .A1(_07881_ ), .A2(_07630_ ), .ZN(_07882_ ) );
NAND2_X1 _15915_ ( .A1(_07239_ ), .A2(_07514_ ), .ZN(_07883_ ) );
NAND3_X1 _15916_ ( .A1(_07882_ ), .A2(_07461_ ), .A3(_07883_ ), .ZN(_07884_ ) );
AND2_X1 _15917_ ( .A1(_07875_ ), .A2(_07884_ ), .ZN(_07885_ ) );
OAI21_X1 _15918_ ( .A(_07131_ ), .B1(_07873_ ), .B2(_07885_ ), .ZN(_07886_ ) );
NAND3_X1 _15919_ ( .A1(_07875_ ), .A2(_07408_ ), .A3(_07884_ ), .ZN(_07887_ ) );
NOR2_X1 _15920_ ( .A1(_07278_ ), .A2(_07696_ ), .ZN(_07888_ ) );
NOR3_X1 _15921_ ( .A1(_07312_ ), .A2(_07320_ ), .A3(_07280_ ), .ZN(_07889_ ) );
OAI21_X1 _15922_ ( .A(_07799_ ), .B1(_07888_ ), .B2(_07889_ ), .ZN(_07890_ ) );
AOI22_X1 _15923_ ( .A1(_04607_ ), .A2(_07327_ ), .B1(_07344_ ), .B2(_07409_ ), .ZN(_07891_ ) );
AND4_X1 _15924_ ( .A1(_07886_ ), .A2(_07887_ ), .A3(_07890_ ), .A4(_07891_ ), .ZN(_07892_ ) );
OR2_X1 _15925_ ( .A1(_07811_ ), .A2(_04603_ ), .ZN(_07893_ ) );
INV_X1 _15926_ ( .A(_07347_ ), .ZN(_07894_ ) );
AOI21_X1 _15927_ ( .A(_04607_ ), .B1(_07893_ ), .B2(_07894_ ), .ZN(_07895_ ) );
AOI211_X1 _15928_ ( .A(_07347_ ), .B(_04608_ ), .C1(_07812_ ), .C2(_04602_ ), .ZN(_07896_ ) );
OAI21_X1 _15929_ ( .A(_07404_ ), .B1(_07895_ ), .B2(_07896_ ), .ZN(_07897_ ) );
OR2_X1 _15930_ ( .A1(_07345_ ), .A2(_07657_ ), .ZN(_07898_ ) );
NAND3_X1 _15931_ ( .A1(_07892_ ), .A2(_07897_ ), .A3(_07898_ ), .ZN(_07899_ ) );
AOI21_X1 _15932_ ( .A(_07870_ ), .B1(_07899_ ), .B2(_07421_ ), .ZN(_07900_ ) );
NAND2_X1 _15933_ ( .A1(_05097_ ), .A2(_07663_ ), .ZN(_07901_ ) );
NAND2_X1 _15934_ ( .A1(_07901_ ), .A2(_07665_ ), .ZN(_07902_ ) );
OAI21_X1 _15935_ ( .A(_07860_ ), .B1(_07900_ ), .B2(_07902_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
OR3_X1 _15936_ ( .A1(_05284_ ), .A2(_05285_ ), .A3(\EX_LS_result_csreg_mem [12] ), .ZN(_07903_ ) );
NAND3_X1 _15937_ ( .A1(_06787_ ), .A2(\mtvec [12] ), .A3(_04987_ ), .ZN(_07904_ ) );
NAND3_X1 _15938_ ( .A1(_06787_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_04991_ ), .ZN(_07905_ ) );
NAND4_X1 _15939_ ( .A1(_05456_ ), .A2(_04896_ ), .A3(\mepc [12] ), .A4(_04992_ ), .ZN(_07906_ ) );
NAND4_X1 _15940_ ( .A1(_07904_ ), .A2(_07905_ ), .A3(_06834_ ), .A4(_07906_ ), .ZN(_07907_ ) );
OAI211_X1 _15941_ ( .A(_06802_ ), .B(_07903_ ), .C1(_07083_ ), .C2(_07907_ ), .ZN(_07908_ ) );
NAND3_X1 _15942_ ( .A1(_07765_ ), .A2(_07764_ ), .A3(_04434_ ), .ZN(_07909_ ) );
NAND3_X1 _15943_ ( .A1(_07862_ ), .A2(_07126_ ), .A3(_07909_ ), .ZN(_07910_ ) );
AOI22_X1 _15944_ ( .A1(_05135_ ), .A2(_07603_ ), .B1(\ID_EX_imm [12] ), .B2(_07539_ ), .ZN(_07911_ ) );
AOI21_X1 _15945_ ( .A(_07531_ ), .B1(_07910_ ), .B2(_07911_ ), .ZN(_07912_ ) );
OR2_X1 _15946_ ( .A1(_07912_ ), .A2(_07662_ ), .ZN(_07913_ ) );
BUF_X4 _15947_ ( .A(_07186_ ), .Z(_07914_ ) );
OAI211_X1 _15948_ ( .A(_07914_ ), .B(_07827_ ), .C1(_07434_ ), .C2(_07544_ ), .ZN(_07915_ ) );
BUF_X2 _15949_ ( .A(_07272_ ), .Z(_07916_ ) );
AND3_X1 _15950_ ( .A1(_07458_ ), .A2(_07578_ ), .A3(_07916_ ), .ZN(_07917_ ) );
OR2_X1 _15951_ ( .A1(_07917_ ), .A2(_07251_ ), .ZN(_07918_ ) );
NAND2_X1 _15952_ ( .A1(_07452_ ), .A2(_07280_ ), .ZN(_07919_ ) );
BUF_X4 _15953_ ( .A(_07323_ ), .Z(_07920_ ) );
NAND3_X1 _15954_ ( .A1(_07729_ ), .A2(_07730_ ), .A3(_07650_ ), .ZN(_07921_ ) );
OR3_X1 _15955_ ( .A1(_07487_ ), .A2(_07491_ ), .A3(_07202_ ), .ZN(_07922_ ) );
OAI211_X1 _15956_ ( .A(_07483_ ), .B(_07258_ ), .C1(_04179_ ), .C2(_07204_ ), .ZN(_07923_ ) );
NAND3_X1 _15957_ ( .A1(_07922_ ), .A2(_07273_ ), .A3(_07923_ ), .ZN(_07924_ ) );
NAND2_X1 _15958_ ( .A1(_07921_ ), .A2(_07924_ ), .ZN(_07925_ ) );
OAI211_X1 _15959_ ( .A(_07919_ ), .B(_07464_ ), .C1(_07920_ ), .C2(_07925_ ), .ZN(_07926_ ) );
NAND2_X1 _15960_ ( .A1(_07918_ ), .A2(_07926_ ), .ZN(_07927_ ) );
AOI21_X1 _15961_ ( .A(_07805_ ), .B1(_07915_ ), .B2(_07927_ ), .ZN(_07928_ ) );
AND3_X1 _15962_ ( .A1(_07918_ ), .A2(_07408_ ), .A3(_07926_ ), .ZN(_07929_ ) );
INV_X1 _15963_ ( .A(_07798_ ), .ZN(_07930_ ) );
OR2_X1 _15964_ ( .A1(_07513_ ), .A2(_07638_ ), .ZN(_07931_ ) );
OAI21_X1 _15965_ ( .A(_07638_ ), .B1(_07475_ ), .B2(_07485_ ), .ZN(_07932_ ) );
AOI21_X1 _15966_ ( .A(_07930_ ), .B1(_07931_ ), .B2(_07932_ ), .ZN(_07933_ ) );
NOR3_X1 _15967_ ( .A1(_07928_ ), .A2(_07929_ ), .A3(_07933_ ), .ZN(_07934_ ) );
AOI21_X1 _15968_ ( .A(_07809_ ), .B1(_07812_ ), .B2(_04602_ ), .ZN(_07935_ ) );
OAI21_X1 _15969_ ( .A(_07935_ ), .B1(_04602_ ), .B2(_07812_ ), .ZN(_07936_ ) );
AND2_X1 _15970_ ( .A1(_04602_ ), .A2(_07327_ ), .ZN(_07937_ ) );
NOR3_X1 _15971_ ( .A1(_04601_ ), .A2(_06840_ ), .A3(_07521_ ), .ZN(_07938_ ) );
AOI21_X1 _15972_ ( .A(_07657_ ), .B1(_04601_ ), .B2(_06840_ ), .ZN(_07939_ ) );
NOR3_X1 _15973_ ( .A1(_07937_ ), .A2(_07938_ ), .A3(_07939_ ), .ZN(_07940_ ) );
NAND3_X1 _15974_ ( .A1(_07934_ ), .A2(_07936_ ), .A3(_07940_ ), .ZN(_07941_ ) );
AOI21_X1 _15975_ ( .A(_07913_ ), .B1(_07941_ ), .B2(_07421_ ), .ZN(_07942_ ) );
OAI21_X1 _15976_ ( .A(_06994_ ), .B1(_05134_ ), .B2(_05663_ ), .ZN(_07943_ ) );
OAI21_X1 _15977_ ( .A(_07908_ ), .B1(_07942_ ), .B2(_07943_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
OR2_X1 _15978_ ( .A1(_03579_ ), .A2(_06700_ ), .ZN(_07944_ ) );
INV_X1 _15979_ ( .A(_04724_ ), .ZN(_07945_ ) );
AND2_X1 _15980_ ( .A1(_04550_ ), .A2(_04546_ ), .ZN(_07946_ ) );
AND3_X1 _15981_ ( .A1(_07946_ ), .A2(_04540_ ), .A3(_04536_ ), .ZN(_07947_ ) );
OAI21_X2 _15982_ ( .A(_07947_ ), .B1(_07386_ ), .B2(_07394_ ), .ZN(_07948_ ) );
AOI21_X1 _15983_ ( .A(_04698_ ), .B1(_04546_ ), .B2(_07398_ ), .ZN(_07949_ ) );
INV_X1 _15984_ ( .A(_04536_ ), .ZN(_07950_ ) );
OR3_X1 _15985_ ( .A1(_07949_ ), .A2(_04695_ ), .A3(_07950_ ), .ZN(_07951_ ) );
NAND2_X1 _15986_ ( .A1(_07149_ ), .A2(_02548_ ), .ZN(_07952_ ) );
INV_X1 _15987_ ( .A(_02522_ ), .ZN(_07953_ ) );
NOR2_X1 _15988_ ( .A1(_04535_ ), .A2(_07953_ ), .ZN(_07954_ ) );
NAND2_X1 _15989_ ( .A1(_04540_ ), .A2(_07954_ ), .ZN(_07955_ ) );
AND3_X1 _15990_ ( .A1(_07951_ ), .A2(_07952_ ), .A3(_07955_ ), .ZN(_07956_ ) );
AND2_X2 _15991_ ( .A1(_07948_ ), .A2(_07956_ ), .ZN(_07957_ ) );
INV_X2 _15992_ ( .A(_07957_ ), .ZN(_07958_ ) );
NAND3_X2 _15993_ ( .A1(_07958_ ), .A2(_04731_ ), .A3(_04738_ ), .ZN(_07959_ ) );
AOI21_X1 _15994_ ( .A(_04736_ ), .B1(_04738_ ), .B2(_04729_ ), .ZN(_07960_ ) );
AOI211_X2 _15995_ ( .A(_04745_ ), .B(_07945_ ), .C1(_07959_ ), .C2(_07960_ ), .ZN(_07961_ ) );
INV_X1 _15996_ ( .A(_07961_ ), .ZN(_07962_ ) );
NOR2_X1 _15997_ ( .A1(_04490_ ), .A2(_04716_ ), .ZN(_07963_ ) );
AOI21_X1 _15998_ ( .A(_07963_ ), .B1(_04717_ ), .B2(_04722_ ), .ZN(_07964_ ) );
AOI21_X2 _15999_ ( .A(_04531_ ), .B1(_07962_ ), .B2(_07964_ ), .ZN(_07965_ ) );
AND2_X1 _16000_ ( .A1(_04524_ ), .A2(_03276_ ), .ZN(_07966_ ) );
AND2_X1 _16001_ ( .A1(_03253_ ), .A2(_04529_ ), .ZN(_07967_ ) );
OR3_X4 _16002_ ( .A1(_07965_ ), .A2(_07966_ ), .A3(_07967_ ), .ZN(_07968_ ) );
NOR2_X1 _16003_ ( .A1(_04524_ ), .A2(_03276_ ), .ZN(_07969_ ) );
INV_X1 _16004_ ( .A(_07969_ ), .ZN(_07970_ ) );
AND3_X2 _16005_ ( .A1(_07968_ ), .A2(_07970_ ), .A3(_04515_ ), .ZN(_07971_ ) );
AOI21_X1 _16006_ ( .A(_04515_ ), .B1(_07968_ ), .B2(_07970_ ), .ZN(_07972_ ) );
OR3_X1 _16007_ ( .A1(_07971_ ), .A2(_07972_ ), .A3(_07809_ ), .ZN(_07973_ ) );
AOI21_X1 _16008_ ( .A(_07523_ ), .B1(_07154_ ), .B2(_03310_ ), .ZN(_07974_ ) );
AND3_X1 _16009_ ( .A1(_07457_ ), .A2(_07272_ ), .A3(_07292_ ), .ZN(_07975_ ) );
NAND2_X1 _16010_ ( .A1(_07975_ ), .A2(_07477_ ), .ZN(_07976_ ) );
NOR3_X1 _16011_ ( .A1(_07976_ ), .A2(_07283_ ), .A3(_07852_ ), .ZN(_07977_ ) );
AOI211_X1 _16012_ ( .A(_07974_ ), .B(_07977_ ), .C1(_04515_ ), .C2(_07326_ ), .ZN(_07978_ ) );
NOR2_X1 _16013_ ( .A1(_07249_ ), .A2(_07255_ ), .ZN(_07979_ ) );
NAND3_X1 _16014_ ( .A1(_07846_ ), .A2(_07849_ ), .A3(_07979_ ), .ZN(_07980_ ) );
NAND3_X1 _16015_ ( .A1(_07456_ ), .A2(_04514_ ), .A3(_04419_ ), .ZN(_07981_ ) );
NAND3_X1 _16016_ ( .A1(_07978_ ), .A2(_07980_ ), .A3(_07981_ ), .ZN(_07982_ ) );
AOI21_X1 _16017_ ( .A(_07802_ ), .B1(_07186_ ), .B2(_07211_ ), .ZN(_07983_ ) );
NOR2_X1 _16018_ ( .A1(_07608_ ), .A2(_07983_ ), .ZN(_07984_ ) );
INV_X1 _16019_ ( .A(_07984_ ), .ZN(_07985_ ) );
NAND3_X1 _16020_ ( .A1(_07914_ ), .A2(_07725_ ), .A3(_07828_ ), .ZN(_07986_ ) );
OR2_X1 _16021_ ( .A1(_07976_ ), .A2(_07283_ ), .ZN(_07987_ ) );
AND2_X1 _16022_ ( .A1(_07986_ ), .A2(_07987_ ), .ZN(_07988_ ) );
AOI21_X1 _16023_ ( .A(_07804_ ), .B1(_07985_ ), .B2(_07988_ ), .ZN(_07989_ ) );
OR3_X1 _16024_ ( .A1(_07437_ ), .A2(_07292_ ), .A3(_07446_ ), .ZN(_07990_ ) );
NOR2_X1 _16025_ ( .A1(_07445_ ), .A2(_07449_ ), .ZN(_07991_ ) );
NAND2_X1 _16026_ ( .A1(_07991_ ), .A2(_07304_ ), .ZN(_07992_ ) );
NAND2_X1 _16027_ ( .A1(_07990_ ), .A2(_07992_ ), .ZN(_07993_ ) );
AOI21_X1 _16028_ ( .A(_07454_ ), .B1(_03310_ ), .B2(_07204_ ), .ZN(_07994_ ) );
NOR2_X1 _16029_ ( .A1(_07453_ ), .A2(_07448_ ), .ZN(_07995_ ) );
MUX2_X1 _16030_ ( .A(_07994_ ), .B(_07995_ ), .S(_07286_ ), .Z(_07996_ ) );
MUX2_X1 _16031_ ( .A(_07993_ ), .B(_07996_ ), .S(_07916_ ), .Z(_07997_ ) );
NOR2_X1 _16032_ ( .A1(_07997_ ), .A2(_07920_ ), .ZN(_07998_ ) );
OR3_X1 _16033_ ( .A1(_07643_ ), .A2(_07644_ ), .A3(_07433_ ), .ZN(_07999_ ) );
OAI21_X1 _16034_ ( .A(_07292_ ), .B1(_07440_ ), .B2(_07438_ ), .ZN(_08000_ ) );
OAI21_X1 _16035_ ( .A(_07286_ ), .B1(_07497_ ), .B2(_07441_ ), .ZN(_08001_ ) );
NAND2_X1 _16036_ ( .A1(_08000_ ), .A2(_08001_ ), .ZN(_08002_ ) );
NAND2_X1 _16037_ ( .A1(_08002_ ), .A2(_07916_ ), .ZN(_08003_ ) );
NAND2_X1 _16038_ ( .A1(_07999_ ), .A2(_08003_ ), .ZN(_08004_ ) );
AOI21_X1 _16039_ ( .A(_07998_ ), .B1(_07920_ ), .B2(_08004_ ), .ZN(_08005_ ) );
AOI211_X1 _16040_ ( .A(_07982_ ), .B(_07989_ ), .C1(_07799_ ), .C2(_08005_ ), .ZN(_08006_ ) );
AOI21_X1 _16041_ ( .A(_07419_ ), .B1(_07973_ ), .B2(_08006_ ), .ZN(_08007_ ) );
AOI22_X1 _16042_ ( .A1(_03515_ ), .A2(_07428_ ), .B1(\ID_EX_imm [30] ), .B2(_07539_ ), .ZN(_08008_ ) );
OAI21_X1 _16043_ ( .A(_04033_ ), .B1(_04458_ ), .B2(_04481_ ), .ZN(_08009_ ) );
NAND2_X1 _16044_ ( .A1(_08009_ ), .A2(_04494_ ), .ZN(_08010_ ) );
AOI21_X1 _16045_ ( .A(_04499_ ), .B1(_08010_ ), .B2(_03893_ ), .ZN(_08011_ ) );
INV_X1 _16046_ ( .A(_03939_ ), .ZN(_08012_ ) );
AOI21_X1 _16047_ ( .A(_07600_ ), .B1(_08011_ ), .B2(_08012_ ), .ZN(_08013_ ) );
OAI21_X1 _16048_ ( .A(_08013_ ), .B1(_08012_ ), .B2(_08011_ ), .ZN(_08014_ ) );
AOI21_X1 _16049_ ( .A(_07531_ ), .B1(_08008_ ), .B2(_08014_ ), .ZN(_08015_ ) );
NOR3_X1 _16050_ ( .A1(_08007_ ), .A2(_07663_ ), .A3(_08015_ ), .ZN(_08016_ ) );
NAND2_X1 _16051_ ( .A1(_03600_ ), .A2(_07663_ ), .ZN(_08017_ ) );
NAND2_X1 _16052_ ( .A1(_08017_ ), .A2(_07665_ ), .ZN(_08018_ ) );
OAI21_X1 _16053_ ( .A(_07944_ ), .B1(_08016_ ), .B2(_08018_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _16054_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_06866_ ), .ZN(_08019_ ) );
OAI211_X1 _16055_ ( .A(_06802_ ), .B(_08019_ ), .C1(_07083_ ), .C2(_06864_ ), .ZN(_08020_ ) );
OR2_X1 _16056_ ( .A1(_05150_ ), .A2(_04782_ ), .ZN(_08021_ ) );
OAI211_X1 _16057_ ( .A(_07914_ ), .B(_07827_ ), .C1(_07543_ ), .C2(_07212_ ), .ZN(_08022_ ) );
NOR3_X1 _16058_ ( .A1(_07274_ ), .A2(_07306_ ), .A3(_07310_ ), .ZN(_08023_ ) );
NOR3_X1 _16059_ ( .A1(_07305_ ), .A2(_07295_ ), .A3(_07257_ ), .ZN(_08024_ ) );
OAI21_X1 _16060_ ( .A(_07261_ ), .B1(_08023_ ), .B2(_08024_ ), .ZN(_08025_ ) );
OAI21_X1 _16061_ ( .A(_07206_ ), .B1(_07782_ ), .B2(_07783_ ), .ZN(_08026_ ) );
NAND3_X1 _16062_ ( .A1(_08025_ ), .A2(_07477_ ), .A3(_08026_ ), .ZN(_08027_ ) );
OAI21_X1 _16063_ ( .A(_07322_ ), .B1(_07549_ ), .B2(_07552_ ), .ZN(_08028_ ) );
AND3_X1 _16064_ ( .A1(_08027_ ), .A2(_08028_ ), .A3(_07249_ ), .ZN(_08029_ ) );
AOI211_X1 _16065_ ( .A(_07249_ ), .B(_07279_ ), .C1(_07556_ ), .C2(_07557_ ), .ZN(_08030_ ) );
NOR2_X1 _16066_ ( .A1(_08029_ ), .A2(_08030_ ), .ZN(_08031_ ) );
AOI21_X1 _16067_ ( .A(_07804_ ), .B1(_08022_ ), .B2(_08031_ ), .ZN(_08032_ ) );
NOR2_X1 _16068_ ( .A1(_08031_ ), .A2(_07852_ ), .ZN(_08033_ ) );
OR2_X1 _16069_ ( .A1(_08032_ ), .A2(_08033_ ), .ZN(_08034_ ) );
NAND3_X1 _16070_ ( .A1(_07573_ ), .A2(_07576_ ), .A3(_07630_ ), .ZN(_08035_ ) );
NAND2_X1 _16071_ ( .A1(_07589_ ), .A2(_07323_ ), .ZN(_08036_ ) );
AOI21_X1 _16072_ ( .A(_07930_ ), .B1(_08035_ ), .B2(_08036_ ), .ZN(_08037_ ) );
NOR3_X1 _16073_ ( .A1(_04612_ ), .A2(_04249_ ), .A3(_07521_ ), .ZN(_08038_ ) );
OAI22_X1 _16074_ ( .A1(_04616_ ), .A2(_07753_ ), .B1(_04614_ ), .B2(_07524_ ), .ZN(_08039_ ) );
NOR4_X1 _16075_ ( .A1(_08034_ ), .A2(_08037_ ), .A3(_08038_ ), .A4(_08039_ ), .ZN(_08040_ ) );
OAI21_X1 _16076_ ( .A(_07379_ ), .B1(_07369_ ), .B2(_07377_ ), .ZN(_08041_ ) );
AOI21_X1 _16077_ ( .A(_04621_ ), .B1(_08041_ ), .B2(_07335_ ), .ZN(_08042_ ) );
NOR2_X1 _16078_ ( .A1(_04619_ ), .A2(_07308_ ), .ZN(_08043_ ) );
OR3_X1 _16079_ ( .A1(_08042_ ), .A2(_04615_ ), .A3(_08043_ ), .ZN(_08044_ ) );
OAI21_X1 _16080_ ( .A(_04615_ ), .B1(_08042_ ), .B2(_08043_ ), .ZN(_08045_ ) );
NAND3_X1 _16081_ ( .A1(_08044_ ), .A2(_07404_ ), .A3(_08045_ ), .ZN(_08046_ ) );
AOI21_X1 _16082_ ( .A(_07419_ ), .B1(_08040_ ), .B2(_08046_ ), .ZN(_08047_ ) );
OAI22_X1 _16083_ ( .A1(_05156_ ), .A2(_07111_ ), .B1(_02968_ ), .B2(_07115_ ), .ZN(_08048_ ) );
AND3_X1 _16084_ ( .A1(_04454_ ), .A2(_04298_ ), .A3(_04320_ ), .ZN(_08049_ ) );
OAI21_X1 _16085_ ( .A(_04272_ ), .B1(_08049_ ), .B2(_04430_ ), .ZN(_08050_ ) );
NAND2_X1 _16086_ ( .A1(_04271_ ), .A2(_03012_ ), .ZN(_08051_ ) );
AND2_X1 _16087_ ( .A1(_08050_ ), .A2(_08051_ ), .ZN(_08052_ ) );
XNOR2_X1 _16088_ ( .A(_08052_ ), .B(_04250_ ), .ZN(_08053_ ) );
AOI21_X1 _16089_ ( .A(_08048_ ), .B1(_08053_ ), .B2(_07126_ ), .ZN(_08054_ ) );
AOI21_X1 _16090_ ( .A(_05495_ ), .B1(_08054_ ), .B2(_05672_ ), .ZN(_08055_ ) );
OAI21_X1 _16091_ ( .A(_08021_ ), .B1(_08047_ ), .B2(_08055_ ), .ZN(_08056_ ) );
OAI21_X1 _16092_ ( .A(_08020_ ), .B1(_08056_ ), .B2(_06698_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OR3_X1 _16093_ ( .A1(_08049_ ), .A2(_04272_ ), .A3(_04430_ ), .ZN(_08057_ ) );
NAND3_X1 _16094_ ( .A1(_08057_ ), .A2(_07125_ ), .A3(_08050_ ), .ZN(_08058_ ) );
AOI22_X1 _16095_ ( .A1(_05206_ ), .A2(_07110_ ), .B1(\ID_EX_imm [10] ), .B2(_07114_ ), .ZN(_08059_ ) );
AOI21_X1 _16096_ ( .A(_07418_ ), .B1(_08058_ ), .B2(_08059_ ), .ZN(_08060_ ) );
OR2_X1 _16097_ ( .A1(_08060_ ), .A2(_04870_ ), .ZN(_08061_ ) );
NAND3_X1 _16098_ ( .A1(_07200_ ), .A2(_07610_ ), .A3(_07543_ ), .ZN(_08062_ ) );
NAND2_X1 _16099_ ( .A1(_07200_ ), .A2(_07212_ ), .ZN(_08063_ ) );
NAND2_X1 _16100_ ( .A1(_08062_ ), .A2(_08063_ ), .ZN(_08064_ ) );
NAND2_X1 _16101_ ( .A1(_08064_ ), .A2(_07827_ ), .ZN(_08065_ ) );
OR3_X1 _16102_ ( .A1(_07626_ ), .A2(_07461_ ), .A3(_07514_ ), .ZN(_08066_ ) );
OAI21_X1 _16103_ ( .A(_07275_ ), .B1(_07490_ ), .B2(_07482_ ), .ZN(_08067_ ) );
OAI21_X1 _16104_ ( .A(_07258_ ), .B1(_07640_ ), .B2(_07480_ ), .ZN(_08068_ ) );
AOI21_X1 _16105_ ( .A(_07478_ ), .B1(_08067_ ), .B2(_08068_ ), .ZN(_08069_ ) );
AOI21_X1 _16106_ ( .A(_07272_ ), .B1(_07830_ ), .B2(_07831_ ), .ZN(_08070_ ) );
OAI21_X1 _16107_ ( .A(_07630_ ), .B1(_08069_ ), .B2(_08070_ ), .ZN(_08071_ ) );
OAI211_X1 _16108_ ( .A(_08071_ ), .B(_07251_ ), .C1(_07620_ ), .C2(_07696_ ), .ZN(_08072_ ) );
AND2_X1 _16109_ ( .A1(_08066_ ), .A2(_08072_ ), .ZN(_08073_ ) );
AOI21_X1 _16110_ ( .A(_07805_ ), .B1(_08065_ ), .B2(_08073_ ), .ZN(_08074_ ) );
AOI21_X1 _16111_ ( .A(_07852_ ), .B1(_08066_ ), .B2(_08072_ ), .ZN(_08075_ ) );
OAI21_X1 _16112_ ( .A(_07697_ ), .B1(_07634_ ), .B2(_07635_ ), .ZN(_08076_ ) );
OAI211_X1 _16113_ ( .A(_08076_ ), .B(_07696_ ), .C1(_07844_ ), .C2(_07697_ ), .ZN(_08077_ ) );
OAI21_X1 _16114_ ( .A(_07920_ ), .B1(_07649_ ), .B2(_07650_ ), .ZN(_08078_ ) );
AND3_X1 _16115_ ( .A1(_08077_ ), .A2(_07799_ ), .A3(_08078_ ), .ZN(_08079_ ) );
NOR3_X1 _16116_ ( .A1(_08074_ ), .A2(_08075_ ), .A3(_08079_ ), .ZN(_08080_ ) );
AND3_X1 _16117_ ( .A1(_08041_ ), .A2(_04621_ ), .A3(_07335_ ), .ZN(_08081_ ) );
OR3_X1 _16118_ ( .A1(_08081_ ), .A2(_08042_ ), .A3(_07809_ ), .ZN(_08082_ ) );
AND2_X1 _16119_ ( .A1(_04620_ ), .A2(_07327_ ), .ZN(_08083_ ) );
NOR3_X1 _16120_ ( .A1(_04619_ ), .A2(_07308_ ), .A3(_07521_ ), .ZN(_08084_ ) );
AOI21_X1 _16121_ ( .A(_07657_ ), .B1(_04619_ ), .B2(_07308_ ), .ZN(_08085_ ) );
NOR3_X1 _16122_ ( .A1(_08083_ ), .A2(_08084_ ), .A3(_08085_ ), .ZN(_08086_ ) );
NAND3_X1 _16123_ ( .A1(_08080_ ), .A2(_08082_ ), .A3(_08086_ ), .ZN(_08087_ ) );
AOI21_X1 _16124_ ( .A(_08061_ ), .B1(_08087_ ), .B2(_07420_ ), .ZN(_08088_ ) );
BUF_X4 _16125_ ( .A(_06694_ ), .Z(_08089_ ) );
OAI21_X1 _16126_ ( .A(_08089_ ), .B1(_05203_ ), .B2(_04783_ ), .ZN(_08090_ ) );
OAI22_X1 _16127_ ( .A1(_08088_ ), .A2(_08090_ ), .B1(_06695_ ), .B2(_05218_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
OAI21_X1 _16128_ ( .A(_07424_ ), .B1(_06886_ ), .B2(_06887_ ), .ZN(_08091_ ) );
AOI21_X1 _16129_ ( .A(_04427_ ), .B1(_04454_ ), .B2(_04320_ ), .ZN(_08092_ ) );
XNOR2_X1 _16130_ ( .A(_08092_ ), .B(_04298_ ), .ZN(_08093_ ) );
NAND2_X1 _16131_ ( .A1(_08093_ ), .A2(_07126_ ), .ZN(_08094_ ) );
AOI22_X1 _16132_ ( .A1(_05232_ ), .A2(_07603_ ), .B1(\ID_EX_imm [9] ), .B2(_07539_ ), .ZN(_08095_ ) );
AOI21_X1 _16133_ ( .A(_07418_ ), .B1(_08094_ ), .B2(_08095_ ), .ZN(_08096_ ) );
OR2_X1 _16134_ ( .A1(_08096_ ), .A2(_07662_ ), .ZN(_08097_ ) );
NAND3_X1 _16135_ ( .A1(_07200_ ), .A2(_07205_ ), .A3(_07543_ ), .ZN(_08098_ ) );
OAI21_X1 _16136_ ( .A(_08063_ ), .B1(_08098_ ), .B2(_07212_ ), .ZN(_08099_ ) );
NAND2_X1 _16137_ ( .A1(_08099_ ), .A2(_07827_ ), .ZN(_08100_ ) );
OAI21_X1 _16138_ ( .A(_07283_ ), .B1(_07684_ ), .B2(_07514_ ), .ZN(_08101_ ) );
AOI21_X1 _16139_ ( .A(_07261_ ), .B1(_07877_ ), .B2(_07878_ ), .ZN(_08102_ ) );
OAI21_X1 _16140_ ( .A(_07274_ ), .B1(_07306_ ), .B2(_07310_ ), .ZN(_08103_ ) );
OAI21_X1 _16141_ ( .A(_07202_ ), .B1(_07309_ ), .B2(_07318_ ), .ZN(_08104_ ) );
AOI21_X1 _16142_ ( .A(_07206_ ), .B1(_08103_ ), .B2(_08104_ ), .ZN(_08105_ ) );
NOR2_X1 _16143_ ( .A1(_08102_ ), .A2(_08105_ ), .ZN(_08106_ ) );
NOR2_X1 _16144_ ( .A1(_08106_ ), .A2(_07322_ ), .ZN(_08107_ ) );
AND3_X1 _16145_ ( .A1(_07676_ ), .A2(_07679_ ), .A3(_07209_ ), .ZN(_08108_ ) );
OAI21_X1 _16146_ ( .A(_07250_ ), .B1(_08107_ ), .B2(_08108_ ), .ZN(_08109_ ) );
NAND2_X1 _16147_ ( .A1(_08101_ ), .A2(_08109_ ), .ZN(_08110_ ) );
AOI21_X1 _16148_ ( .A(_07804_ ), .B1(_08100_ ), .B2(_08110_ ), .ZN(_08111_ ) );
AND3_X1 _16149_ ( .A1(_08101_ ), .A2(_07407_ ), .A3(_08109_ ), .ZN(_08112_ ) );
OAI21_X1 _16150_ ( .A(_07630_ ), .B1(_07689_ ), .B2(_07690_ ), .ZN(_08113_ ) );
NAND3_X1 _16151_ ( .A1(_07277_ ), .A2(_07323_ ), .A3(_07916_ ), .ZN(_08114_ ) );
AOI21_X1 _16152_ ( .A(_07930_ ), .B1(_08113_ ), .B2(_08114_ ), .ZN(_08115_ ) );
OR3_X1 _16153_ ( .A1(_08111_ ), .A2(_08112_ ), .A3(_08115_ ), .ZN(_08116_ ) );
OAI21_X1 _16154_ ( .A(_04580_ ), .B1(_07369_ ), .B2(_07377_ ), .ZN(_08117_ ) );
INV_X1 _16155_ ( .A(_07333_ ), .ZN(_08118_ ) );
AND3_X1 _16156_ ( .A1(_08117_ ), .A2(_04586_ ), .A3(_08118_ ), .ZN(_08119_ ) );
AOI21_X1 _16157_ ( .A(_04586_ ), .B1(_08117_ ), .B2(_08118_ ), .ZN(_08120_ ) );
NOR3_X1 _16158_ ( .A1(_08119_ ), .A2(_08120_ ), .A3(_07808_ ), .ZN(_08121_ ) );
AOI22_X1 _16159_ ( .A1(_07332_ ), .A2(_07409_ ), .B1(_07334_ ), .B2(_07329_ ), .ZN(_08122_ ) );
OAI21_X1 _16160_ ( .A(_08122_ ), .B1(_04586_ ), .B2(_07753_ ), .ZN(_08123_ ) );
OR3_X1 _16161_ ( .A1(_08116_ ), .A2(_08121_ ), .A3(_08123_ ), .ZN(_08124_ ) );
BUF_X4 _16162_ ( .A(_07420_ ), .Z(_08125_ ) );
AOI21_X1 _16163_ ( .A(_08097_ ), .B1(_08124_ ), .B2(_08125_ ), .ZN(_08126_ ) );
NAND2_X1 _16164_ ( .A1(_05228_ ), .A2(_07663_ ), .ZN(_08127_ ) );
NAND2_X1 _16165_ ( .A1(_08127_ ), .A2(_07665_ ), .ZN(_08128_ ) );
OAI21_X1 _16166_ ( .A(_08091_ ), .B1(_08126_ ), .B2(_08128_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _16167_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_06606_ ), .ZN(_08129_ ) );
OAI211_X1 _16168_ ( .A(_06802_ ), .B(_08129_ ), .C1(_07083_ ), .C2(_06898_ ), .ZN(_08130_ ) );
AOI21_X1 _16169_ ( .A(_07600_ ), .B1(_04454_ ), .B2(_04320_ ), .ZN(_08131_ ) );
OAI21_X1 _16170_ ( .A(_08131_ ), .B1(_04320_ ), .B2(_04454_ ), .ZN(_08132_ ) );
AOI22_X1 _16171_ ( .A1(_05265_ ), .A2(_07603_ ), .B1(\ID_EX_imm [8] ), .B2(_07114_ ), .ZN(_08133_ ) );
AOI21_X1 _16172_ ( .A(_07418_ ), .B1(_08132_ ), .B2(_08133_ ), .ZN(_08134_ ) );
OR2_X1 _16173_ ( .A1(_08134_ ), .A2(_07662_ ), .ZN(_08135_ ) );
NOR2_X1 _16174_ ( .A1(_07134_ ), .A2(_07280_ ), .ZN(_08136_ ) );
INV_X1 _16175_ ( .A(_08136_ ), .ZN(_08137_ ) );
NAND4_X1 _16176_ ( .A1(_07914_ ), .A2(_07802_ ), .A3(_08137_ ), .A4(_07725_ ), .ZN(_08138_ ) );
OAI21_X1 _16177_ ( .A(_07283_ ), .B1(_07734_ ), .B2(_07514_ ), .ZN(_08139_ ) );
NAND3_X1 _16178_ ( .A1(_07728_ ), .A2(_07279_ ), .A3(_07731_ ), .ZN(_08140_ ) );
OAI21_X1 _16179_ ( .A(_07265_ ), .B1(_07640_ ), .B2(_07480_ ), .ZN(_08141_ ) );
OAI21_X1 _16180_ ( .A(_07258_ ), .B1(_07479_ ), .B2(_07468_ ), .ZN(_08142_ ) );
NAND2_X1 _16181_ ( .A1(_08141_ ), .A2(_08142_ ), .ZN(_08143_ ) );
NAND2_X1 _16182_ ( .A1(_08143_ ), .A2(_07272_ ), .ZN(_08144_ ) );
NAND3_X1 _16183_ ( .A1(_07922_ ), .A2(_07478_ ), .A3(_07923_ ), .ZN(_08145_ ) );
NAND3_X1 _16184_ ( .A1(_08144_ ), .A2(_08145_ ), .A3(_07477_ ), .ZN(_08146_ ) );
NAND3_X1 _16185_ ( .A1(_08140_ ), .A2(_07250_ ), .A3(_08146_ ), .ZN(_08147_ ) );
NAND2_X1 _16186_ ( .A1(_08139_ ), .A2(_08147_ ), .ZN(_08148_ ) );
AOI21_X1 _16187_ ( .A(_07805_ ), .B1(_08138_ ), .B2(_08148_ ), .ZN(_08149_ ) );
NAND2_X1 _16188_ ( .A1(_08117_ ), .A2(_07403_ ), .ZN(_08150_ ) );
AOI21_X1 _16189_ ( .A(_08150_ ), .B1(_04581_ ), .B2(_07378_ ), .ZN(_08151_ ) );
AND3_X1 _16190_ ( .A1(_08139_ ), .A2(_07407_ ), .A3(_08147_ ), .ZN(_08152_ ) );
NOR3_X1 _16191_ ( .A1(_04579_ ), .A2(_04679_ ), .A3(_07521_ ), .ZN(_08153_ ) );
OAI21_X1 _16192_ ( .A(_07433_ ), .B1(_07469_ ), .B2(_07473_ ), .ZN(_08154_ ) );
OAI211_X1 _16193_ ( .A(_08154_ ), .B(_07477_ ), .C1(_07273_ ), .C2(_07512_ ), .ZN(_08155_ ) );
OAI21_X1 _16194_ ( .A(_07279_ ), .B1(_07505_ ), .B2(_07301_ ), .ZN(_08156_ ) );
NAND3_X1 _16195_ ( .A1(_08155_ ), .A2(_07799_ ), .A3(_08156_ ), .ZN(_08157_ ) );
NAND2_X1 _16196_ ( .A1(_04580_ ), .A2(_07326_ ), .ZN(_08158_ ) );
OAI21_X1 _16197_ ( .A(_07329_ ), .B1(_04680_ ), .B2(_02938_ ), .ZN(_08159_ ) );
NAND3_X1 _16198_ ( .A1(_08157_ ), .A2(_08158_ ), .A3(_08159_ ), .ZN(_08160_ ) );
OR3_X1 _16199_ ( .A1(_08152_ ), .A2(_08153_ ), .A3(_08160_ ), .ZN(_08161_ ) );
OR3_X1 _16200_ ( .A1(_08149_ ), .A2(_08151_ ), .A3(_08161_ ), .ZN(_08162_ ) );
AOI21_X1 _16201_ ( .A(_08135_ ), .B1(_08162_ ), .B2(_08125_ ), .ZN(_08163_ ) );
OAI21_X1 _16202_ ( .A(_06994_ ), .B1(_05264_ ), .B2(_05663_ ), .ZN(_08164_ ) );
OAI21_X1 _16203_ ( .A(_08130_ ), .B1(_08163_ ), .B2(_08164_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
OR2_X1 _16204_ ( .A1(_05288_ ), .A2(_06700_ ), .ZN(_08165_ ) );
OR2_X1 _16205_ ( .A1(_04442_ ), .A2(_04445_ ), .ZN(_08166_ ) );
AOI21_X1 _16206_ ( .A(_04451_ ), .B1(_08166_ ), .B2(_04413_ ), .ZN(_08167_ ) );
INV_X1 _16207_ ( .A(_04367_ ), .ZN(_08168_ ) );
OR2_X1 _16208_ ( .A1(_08167_ ), .A2(_08168_ ), .ZN(_08169_ ) );
INV_X1 _16209_ ( .A(_04343_ ), .ZN(_08170_ ) );
AND3_X1 _16210_ ( .A1(_08169_ ), .A2(_08170_ ), .A3(_04365_ ), .ZN(_08171_ ) );
AOI21_X1 _16211_ ( .A(_08170_ ), .B1(_08169_ ), .B2(_04365_ ), .ZN(_08172_ ) );
OR3_X1 _16212_ ( .A1(_08171_ ), .A2(_08172_ ), .A3(_07599_ ), .ZN(_08173_ ) );
AOI22_X1 _16213_ ( .A1(_05292_ ), .A2(_07603_ ), .B1(\ID_EX_imm [7] ), .B2(_07114_ ), .ZN(_08174_ ) );
AOI21_X1 _16214_ ( .A(_07418_ ), .B1(_08173_ ), .B2(_08174_ ), .ZN(_08175_ ) );
OR2_X1 _16215_ ( .A1(_08175_ ), .A2(_07662_ ), .ZN(_08176_ ) );
NAND4_X1 _16216_ ( .A1(_07914_ ), .A2(_07802_ ), .A3(_07544_ ), .A4(_07725_ ), .ZN(_08177_ ) );
MUX2_X1 _16217_ ( .A(_07788_ ), .B(_07780_ ), .S(_07476_ ), .Z(_08178_ ) );
OR2_X1 _16218_ ( .A1(_08178_ ), .A2(_07249_ ), .ZN(_08179_ ) );
OR3_X1 _16219_ ( .A1(_08023_ ), .A2(_08024_ ), .A3(_07271_ ), .ZN(_08180_ ) );
NOR3_X1 _16220_ ( .A1(_07313_ ), .A2(_07265_ ), .A3(_07317_ ), .ZN(_08181_ ) );
NOR3_X1 _16221_ ( .A1(_07309_ ), .A2(_07318_ ), .A3(_07202_ ), .ZN(_08182_ ) );
NOR2_X1 _16222_ ( .A1(_08181_ ), .A2(_08182_ ), .ZN(_08183_ ) );
INV_X1 _16223_ ( .A(_08183_ ), .ZN(_08184_ ) );
OAI211_X1 _16224_ ( .A(_08180_ ), .B(_07477_ ), .C1(_07301_ ), .C2(_08184_ ), .ZN(_08185_ ) );
OAI211_X1 _16225_ ( .A(_08185_ ), .B(_07250_ ), .C1(_07578_ ), .C2(_07786_ ), .ZN(_08186_ ) );
NAND2_X1 _16226_ ( .A1(_08179_ ), .A2(_08186_ ), .ZN(_08187_ ) );
AOI21_X1 _16227_ ( .A(_07805_ ), .B1(_08177_ ), .B2(_08187_ ), .ZN(_08188_ ) );
AND3_X1 _16228_ ( .A1(_07363_ ), .A2(_07354_ ), .A3(_07368_ ), .ZN(_08189_ ) );
OAI21_X1 _16229_ ( .A(_04670_ ), .B1(_08189_ ), .B2(_07375_ ), .ZN(_08190_ ) );
INV_X1 _16230_ ( .A(_07371_ ), .ZN(_08191_ ) );
AND3_X1 _16231_ ( .A1(_08190_ ), .A2(_04672_ ), .A3(_08191_ ), .ZN(_08192_ ) );
AOI21_X1 _16232_ ( .A(_04672_ ), .B1(_08190_ ), .B2(_08191_ ), .ZN(_08193_ ) );
NOR3_X1 _16233_ ( .A1(_08192_ ), .A2(_08193_ ), .A3(_07808_ ), .ZN(_08194_ ) );
AND3_X1 _16234_ ( .A1(_08179_ ), .A2(_07406_ ), .A3(_08186_ ), .ZN(_08195_ ) );
AOI21_X1 _16235_ ( .A(_07524_ ), .B1(_04665_ ), .B2(_02912_ ), .ZN(_08196_ ) );
NOR3_X1 _16236_ ( .A1(_07793_ ), .A2(_07279_ ), .A3(_07930_ ), .ZN(_08197_ ) );
AND2_X1 _16237_ ( .A1(_04666_ ), .A2(_04506_ ), .ZN(_08198_ ) );
NOR3_X1 _16238_ ( .A1(_04665_ ), .A2(_02912_ ), .A3(_04420_ ), .ZN(_08199_ ) );
OR3_X1 _16239_ ( .A1(_08197_ ), .A2(_08198_ ), .A3(_08199_ ), .ZN(_08200_ ) );
OR3_X1 _16240_ ( .A1(_08195_ ), .A2(_08196_ ), .A3(_08200_ ), .ZN(_08201_ ) );
OR3_X1 _16241_ ( .A1(_08188_ ), .A2(_08194_ ), .A3(_08201_ ), .ZN(_08202_ ) );
AOI21_X1 _16242_ ( .A(_08176_ ), .B1(_08202_ ), .B2(_08125_ ), .ZN(_08203_ ) );
OAI21_X1 _16243_ ( .A(_06994_ ), .B1(_05295_ ), .B2(_05663_ ), .ZN(_08204_ ) );
OAI21_X1 _16244_ ( .A(_08165_ ), .B1(_08203_ ), .B2(_08204_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _16245_ ( .A1(_08167_ ), .A2(_08168_ ), .ZN(_08205_ ) );
NAND3_X1 _16246_ ( .A1(_08169_ ), .A2(_07126_ ), .A3(_08205_ ), .ZN(_08206_ ) );
NAND3_X1 _16247_ ( .A1(_05319_ ), .A2(_03428_ ), .A3(_07428_ ), .ZN(_08207_ ) );
NAND3_X1 _16248_ ( .A1(_07112_ ), .A2(\ID_EX_imm [6] ), .A3(_07109_ ), .ZN(_08208_ ) );
NAND3_X1 _16249_ ( .A1(_08206_ ), .A2(_08207_ ), .A3(_08208_ ), .ZN(_08209_ ) );
AOI21_X1 _16250_ ( .A(_05180_ ), .B1(_08209_ ), .B2(_07417_ ), .ZN(_08210_ ) );
AND4_X1 _16251_ ( .A1(_07544_ ), .A2(_07200_ ), .A3(_07827_ ), .A4(_07828_ ), .ZN(_08211_ ) );
MUX2_X1 _16252_ ( .A(_07975_ ), .B(_07837_ ), .S(_07477_ ), .Z(_08212_ ) );
NAND2_X1 _16253_ ( .A1(_08212_ ), .A2(_07284_ ), .ZN(_08213_ ) );
OAI211_X1 _16254_ ( .A(_07832_ ), .B(_07323_ ), .C1(_07833_ ), .C2(_07916_ ), .ZN(_08214_ ) );
OAI21_X1 _16255_ ( .A(_07292_ ), .B1(_07467_ ), .B2(_07471_ ), .ZN(_08215_ ) );
OAI21_X1 _16256_ ( .A(_07275_ ), .B1(_07479_ ), .B2(_07468_ ), .ZN(_08216_ ) );
AND3_X1 _16257_ ( .A1(_08215_ ), .A2(_07916_ ), .A3(_08216_ ), .ZN(_08217_ ) );
NAND3_X1 _16258_ ( .A1(_08067_ ), .A2(_08068_ ), .A3(_07650_ ), .ZN(_08218_ ) );
NAND2_X1 _16259_ ( .A1(_08218_ ), .A2(_07630_ ), .ZN(_08219_ ) );
OAI211_X1 _16260_ ( .A(_08214_ ), .B(_07251_ ), .C1(_08217_ ), .C2(_08219_ ), .ZN(_08220_ ) );
NAND2_X1 _16261_ ( .A1(_08213_ ), .A2(_08220_ ), .ZN(_08221_ ) );
OAI21_X1 _16262_ ( .A(_07131_ ), .B1(_08211_ ), .B2(_08221_ ), .ZN(_08222_ ) );
OR3_X1 _16263_ ( .A1(_08189_ ), .A2(_04670_ ), .A3(_07375_ ), .ZN(_08223_ ) );
NAND3_X1 _16264_ ( .A1(_08223_ ), .A2(_07404_ ), .A3(_08190_ ), .ZN(_08224_ ) );
AOI21_X1 _16265_ ( .A(_07524_ ), .B1(_04669_ ), .B2(_07314_ ), .ZN(_08225_ ) );
NOR3_X1 _16266_ ( .A1(_07845_ ), .A2(_07514_ ), .A3(_07930_ ), .ZN(_08226_ ) );
AND2_X1 _16267_ ( .A1(_04670_ ), .A2(_04506_ ), .ZN(_08227_ ) );
NOR3_X1 _16268_ ( .A1(_04669_ ), .A2(_07314_ ), .A3(_04420_ ), .ZN(_08228_ ) );
OR3_X1 _16269_ ( .A1(_08226_ ), .A2(_08227_ ), .A3(_08228_ ), .ZN(_08229_ ) );
AOI211_X1 _16270_ ( .A(_08225_ ), .B(_08229_ ), .C1(_08221_ ), .C2(_07408_ ), .ZN(_08230_ ) );
AND3_X1 _16271_ ( .A1(_08222_ ), .A2(_08224_ ), .A3(_08230_ ), .ZN(_08231_ ) );
OAI21_X1 _16272_ ( .A(_08210_ ), .B1(_08231_ ), .B2(_07419_ ), .ZN(_08232_ ) );
OR2_X1 _16273_ ( .A1(_05318_ ), .A2(_04831_ ), .ZN(_08233_ ) );
NAND3_X1 _16274_ ( .A1(_08232_ ), .A2(_06695_ ), .A3(_08233_ ), .ZN(_08234_ ) );
NAND2_X1 _16275_ ( .A1(_06928_ ), .A2(_06706_ ), .ZN(_08235_ ) );
NAND2_X1 _16276_ ( .A1(_08234_ ), .A2(_08235_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
NOR2_X1 _16277_ ( .A1(_06939_ ), .A2(_06940_ ), .ZN(_08236_ ) );
AND2_X1 _16278_ ( .A1(_05332_ ), .A2(_02415_ ), .ZN(_08237_ ) );
NOR3_X1 _16279_ ( .A1(_07366_ ), .A2(_07367_ ), .A3(_07753_ ), .ZN(_08238_ ) );
AND4_X1 _16280_ ( .A1(_07208_ ), .A2(_07199_ ), .A3(_07212_ ), .A4(_07827_ ), .ZN(_08239_ ) );
NAND2_X1 _16281_ ( .A1(_07248_ ), .A2(_07283_ ), .ZN(_08240_ ) );
NOR3_X1 _16282_ ( .A1(_07274_ ), .A2(_07315_ ), .A3(_07268_ ), .ZN(_08241_ ) );
NOR3_X1 _16283_ ( .A1(_07313_ ), .A2(_07317_ ), .A3(_07257_ ), .ZN(_08242_ ) );
OAI21_X1 _16284_ ( .A(_07271_ ), .B1(_08241_ ), .B2(_08242_ ), .ZN(_08243_ ) );
NAND3_X1 _16285_ ( .A1(_08103_ ), .A2(_08104_ ), .A3(_07444_ ), .ZN(_08244_ ) );
NAND3_X1 _16286_ ( .A1(_08243_ ), .A2(_07476_ ), .A3(_08244_ ), .ZN(_08245_ ) );
OAI211_X1 _16287_ ( .A(_07249_ ), .B(_08245_ ), .C1(_07881_ ), .C2(_07476_ ), .ZN(_08246_ ) );
NAND2_X1 _16288_ ( .A1(_08240_ ), .A2(_08246_ ), .ZN(_08247_ ) );
OAI21_X1 _16289_ ( .A(_07130_ ), .B1(_08239_ ), .B2(_08247_ ), .ZN(_08248_ ) );
NAND2_X1 _16290_ ( .A1(_08247_ ), .A2(_07406_ ), .ZN(_08249_ ) );
NAND2_X1 _16291_ ( .A1(_08248_ ), .A2(_08249_ ), .ZN(_08250_ ) );
OAI22_X1 _16292_ ( .A1(_07372_ ), .A2(_04420_ ), .B1(_07367_ ), .B2(_07523_ ), .ZN(_08251_ ) );
NOR3_X1 _16293_ ( .A1(_07278_ ), .A2(_07323_ ), .A3(_07930_ ), .ZN(_08252_ ) );
OR4_X1 _16294_ ( .A1(_08238_ ), .A2(_08250_ ), .A3(_08251_ ), .A4(_08252_ ), .ZN(_08253_ ) );
NAND2_X1 _16295_ ( .A1(_07363_ ), .A2(_07354_ ), .ZN(_00304_ ) );
NOR2_X1 _16296_ ( .A1(_00304_ ), .A2(_07365_ ), .ZN(_00305_ ) );
NOR3_X1 _16297_ ( .A1(_00305_ ), .A2(_04626_ ), .A3(_07373_ ), .ZN(_00306_ ) );
NOR2_X1 _16298_ ( .A1(_00306_ ), .A2(_07808_ ), .ZN(_00307_ ) );
OAI21_X1 _16299_ ( .A(_04626_ ), .B1(_00305_ ), .B2(_07373_ ), .ZN(_00308_ ) );
AND2_X1 _16300_ ( .A1(_00307_ ), .A2(_00308_ ), .ZN(_00309_ ) );
OAI21_X1 _16301_ ( .A(_07420_ ), .B1(_08253_ ), .B2(_00309_ ), .ZN(_00310_ ) );
AND2_X1 _16302_ ( .A1(_08166_ ), .A2(_04390_ ), .ZN(_00311_ ) );
OR3_X1 _16303_ ( .A1(_00311_ ), .A2(_04412_ ), .A3(_04448_ ), .ZN(_00312_ ) );
OAI21_X1 _16304_ ( .A(_04412_ ), .B1(_00311_ ), .B2(_04448_ ), .ZN(_00313_ ) );
NAND3_X1 _16305_ ( .A1(_00312_ ), .A2(_07125_ ), .A3(_00313_ ), .ZN(_00314_ ) );
AOI22_X1 _16306_ ( .A1(_05336_ ), .A2(_07110_ ), .B1(\ID_EX_imm [5] ), .B2(_07114_ ), .ZN(_00315_ ) );
AOI21_X1 _16307_ ( .A(_07418_ ), .B1(_00314_ ), .B2(_00315_ ), .ZN(_00316_ ) );
NOR2_X1 _16308_ ( .A1(_00316_ ), .A2(_04870_ ), .ZN(_00317_ ) );
AOI21_X1 _16309_ ( .A(_08237_ ), .B1(_00310_ ), .B2(_00317_ ), .ZN(_00318_ ) );
MUX2_X1 _16310_ ( .A(_08236_ ), .B(_00318_ ), .S(_06700_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
NOR3_X1 _16311_ ( .A1(_04442_ ), .A2(_04390_ ), .A3(_04445_ ), .ZN(_00319_ ) );
NOR3_X1 _16312_ ( .A1(_00311_ ), .A2(_00319_ ), .A3(_07600_ ), .ZN(_00320_ ) );
OAI22_X1 _16313_ ( .A1(_05372_ ), .A2(_07111_ ), .B1(_02856_ ), .B2(_07115_ ), .ZN(_00321_ ) );
OAI21_X1 _16314_ ( .A(_07417_ ), .B1(_00320_ ), .B2(_00321_ ), .ZN(_00322_ ) );
AND2_X1 _16315_ ( .A1(_00322_ ), .A2(_04782_ ), .ZN(_00323_ ) );
NAND4_X1 _16316_ ( .A1(_07914_ ), .A2(_07434_ ), .A3(_07544_ ), .A4(_07827_ ), .ZN(_00324_ ) );
AND2_X1 _16317_ ( .A1(_07460_ ), .A2(_07688_ ), .ZN(_00325_ ) );
AND3_X1 _16318_ ( .A1(_08141_ ), .A2(_08142_ ), .A3(_07478_ ), .ZN(_00326_ ) );
NOR3_X1 _16319_ ( .A1(_07507_ ), .A2(_07265_ ), .A3(_07470_ ), .ZN(_00327_ ) );
NOR3_X1 _16320_ ( .A1(_07467_ ), .A2(_07472_ ), .A3(_07471_ ), .ZN(_00328_ ) );
NOR2_X1 _16321_ ( .A1(_00327_ ), .A2(_00328_ ), .ZN(_00329_ ) );
INV_X1 _16322_ ( .A(_00329_ ), .ZN(_00330_ ) );
AOI211_X1 _16323_ ( .A(_07279_ ), .B(_00326_ ), .C1(_00330_ ), .C2(_07916_ ), .ZN(_00331_ ) );
AOI211_X1 _16324_ ( .A(_07688_ ), .B(_00331_ ), .C1(_07280_ ), .C2(_07925_ ), .ZN(_00332_ ) );
NOR2_X1 _16325_ ( .A1(_00325_ ), .A2(_00332_ ), .ZN(_00333_ ) );
AOI21_X1 _16326_ ( .A(_07805_ ), .B1(_00324_ ), .B2(_00333_ ), .ZN(_00334_ ) );
AOI21_X1 _16327_ ( .A(_07808_ ), .B1(_00304_ ), .B2(_07365_ ), .ZN(_00335_ ) );
OAI21_X1 _16328_ ( .A(_00335_ ), .B1(_07365_ ), .B2(_00304_ ), .ZN(_00336_ ) );
AND2_X1 _16329_ ( .A1(_07464_ ), .A2(_02860_ ), .ZN(_00337_ ) );
OAI221_X1 _16330_ ( .A(_00336_ ), .B1(_00337_ ), .B2(_07657_ ), .C1(_00333_ ), .C2(_07852_ ), .ZN(_00338_ ) );
OR3_X1 _16331_ ( .A1(_07513_ ), .A2(_07280_ ), .A3(_07930_ ), .ZN(_00339_ ) );
OAI221_X1 _16332_ ( .A(_00339_ ), .B1(_07374_ ), .B2(_07521_ ), .C1(_07365_ ), .C2(_07753_ ), .ZN(_00340_ ) );
NOR3_X1 _16333_ ( .A1(_00334_ ), .A2(_00338_ ), .A3(_00340_ ), .ZN(_00341_ ) );
OAI21_X1 _16334_ ( .A(_00323_ ), .B1(_00341_ ), .B2(_07419_ ), .ZN(_00342_ ) );
NAND2_X1 _16335_ ( .A1(_05370_ ), .A2(_07663_ ), .ZN(_00343_ ) );
NAND3_X1 _16336_ ( .A1(_00342_ ), .A2(_06695_ ), .A3(_00343_ ), .ZN(_00344_ ) );
OAI211_X1 _16337_ ( .A(_07424_ ), .B(_06952_ ), .C1(_06822_ ), .C2(_05362_ ), .ZN(_00345_ ) );
NAND2_X1 _16338_ ( .A1(_00344_ ), .A2(_00345_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
OR2_X1 _16339_ ( .A1(_04439_ ), .A2(_04441_ ), .ZN(_00346_ ) );
INV_X1 _16340_ ( .A(_04443_ ), .ZN(_00347_ ) );
AND3_X1 _16341_ ( .A1(_00346_ ), .A2(_04440_ ), .A3(_00347_ ), .ZN(_00348_ ) );
AOI21_X1 _16342_ ( .A(_04440_ ), .B1(_00346_ ), .B2(_00347_ ), .ZN(_00349_ ) );
OR3_X1 _16343_ ( .A1(_00348_ ), .A2(_00349_ ), .A3(_07600_ ), .ZN(_00350_ ) );
AOI22_X1 _16344_ ( .A1(_05388_ ), .A2(_07428_ ), .B1(\ID_EX_imm [3] ), .B2(_07539_ ), .ZN(_00351_ ) );
AOI21_X1 _16345_ ( .A(_07531_ ), .B1(_00350_ ), .B2(_00351_ ), .ZN(_00352_ ) );
NOR2_X1 _16346_ ( .A1(_00352_ ), .A2(_05180_ ), .ZN(_00353_ ) );
NAND4_X1 _16347_ ( .A1(_07914_ ), .A2(_07543_ ), .A3(_07544_ ), .A4(_07827_ ), .ZN(_00354_ ) );
NOR2_X1 _16348_ ( .A1(_07315_ ), .A2(_07268_ ), .ZN(_00355_ ) );
NOR2_X1 _16349_ ( .A1(_07256_ ), .A2(_07263_ ), .ZN(_00356_ ) );
MUX2_X1 _16350_ ( .A(_00355_ ), .B(_00356_ ), .S(_07257_ ), .Z(_00357_ ) );
AND2_X1 _16351_ ( .A1(_00357_ ), .A2(_07261_ ), .ZN(_00358_ ) );
AOI211_X1 _16352_ ( .A(_07322_ ), .B(_00358_ ), .C1(_07650_ ), .C2(_08184_ ), .ZN(_00359_ ) );
AND3_X1 _16353_ ( .A1(_08025_ ), .A2(_07322_ ), .A3(_08026_ ), .ZN(_00360_ ) );
OR3_X1 _16354_ ( .A1(_00359_ ), .A2(_07283_ ), .A3(_00360_ ), .ZN(_00361_ ) );
NAND2_X1 _16355_ ( .A1(_07559_ ), .A2(_07688_ ), .ZN(_00362_ ) );
AND2_X1 _16356_ ( .A1(_00361_ ), .A2(_00362_ ), .ZN(_00363_ ) );
AOI21_X1 _16357_ ( .A(_07805_ ), .B1(_00354_ ), .B2(_00363_ ), .ZN(_00364_ ) );
NOR2_X1 _16358_ ( .A1(_07362_ ), .A2(_04656_ ), .ZN(_00365_ ) );
OAI21_X1 _16359_ ( .A(_04636_ ), .B1(_00365_ ), .B2(_07355_ ), .ZN(_00366_ ) );
OAI221_X1 _16360_ ( .A(_07356_ ), .B1(_04657_ ), .B2(_04658_ ), .C1(_07362_ ), .C2(_04656_ ), .ZN(_00367_ ) );
AND3_X1 _16361_ ( .A1(_00366_ ), .A2(_07403_ ), .A3(_00367_ ), .ZN(_00368_ ) );
AND3_X1 _16362_ ( .A1(_07589_ ), .A2(_07477_ ), .A3(_07799_ ), .ZN(_00369_ ) );
AOI221_X4 _16363_ ( .A(_00369_ ), .B1(_04657_ ), .B2(_04419_ ), .C1(_04636_ ), .C2(_04506_ ), .ZN(_00370_ ) );
OAI221_X1 _16364_ ( .A(_00370_ ), .B1(_04658_ ), .B2(_07657_ ), .C1(_00363_ ), .C2(_07852_ ), .ZN(_00371_ ) );
NOR3_X1 _16365_ ( .A1(_00364_ ), .A2(_00368_ ), .A3(_00371_ ), .ZN(_00372_ ) );
OAI21_X1 _16366_ ( .A(_00353_ ), .B1(_00372_ ), .B2(_07419_ ), .ZN(_00373_ ) );
NAND3_X1 _16367_ ( .A1(_05383_ ), .A2(\ID_EX_typ [7] ), .A3(_02413_ ), .ZN(_00374_ ) );
NAND3_X1 _16368_ ( .A1(_00373_ ), .A2(_07665_ ), .A3(_00374_ ), .ZN(_00375_ ) );
NAND3_X1 _16369_ ( .A1(_05364_ ), .A2(_05365_ ), .A3(_06579_ ), .ZN(_00376_ ) );
AND3_X1 _16370_ ( .A1(_06716_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_04896_ ), .ZN(_00377_ ) );
INV_X1 _16371_ ( .A(_00377_ ), .ZN(_00378_ ) );
NAND3_X1 _16372_ ( .A1(_06787_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_04991_ ), .ZN(_00379_ ) );
NAND3_X1 _16373_ ( .A1(_06787_ ), .A2(\mtvec [3] ), .A3(_04987_ ), .ZN(_00380_ ) );
NAND4_X1 _16374_ ( .A1(_05456_ ), .A2(_04896_ ), .A3(\mepc [3] ), .A4(_04992_ ), .ZN(_00381_ ) );
NAND4_X1 _16375_ ( .A1(_00378_ ), .A2(_00379_ ), .A3(_00380_ ), .A4(_00381_ ), .ZN(_00382_ ) );
OAI211_X1 _16376_ ( .A(_07424_ ), .B(_00376_ ), .C1(_06822_ ), .C2(_00382_ ), .ZN(_00383_ ) );
NAND2_X1 _16377_ ( .A1(_00375_ ), .A2(_00383_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
OAI21_X1 _16378_ ( .A(_07424_ ), .B1(_06973_ ), .B2(_06974_ ), .ZN(_00384_ ) );
NAND2_X1 _16379_ ( .A1(_04439_ ), .A2(_04441_ ), .ZN(_00385_ ) );
NAND3_X1 _16380_ ( .A1(_00346_ ), .A2(_07125_ ), .A3(_00385_ ), .ZN(_00386_ ) );
AOI22_X1 _16381_ ( .A1(_05414_ ), .A2(_07603_ ), .B1(\ID_EX_imm [2] ), .B2(_07114_ ), .ZN(_00387_ ) );
AOI21_X1 _16382_ ( .A(_07418_ ), .B1(_00386_ ), .B2(_00387_ ), .ZN(_00388_ ) );
OR2_X1 _16383_ ( .A1(_00388_ ), .A2(_07662_ ), .ZN(_00389_ ) );
NAND2_X1 _16384_ ( .A1(_07627_ ), .A2(_07688_ ), .ZN(_00390_ ) );
NOR3_X1 _16385_ ( .A1(_07507_ ), .A2(_07470_ ), .A3(_07258_ ), .ZN(_00391_ ) );
NOR2_X1 _16386_ ( .A1(_07506_ ), .A2(_07510_ ), .ZN(_00392_ ) );
AOI211_X1 _16387_ ( .A(_07478_ ), .B(_00391_ ), .C1(_07304_ ), .C2(_00392_ ), .ZN(_00393_ ) );
AOI21_X1 _16388_ ( .A(_07433_ ), .B1(_08215_ ), .B2(_08216_ ), .ZN(_00394_ ) );
OAI21_X1 _16389_ ( .A(_07578_ ), .B1(_00393_ ), .B2(_00394_ ), .ZN(_00395_ ) );
OAI21_X1 _16390_ ( .A(_07279_ ), .B1(_08069_ ), .B2(_08070_ ), .ZN(_00396_ ) );
NAND3_X1 _16391_ ( .A1(_00395_ ), .A2(_07461_ ), .A3(_00396_ ), .ZN(_00397_ ) );
AOI21_X1 _16392_ ( .A(_07852_ ), .B1(_00390_ ), .B2(_00397_ ), .ZN(_00398_ ) );
NOR4_X1 _16393_ ( .A1(_07649_ ), .A2(_07688_ ), .A3(_07323_ ), .A4(_07650_ ), .ZN(_00399_ ) );
AND2_X1 _16394_ ( .A1(_07186_ ), .A2(_07543_ ), .ZN(_00400_ ) );
NAND4_X1 _16395_ ( .A1(_00400_ ), .A2(_07610_ ), .A3(_07544_ ), .A4(_07827_ ), .ZN(_00401_ ) );
NAND3_X1 _16396_ ( .A1(_00401_ ), .A2(_00397_ ), .A3(_00390_ ), .ZN(_00402_ ) );
AOI221_X4 _16397_ ( .A(_00398_ ), .B1(_07254_ ), .B2(_00399_ ), .C1(_00402_ ), .C2(_07130_ ), .ZN(_00403_ ) );
AOI21_X1 _16398_ ( .A(_07809_ ), .B1(_07362_ ), .B2(_04656_ ), .ZN(_00404_ ) );
OAI21_X1 _16399_ ( .A(_00404_ ), .B1(_04656_ ), .B2(_07362_ ), .ZN(_00405_ ) );
AOI21_X1 _16400_ ( .A(_07524_ ), .B1(_07697_ ), .B2(_04108_ ), .ZN(_00406_ ) );
AOI221_X4 _16401_ ( .A(_00406_ ), .B1(_07355_ ), .B2(_04419_ ), .C1(_04655_ ), .C2(_07326_ ), .ZN(_00407_ ) );
NAND3_X1 _16402_ ( .A1(_00403_ ), .A2(_00405_ ), .A3(_00407_ ), .ZN(_00408_ ) );
AOI21_X1 _16403_ ( .A(_00389_ ), .B1(_00408_ ), .B2(_08125_ ), .ZN(_00409_ ) );
OAI21_X1 _16404_ ( .A(_08089_ ), .B1(_05453_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00410_ ) );
OAI21_X1 _16405_ ( .A(_00384_ ), .B1(_00409_ ), .B2(_00410_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
OAI211_X1 _16406_ ( .A(_06802_ ), .B(_06989_ ), .C1(_06822_ ), .C2(_06985_ ), .ZN(_00411_ ) );
NOR2_X1 _16407_ ( .A1(_04793_ ), .A2(_07111_ ), .ZN(_00412_ ) );
AND2_X1 _16408_ ( .A1(_08010_ ), .A2(_03870_ ), .ZN(_00413_ ) );
NOR2_X1 _16409_ ( .A1(_04750_ ), .A2(_03869_ ), .ZN(_00414_ ) );
OR3_X1 _16410_ ( .A1(_00413_ ), .A2(_00414_ ), .A3(_03892_ ), .ZN(_00415_ ) );
OAI21_X1 _16411_ ( .A(_03892_ ), .B1(_00413_ ), .B2(_00414_ ), .ZN(_00416_ ) );
AND3_X1 _16412_ ( .A1(_00415_ ), .A2(_07125_ ), .A3(_00416_ ), .ZN(_00417_ ) );
AND3_X1 _16413_ ( .A1(_07112_ ), .A2(\ID_EX_imm [29] ), .A3(_07109_ ), .ZN(_00418_ ) );
NOR3_X1 _16414_ ( .A1(_00412_ ), .A2(_00417_ ), .A3(_00418_ ), .ZN(_00419_ ) );
AOI21_X1 _16415_ ( .A(_05495_ ), .B1(_00419_ ), .B2(_05672_ ), .ZN(_00420_ ) );
OR3_X1 _16416_ ( .A1(_07965_ ), .A2(_04525_ ), .A3(_07967_ ), .ZN(_00421_ ) );
OAI21_X1 _16417_ ( .A(_04525_ ), .B1(_07965_ ), .B2(_07967_ ), .ZN(_00422_ ) );
NAND3_X1 _16418_ ( .A1(_00421_ ), .A2(_07404_ ), .A3(_00422_ ), .ZN(_00423_ ) );
AOI22_X1 _16419_ ( .A1(_04525_ ), .A2(_07327_ ), .B1(_07970_ ), .B2(_07329_ ), .ZN(_00424_ ) );
NAND3_X1 _16420_ ( .A1(_04524_ ), .A2(_03276_ ), .A3(_07409_ ), .ZN(_00425_ ) );
AND2_X1 _16421_ ( .A1(_00424_ ), .A2(_00425_ ), .ZN(_00426_ ) );
NOR4_X1 _16422_ ( .A1(_07170_ ), .A2(_07198_ ), .A3(_07138_ ), .A4(_07872_ ), .ZN(_00427_ ) );
AND2_X1 _16423_ ( .A1(_07200_ ), .A2(_07725_ ), .ZN(_00428_ ) );
AOI21_X1 _16424_ ( .A(_00427_ ), .B1(_00428_ ), .B2(_07802_ ), .ZN(_00429_ ) );
NAND2_X1 _16425_ ( .A1(_07874_ ), .A2(_07560_ ), .ZN(_00430_ ) );
AOI21_X1 _16426_ ( .A(_07805_ ), .B1(_00429_ ), .B2(_00430_ ), .ZN(_00431_ ) );
OAI21_X1 _16427_ ( .A(_07284_ ), .B1(_07888_ ), .B2(_07889_ ), .ZN(_00432_ ) );
OR3_X1 _16428_ ( .A1(_07230_ ), .A2(_07235_ ), .A3(_07258_ ), .ZN(_00433_ ) );
OR3_X1 _16429_ ( .A1(_07275_ ), .A2(_07236_ ), .A3(_07226_ ), .ZN(_00434_ ) );
AOI21_X1 _16430_ ( .A(_07273_ ), .B1(_00433_ ), .B2(_00434_ ), .ZN(_00435_ ) );
OAI21_X1 _16431_ ( .A(_07286_ ), .B1(_07217_ ), .B2(_07223_ ), .ZN(_00436_ ) );
OAI21_X1 _16432_ ( .A(_07292_ ), .B1(_07218_ ), .B2(_07244_ ), .ZN(_00437_ ) );
AND3_X1 _16433_ ( .A1(_00436_ ), .A2(_00437_ ), .A3(_07433_ ), .ZN(_00438_ ) );
OR3_X1 _16434_ ( .A1(_00435_ ), .A2(_00438_ ), .A3(_07514_ ), .ZN(_00439_ ) );
OAI211_X1 _16435_ ( .A(_00439_ ), .B(_07560_ ), .C1(_07638_ ), .C2(_07303_ ), .ZN(_00440_ ) );
AOI21_X1 _16436_ ( .A(_07255_ ), .B1(_00432_ ), .B2(_00440_ ), .ZN(_00441_ ) );
AND3_X1 _16437_ ( .A1(_07874_ ), .A2(_07560_ ), .A3(_07407_ ), .ZN(_00442_ ) );
NOR3_X1 _16438_ ( .A1(_00431_ ), .A2(_00441_ ), .A3(_00442_ ), .ZN(_00443_ ) );
NAND3_X1 _16439_ ( .A1(_00423_ ), .A2(_00426_ ), .A3(_00443_ ), .ZN(_00444_ ) );
AOI21_X1 _16440_ ( .A(_00420_ ), .B1(_00444_ ), .B2(_08125_ ), .ZN(_00445_ ) );
OAI21_X1 _16441_ ( .A(_08089_ ), .B1(_04821_ ), .B2(_05663_ ), .ZN(_00446_ ) );
OAI21_X1 _16442_ ( .A(_00411_ ), .B1(_00445_ ), .B2(_00446_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
NAND3_X1 _16443_ ( .A1(_06997_ ), .A2(_06706_ ), .A3(_07002_ ), .ZN(_00447_ ) );
OAI21_X1 _16444_ ( .A(_07125_ ), .B1(_04057_ ), .B2(_04082_ ), .ZN(_00448_ ) );
OAI22_X1 _16445_ ( .A1(_04438_ ), .A2(_00448_ ), .B1(_02780_ ), .B2(_07115_ ), .ZN(_00449_ ) );
AOI21_X1 _16446_ ( .A(_00449_ ), .B1(_05434_ ), .B2(_07428_ ), .ZN(_00450_ ) );
AOI21_X1 _16447_ ( .A(_05495_ ), .B1(_00450_ ), .B2(_05672_ ), .ZN(_00451_ ) );
NOR4_X1 _16448_ ( .A1(_08098_ ), .A2(_07187_ ), .A3(_07210_ ), .A4(_07138_ ), .ZN(_00452_ ) );
NAND2_X1 _16449_ ( .A1(_07685_ ), .A2(_07284_ ), .ZN(_00453_ ) );
OAI21_X1 _16450_ ( .A(_07304_ ), .B1(_07259_ ), .B2(_07276_ ), .ZN(_00454_ ) );
OAI211_X1 _16451_ ( .A(_00454_ ), .B(_07273_ ), .C1(_00356_ ), .C2(_07304_ ), .ZN(_00455_ ) );
OAI21_X1 _16452_ ( .A(_07650_ ), .B1(_08241_ ), .B2(_08242_ ), .ZN(_00456_ ) );
NAND3_X1 _16453_ ( .A1(_00455_ ), .A2(_00456_ ), .A3(_07630_ ), .ZN(_00457_ ) );
OAI211_X1 _16454_ ( .A(_00457_ ), .B(_07251_ ), .C1(_08106_ ), .C2(_07696_ ), .ZN(_00458_ ) );
NAND2_X1 _16455_ ( .A1(_00453_ ), .A2(_00458_ ), .ZN(_00459_ ) );
OAI21_X1 _16456_ ( .A(_07131_ ), .B1(_00452_ ), .B2(_00459_ ), .ZN(_00460_ ) );
OAI21_X1 _16457_ ( .A(_07403_ ), .B1(_04649_ ), .B2(_07360_ ), .ZN(_00461_ ) );
OR2_X1 _16458_ ( .A1(_00461_ ), .A2(_07361_ ), .ZN(_00462_ ) );
NAND2_X1 _16459_ ( .A1(_00459_ ), .A2(_07408_ ), .ZN(_00463_ ) );
AND4_X1 _16460_ ( .A1(_07251_ ), .A2(_07696_ ), .A3(_07697_ ), .A4(_07277_ ), .ZN(_00464_ ) );
NAND2_X1 _16461_ ( .A1(_00464_ ), .A2(_07254_ ), .ZN(_00465_ ) );
NAND2_X1 _16462_ ( .A1(_07357_ ), .A2(_07409_ ), .ZN(_00466_ ) );
AOI22_X1 _16463_ ( .A1(_04649_ ), .A2(_07326_ ), .B1(_07359_ ), .B2(_07329_ ), .ZN(_00467_ ) );
AND4_X1 _16464_ ( .A1(_00463_ ), .A2(_00465_ ), .A3(_00466_ ), .A4(_00467_ ), .ZN(_00468_ ) );
NAND3_X1 _16465_ ( .A1(_00460_ ), .A2(_00462_ ), .A3(_00468_ ), .ZN(_00469_ ) );
AOI21_X1 _16466_ ( .A(_00451_ ), .B1(_00469_ ), .B2(_08125_ ), .ZN(_00470_ ) );
OAI21_X1 _16467_ ( .A(_08089_ ), .B1(_05453_ ), .B2(\ID_EX_pc [1] ), .ZN(_00471_ ) );
OAI21_X1 _16468_ ( .A(_00447_ ), .B1(_00470_ ), .B2(_00471_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
NOR3_X1 _16469_ ( .A1(_04749_ ), .A2(_04760_ ), .A3(_07415_ ), .ZN(_00472_ ) );
NAND3_X1 _16470_ ( .A1(_07112_ ), .A2(\ID_EX_imm [0] ), .A3(_07109_ ), .ZN(_00473_ ) );
OAI21_X1 _16471_ ( .A(_00473_ ), .B1(_07111_ ), .B2(_05489_ ), .ZN(_00474_ ) );
AOI21_X1 _16472_ ( .A(_07600_ ), .B1(_04082_ ), .B2(_04083_ ), .ZN(_00475_ ) );
NOR3_X1 _16473_ ( .A1(_00472_ ), .A2(_00474_ ), .A3(_00475_ ), .ZN(_00476_ ) );
OAI211_X1 _16474_ ( .A(_04757_ ), .B(_04761_ ), .C1(_07174_ ), .C2(_04758_ ), .ZN(_00477_ ) );
NOR3_X1 _16475_ ( .A1(_04749_ ), .A2(_04754_ ), .A3(_00477_ ), .ZN(_00478_ ) );
AND4_X1 _16476_ ( .A1(_07254_ ), .A2(_07696_ ), .A3(_07461_ ), .A4(_07745_ ), .ZN(_00479_ ) );
NOR2_X1 _16477_ ( .A1(_00478_ ), .A2(_00479_ ), .ZN(_00480_ ) );
NOR4_X1 _16478_ ( .A1(_07170_ ), .A2(_07185_ ), .A3(_04661_ ), .A4(_07182_ ), .ZN(_00481_ ) );
OR2_X1 _16479_ ( .A1(_07735_ ), .A2(_07250_ ), .ZN(_00482_ ) );
NAND3_X1 _16480_ ( .A1(_08144_ ), .A2(_08145_ ), .A3(_07279_ ), .ZN(_00483_ ) );
NOR3_X1 _16481_ ( .A1(_07506_ ), .A2(_07472_ ), .A3(_07510_ ), .ZN(_00484_ ) );
AND2_X1 _16482_ ( .A1(_07204_ ), .A2(_04650_ ), .ZN(_00485_ ) );
NOR3_X1 _16483_ ( .A1(_00485_ ), .A2(_07265_ ), .A3(_07509_ ), .ZN(_00486_ ) );
OR3_X1 _16484_ ( .A1(_00484_ ), .A2(_00486_ ), .A3(_07206_ ), .ZN(_00487_ ) );
OAI21_X1 _16485_ ( .A(_00487_ ), .B1(_07273_ ), .B2(_00330_ ), .ZN(_00488_ ) );
OAI211_X1 _16486_ ( .A(_07461_ ), .B(_00483_ ), .C1(_00488_ ), .C2(_07514_ ), .ZN(_00489_ ) );
NAND2_X1 _16487_ ( .A1(_00482_ ), .A2(_00489_ ), .ZN(_00490_ ) );
INV_X1 _16488_ ( .A(_00490_ ), .ZN(_00491_ ) );
OAI21_X1 _16489_ ( .A(_07130_ ), .B1(_00481_ ), .B2(_00491_ ), .ZN(_00492_ ) );
OAI211_X1 _16490_ ( .A(_00480_ ), .B(_00492_ ), .C1(_07852_ ), .C2(_00490_ ), .ZN(_00493_ ) );
NOR3_X1 _16491_ ( .A1(_00485_ ), .A2(_07360_ ), .A3(_07808_ ), .ZN(_00494_ ) );
OAI21_X1 _16492_ ( .A(_07326_ ), .B1(_04653_ ), .B2(_07503_ ), .ZN(_00495_ ) );
NAND3_X1 _16493_ ( .A1(_07242_ ), .A2(_04058_ ), .A3(_07409_ ), .ZN(_00496_ ) );
OAI211_X1 _16494_ ( .A(_00495_ ), .B(_00496_ ), .C1(_07657_ ), .C2(_00485_ ), .ZN(_00497_ ) );
NOR3_X1 _16495_ ( .A1(_00493_ ), .A2(_00494_ ), .A3(_00497_ ), .ZN(_00498_ ) );
OAI221_X1 _16496_ ( .A(_04783_ ), .B1(_07531_ ), .B2(_00476_ ), .C1(_00498_ ), .C2(_07419_ ), .ZN(_00499_ ) );
NAND4_X1 _16497_ ( .A1(_05488_ ), .A2(_04920_ ), .A3(\ID_EX_typ [7] ), .A4(\ID_EX_typ [5] ), .ZN(_00500_ ) );
NAND3_X1 _16498_ ( .A1(_00499_ ), .A2(_07665_ ), .A3(_00500_ ), .ZN(_00501_ ) );
OR2_X1 _16499_ ( .A1(_07016_ ), .A2(_06700_ ), .ZN(_00502_ ) );
NAND2_X1 _16500_ ( .A1(_00501_ ), .A2(_00502_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
OR2_X1 _16501_ ( .A1(_07028_ ), .A2(_06700_ ), .ZN(_00503_ ) );
NAND2_X1 _16502_ ( .A1(_05183_ ), .A2(_07428_ ), .ZN(_00504_ ) );
NOR2_X1 _16503_ ( .A1(_08010_ ), .A2(_03870_ ), .ZN(_00505_ ) );
OR3_X1 _16504_ ( .A1(_00413_ ), .A2(_00505_ ), .A3(_07599_ ), .ZN(_00506_ ) );
NAND3_X1 _16505_ ( .A1(_07112_ ), .A2(\ID_EX_imm [28] ), .A3(_07109_ ), .ZN(_00507_ ) );
AND3_X1 _16506_ ( .A1(_00504_ ), .A2(_00506_ ), .A3(_00507_ ), .ZN(_00508_ ) );
AOI21_X1 _16507_ ( .A(_05495_ ), .B1(_00508_ ), .B2(_05672_ ), .ZN(_00509_ ) );
AND3_X1 _16508_ ( .A1(_07962_ ), .A2(_04531_ ), .A3(_07964_ ), .ZN(_00510_ ) );
OR3_X1 _16509_ ( .A1(_00510_ ), .A2(_07965_ ), .A3(_07809_ ), .ZN(_00511_ ) );
AOI21_X1 _16510_ ( .A(_07560_ ), .B1(_07931_ ), .B2(_07932_ ), .ZN(_00512_ ) );
OAI21_X1 _16511_ ( .A(_07286_ ), .B1(_07440_ ), .B2(_07438_ ), .ZN(_00513_ ) );
OAI21_X1 _16512_ ( .A(_07304_ ), .B1(_07437_ ), .B2(_07446_ ), .ZN(_00514_ ) );
AND3_X1 _16513_ ( .A1(_00513_ ), .A2(_00514_ ), .A3(_07650_ ), .ZN(_00515_ ) );
MUX2_X1 _16514_ ( .A(_07991_ ), .B(_07995_ ), .S(_07304_ ), .Z(_00516_ ) );
AOI211_X1 _16515_ ( .A(_07920_ ), .B(_00515_ ), .C1(_07697_ ), .C2(_00516_ ), .ZN(_00517_ ) );
AOI21_X1 _16516_ ( .A(_07638_ ), .B1(_07493_ ), .B2(_07500_ ), .ZN(_00518_ ) );
NOR3_X1 _16517_ ( .A1(_00517_ ), .A2(_07284_ ), .A3(_00518_ ), .ZN(_00519_ ) );
OAI21_X1 _16518_ ( .A(_07254_ ), .B1(_00512_ ), .B2(_00519_ ), .ZN(_00520_ ) );
NAND4_X1 _16519_ ( .A1(_07914_ ), .A2(_07434_ ), .A3(_07210_ ), .A4(_07725_ ), .ZN(_00521_ ) );
NAND2_X1 _16520_ ( .A1(_07917_ ), .A2(_07251_ ), .ZN(_00522_ ) );
NAND2_X1 _16521_ ( .A1(_00521_ ), .A2(_00522_ ), .ZN(_00523_ ) );
OAI21_X1 _16522_ ( .A(_07131_ ), .B1(_07984_ ), .B2(_00523_ ), .ZN(_00524_ ) );
NAND3_X1 _16523_ ( .A1(_07917_ ), .A2(_07560_ ), .A3(_07407_ ), .ZN(_00525_ ) );
OAI21_X1 _16524_ ( .A(_07329_ ), .B1(_03253_ ), .B2(_04529_ ), .ZN(_00526_ ) );
AOI22_X1 _16525_ ( .A1(_04530_ ), .A2(_07326_ ), .B1(_07967_ ), .B2(_04419_ ), .ZN(_00527_ ) );
AND4_X1 _16526_ ( .A1(_00524_ ), .A2(_00525_ ), .A3(_00526_ ), .A4(_00527_ ), .ZN(_00528_ ) );
NAND3_X1 _16527_ ( .A1(_00511_ ), .A2(_00520_ ), .A3(_00528_ ), .ZN(_00529_ ) );
AOI21_X1 _16528_ ( .A(_00509_ ), .B1(_00529_ ), .B2(_08125_ ), .ZN(_00530_ ) );
OAI21_X1 _16529_ ( .A(_08089_ ), .B1(_05182_ ), .B2(_05663_ ), .ZN(_00531_ ) );
OAI21_X1 _16530_ ( .A(_00503_ ), .B1(_00530_ ), .B2(_00531_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _16531_ ( .A1(_05466_ ), .A2(_05180_ ), .ZN(_00532_ ) );
NOR2_X1 _16532_ ( .A1(_04458_ ), .A2(_04481_ ), .ZN(_00533_ ) );
INV_X1 _16533_ ( .A(_03962_ ), .ZN(_00534_ ) );
NOR2_X1 _16534_ ( .A1(_00533_ ), .A2(_00534_ ), .ZN(_00535_ ) );
NOR3_X1 _16535_ ( .A1(_00535_ ), .A2(_04485_ ), .A3(_04484_ ), .ZN(_00536_ ) );
AOI21_X1 _16536_ ( .A(_00536_ ), .B1(_04488_ ), .B2(_03984_ ), .ZN(_00537_ ) );
AND2_X1 _16537_ ( .A1(_00537_ ), .A2(_04032_ ), .ZN(_00538_ ) );
OR3_X1 _16538_ ( .A1(_00538_ ), .A2(_04010_ ), .A3(_04492_ ), .ZN(_00539_ ) );
OAI21_X1 _16539_ ( .A(_04010_ ), .B1(_00538_ ), .B2(_04492_ ), .ZN(_00540_ ) );
AND3_X1 _16540_ ( .A1(_00539_ ), .A2(_07126_ ), .A3(_00540_ ), .ZN(_00541_ ) );
OAI22_X1 _16541_ ( .A1(_05470_ ), .A2(_07111_ ), .B1(_02484_ ), .B2(_07115_ ), .ZN(_00542_ ) );
OAI21_X1 _16542_ ( .A(_07417_ ), .B1(_00541_ ), .B2(_00542_ ), .ZN(_00543_ ) );
NAND2_X1 _16543_ ( .A1(_00543_ ), .A2(_04783_ ), .ZN(_00544_ ) );
AOI21_X1 _16544_ ( .A(_07945_ ), .B1(_07959_ ), .B2(_07960_ ), .ZN(_00545_ ) );
OR3_X1 _16545_ ( .A1(_00545_ ), .A2(_04717_ ), .A3(_04722_ ), .ZN(_00546_ ) );
OAI21_X1 _16546_ ( .A(_04717_ ), .B1(_00545_ ), .B2(_04722_ ), .ZN(_00547_ ) );
NAND3_X1 _16547_ ( .A1(_00546_ ), .A2(_07404_ ), .A3(_00547_ ), .ZN(_00548_ ) );
AND3_X1 _16548_ ( .A1(_07186_ ), .A2(_07543_ ), .A3(_07725_ ), .ZN(_00549_ ) );
AOI21_X1 _16549_ ( .A(_07322_ ), .B1(_07556_ ), .B2(_07557_ ), .ZN(_00550_ ) );
AND2_X1 _16550_ ( .A1(_00550_ ), .A2(_07249_ ), .ZN(_00551_ ) );
NOR2_X1 _16551_ ( .A1(_00549_ ), .A2(_00551_ ), .ZN(_00552_ ) );
AOI21_X1 _16552_ ( .A(_07804_ ), .B1(_07985_ ), .B2(_00552_ ), .ZN(_00553_ ) );
AND3_X1 _16553_ ( .A1(_00550_ ), .A2(_07461_ ), .A3(_07407_ ), .ZN(_00554_ ) );
OR2_X1 _16554_ ( .A1(_00553_ ), .A2(_00554_ ), .ZN(_00555_ ) );
OAI21_X1 _16555_ ( .A(_07292_ ), .B1(_07230_ ), .B2(_07235_ ), .ZN(_00556_ ) );
OAI21_X1 _16556_ ( .A(_07286_ ), .B1(_07287_ ), .B2(_07231_ ), .ZN(_00557_ ) );
NAND2_X1 _16557_ ( .A1(_00556_ ), .A2(_00557_ ), .ZN(_00558_ ) );
OAI21_X1 _16558_ ( .A(_07578_ ), .B1(_00558_ ), .B2(_07273_ ), .ZN(_00559_ ) );
OAI21_X1 _16559_ ( .A(_07292_ ), .B1(_07217_ ), .B2(_07223_ ), .ZN(_00560_ ) );
OAI21_X1 _16560_ ( .A(_07275_ ), .B1(_07236_ ), .B2(_07226_ ), .ZN(_00561_ ) );
AND3_X1 _16561_ ( .A1(_00560_ ), .A2(_07262_ ), .A3(_00561_ ), .ZN(_00562_ ) );
OAI21_X1 _16562_ ( .A(_07799_ ), .B1(_00559_ ), .B2(_00562_ ), .ZN(_00563_ ) );
AOI21_X1 _16563_ ( .A(_00563_ ), .B1(_07920_ ), .B2(_07585_ ), .ZN(_00564_ ) );
INV_X1 _16564_ ( .A(_07979_ ), .ZN(_00565_ ) );
AOI21_X1 _16565_ ( .A(_00565_ ), .B1(_08035_ ), .B2(_08036_ ), .ZN(_00566_ ) );
OR2_X1 _16566_ ( .A1(_00564_ ), .A2(_00566_ ), .ZN(_00567_ ) );
AND3_X1 _16567_ ( .A1(_04716_ ), .A2(_02483_ ), .A3(_02493_ ), .ZN(_00568_ ) );
NOR3_X1 _16568_ ( .A1(_07963_ ), .A2(_00568_ ), .A3(_07753_ ), .ZN(_00569_ ) );
OR3_X1 _16569_ ( .A1(_04490_ ), .A2(_04716_ ), .A3(_04420_ ), .ZN(_00570_ ) );
OAI21_X1 _16570_ ( .A(_00570_ ), .B1(_00568_ ), .B2(_07657_ ), .ZN(_00571_ ) );
NOR4_X1 _16571_ ( .A1(_00555_ ), .A2(_00567_ ), .A3(_00569_ ), .A4(_00571_ ), .ZN(_00572_ ) );
AOI21_X1 _16572_ ( .A(_07419_ ), .B1(_00548_ ), .B2(_00572_ ), .ZN(_00573_ ) );
OAI211_X1 _16573_ ( .A(_06994_ ), .B(_00532_ ), .C1(_00544_ ), .C2(_00573_ ), .ZN(_00574_ ) );
AND3_X1 _16574_ ( .A1(_05046_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_06446_ ), .ZN(_00575_ ) );
NAND4_X1 _16575_ ( .A1(_04896_ ), .A2(_04897_ ), .A3(\mycsreg.CSReg[3][27] ), .A4(_04992_ ), .ZN(_00576_ ) );
NAND4_X1 _16576_ ( .A1(_04987_ ), .A2(\mtvec [27] ), .A3(_04992_ ), .A4(_04993_ ), .ZN(_00577_ ) );
NAND4_X1 _16577_ ( .A1(_03552_ ), .A2(_05458_ ), .A3(_00576_ ), .A4(_00577_ ), .ZN(_00578_ ) );
AND4_X1 _16578_ ( .A1(\mycsreg.CSReg[0][27] ), .A2(_04991_ ), .A3(_04992_ ), .A4(_04993_ ), .ZN(_00579_ ) );
NOR2_X1 _16579_ ( .A1(_00578_ ), .A2(_00579_ ), .ZN(_00580_ ) );
AOI21_X1 _16580_ ( .A(_00580_ ), .B1(_05046_ ), .B2(_06446_ ), .ZN(_00581_ ) );
OAI21_X1 _16581_ ( .A(_06706_ ), .B1(_00575_ ), .B2(_00581_ ), .ZN(_00582_ ) );
NAND2_X1 _16582_ ( .A1(_00574_ ), .A2(_00582_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
NAND3_X1 _16583_ ( .A1(_07047_ ), .A2(_06706_ ), .A3(_07052_ ), .ZN(_00583_ ) );
NOR2_X1 _16584_ ( .A1(_00537_ ), .A2(_04032_ ), .ZN(_00584_ ) );
NOR3_X1 _16585_ ( .A1(_00538_ ), .A2(_00584_ ), .A3(_07600_ ), .ZN(_00585_ ) );
OAI22_X1 _16586_ ( .A1(_05500_ ), .A2(_07111_ ), .B1(_04719_ ), .B2(_07115_ ), .ZN(_00586_ ) );
OAI21_X1 _16587_ ( .A(_07417_ ), .B1(_00585_ ), .B2(_00586_ ), .ZN(_00587_ ) );
NAND2_X1 _16588_ ( .A1(_00587_ ), .A2(_04831_ ), .ZN(_00588_ ) );
AND3_X1 _16589_ ( .A1(_07959_ ), .A2(_07945_ ), .A3(_07960_ ), .ZN(_00589_ ) );
NOR3_X1 _16590_ ( .A1(_00589_ ), .A2(_00545_ ), .A3(_07809_ ), .ZN(_00590_ ) );
NAND3_X1 _16591_ ( .A1(_08077_ ), .A2(_07979_ ), .A3(_08078_ ), .ZN(_00591_ ) );
OR3_X1 _16592_ ( .A1(_04721_ ), .A2(_03227_ ), .A3(_07521_ ), .ZN(_00592_ ) );
AND3_X1 _16593_ ( .A1(_08000_ ), .A2(_07301_ ), .A3(_08001_ ), .ZN(_00593_ ) );
AOI21_X1 _16594_ ( .A(_00593_ ), .B1(_07697_ ), .B2(_07993_ ), .ZN(_00594_ ) );
MUX2_X1 _16595_ ( .A(_07646_ ), .B(_00594_ ), .S(_07696_ ), .Z(_00595_ ) );
OAI211_X1 _16596_ ( .A(_00591_ ), .B(_00592_ ), .C1(_00595_ ), .C2(_07930_ ), .ZN(_00596_ ) );
AND3_X1 _16597_ ( .A1(_07199_ ), .A2(_07610_ ), .A3(_07543_ ), .ZN(_00597_ ) );
NOR2_X1 _16598_ ( .A1(_07626_ ), .A2(_07322_ ), .ZN(_00598_ ) );
AOI22_X1 _16599_ ( .A1(_07607_ ), .A2(_00597_ ), .B1(_07250_ ), .B2(_00598_ ), .ZN(_00599_ ) );
AOI21_X1 _16600_ ( .A(_07804_ ), .B1(_07985_ ), .B2(_00599_ ), .ZN(_00600_ ) );
AND3_X1 _16601_ ( .A1(_00598_ ), .A2(_07250_ ), .A3(_07406_ ), .ZN(_00601_ ) );
NOR3_X1 _16602_ ( .A1(_04722_ ), .A2(_04723_ ), .A3(_07753_ ), .ZN(_00602_ ) );
AOI21_X1 _16603_ ( .A(_07523_ ), .B1(_04721_ ), .B2(_03227_ ), .ZN(_00603_ ) );
OR4_X1 _16604_ ( .A1(_00600_ ), .A2(_00601_ ), .A3(_00602_ ), .A4(_00603_ ), .ZN(_00604_ ) );
OR3_X1 _16605_ ( .A1(_00590_ ), .A2(_00596_ ), .A3(_00604_ ), .ZN(_00605_ ) );
AOI21_X1 _16606_ ( .A(_00588_ ), .B1(_00605_ ), .B2(_08125_ ), .ZN(_00606_ ) );
OAI21_X1 _16607_ ( .A(_08089_ ), .B1(_05502_ ), .B2(_04783_ ), .ZN(_00607_ ) );
OAI21_X1 _16608_ ( .A(_00583_ ), .B1(_00606_ ), .B2(_00607_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
NAND3_X1 _16609_ ( .A1(_05532_ ), .A2(_06706_ ), .A3(_05538_ ), .ZN(_00608_ ) );
OAI22_X1 _16610_ ( .A1(_05530_ ), .A2(_07111_ ), .B1(_03224_ ), .B2(_07115_ ), .ZN(_00609_ ) );
OR3_X1 _16611_ ( .A1(_00535_ ), .A2(_03985_ ), .A3(_04484_ ), .ZN(_00610_ ) );
OAI21_X1 _16612_ ( .A(_03985_ ), .B1(_00535_ ), .B2(_04484_ ), .ZN(_00611_ ) );
AND3_X1 _16613_ ( .A1(_00610_ ), .A2(_07125_ ), .A3(_00611_ ), .ZN(_00612_ ) );
OAI21_X1 _16614_ ( .A(_07417_ ), .B1(_00609_ ), .B2(_00612_ ), .ZN(_00613_ ) );
NAND2_X1 _16615_ ( .A1(_00613_ ), .A2(_04831_ ), .ZN(_00614_ ) );
AOI21_X1 _16616_ ( .A(_00565_ ), .B1(_08113_ ), .B2(_08114_ ), .ZN(_00615_ ) );
NOR3_X1 _16617_ ( .A1(_07684_ ), .A2(_07688_ ), .A3(_07323_ ), .ZN(_00616_ ) );
NAND2_X1 _16618_ ( .A1(_00616_ ), .A2(_07407_ ), .ZN(_00617_ ) );
NOR4_X1 _16619_ ( .A1(_08098_ ), .A2(_07188_ ), .A3(_07212_ ), .A4(_07138_ ), .ZN(_00618_ ) );
NOR3_X1 _16620_ ( .A1(_07984_ ), .A2(_00618_ ), .A3(_00616_ ), .ZN(_00619_ ) );
OAI21_X1 _16621_ ( .A(_00617_ ), .B1(_00619_ ), .B2(_07805_ ), .ZN(_00620_ ) );
OR3_X1 _16622_ ( .A1(_07288_ ), .A2(_07293_ ), .A3(_07916_ ), .ZN(_00621_ ) );
NAND3_X1 _16623_ ( .A1(_00433_ ), .A2(_00434_ ), .A3(_07697_ ), .ZN(_00622_ ) );
NAND3_X1 _16624_ ( .A1(_00621_ ), .A2(_07638_ ), .A3(_00622_ ), .ZN(_00623_ ) );
OAI21_X1 _16625_ ( .A(_00623_ ), .B1(_07638_ ), .B2(_07694_ ), .ZN(_00624_ ) );
AOI211_X1 _16626_ ( .A(_00615_ ), .B(_00620_ ), .C1(_07799_ ), .C2(_00624_ ), .ZN(_00625_ ) );
OR2_X1 _16627_ ( .A1(_07957_ ), .A2(_04732_ ), .ZN(_00626_ ) );
INV_X1 _16628_ ( .A(_04729_ ), .ZN(_00627_ ) );
AND3_X1 _16629_ ( .A1(_00626_ ), .A2(_00627_ ), .A3(_04739_ ), .ZN(_00628_ ) );
AOI21_X1 _16630_ ( .A(_04739_ ), .B1(_00626_ ), .B2(_00627_ ), .ZN(_00629_ ) );
OR3_X1 _16631_ ( .A1(_00628_ ), .A2(_00629_ ), .A3(_07809_ ), .ZN(_00630_ ) );
NOR3_X1 _16632_ ( .A1(_04736_ ), .A2(_04737_ ), .A3(_07753_ ), .ZN(_00631_ ) );
AOI21_X1 _16633_ ( .A(_07657_ ), .B1(_04735_ ), .B2(_04488_ ), .ZN(_00632_ ) );
NOR3_X1 _16634_ ( .A1(_04735_ ), .A2(_04488_ ), .A3(_07521_ ), .ZN(_00633_ ) );
NOR3_X1 _16635_ ( .A1(_00631_ ), .A2(_00632_ ), .A3(_00633_ ), .ZN(_00634_ ) );
NAND3_X1 _16636_ ( .A1(_00625_ ), .A2(_00630_ ), .A3(_00634_ ), .ZN(_00635_ ) );
AOI21_X1 _16637_ ( .A(_00614_ ), .B1(_00635_ ), .B2(_08125_ ), .ZN(_00636_ ) );
OAI21_X1 _16638_ ( .A(_08089_ ), .B1(_05525_ ), .B2(_04783_ ), .ZN(_00637_ ) );
OAI21_X1 _16639_ ( .A(_00608_ ), .B1(_00636_ ), .B2(_00637_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
OR2_X1 _16640_ ( .A1(_07071_ ), .A2(_06694_ ), .ZN(_00638_ ) );
NAND2_X1 _16641_ ( .A1(_05557_ ), .A2(_07428_ ), .ZN(_00639_ ) );
OAI21_X1 _16642_ ( .A(_00639_ ), .B1(_03173_ ), .B2(_07115_ ), .ZN(_00640_ ) );
OAI21_X1 _16643_ ( .A(_07125_ ), .B1(_00533_ ), .B2(_00534_ ), .ZN(_00641_ ) );
AOI21_X1 _16644_ ( .A(_00641_ ), .B1(_00534_ ), .B2(_00533_ ), .ZN(_00642_ ) );
OAI21_X1 _16645_ ( .A(_07417_ ), .B1(_00640_ ), .B2(_00642_ ), .ZN(_00643_ ) );
NAND2_X1 _16646_ ( .A1(_00643_ ), .A2(_04831_ ), .ZN(_00644_ ) );
AOI21_X1 _16647_ ( .A(_07809_ ), .B1(_07958_ ), .B2(_04731_ ), .ZN(_00645_ ) );
OAI21_X1 _16648_ ( .A(_00645_ ), .B1(_04731_ ), .B2(_07958_ ), .ZN(_00646_ ) );
OAI211_X1 _16649_ ( .A(_07914_ ), .B(_07725_ ), .C1(_07802_ ), .C2(_08137_ ), .ZN(_00647_ ) );
INV_X1 _16650_ ( .A(_00647_ ), .ZN(_00648_ ) );
NOR3_X1 _16651_ ( .A1(_07734_ ), .A2(_07284_ ), .A3(_07920_ ), .ZN(_00649_ ) );
OAI21_X1 _16652_ ( .A(_07131_ ), .B1(_00648_ ), .B2(_00649_ ), .ZN(_00650_ ) );
NAND2_X1 _16653_ ( .A1(_00649_ ), .A2(_07408_ ), .ZN(_00651_ ) );
NAND3_X1 _16654_ ( .A1(_08155_ ), .A2(_07979_ ), .A3(_08156_ ), .ZN(_00652_ ) );
NAND2_X1 _16655_ ( .A1(_00651_ ), .A2(_00652_ ), .ZN(_00653_ ) );
NOR3_X1 _16656_ ( .A1(_04728_ ), .A2(_04483_ ), .A3(_07521_ ), .ZN(_00654_ ) );
OAI22_X1 _16657_ ( .A1(_04732_ ), .A2(_07753_ ), .B1(_04730_ ), .B2(_07524_ ), .ZN(_00655_ ) );
OR3_X1 _16658_ ( .A1(_07741_ ), .A2(_07742_ ), .A3(_07630_ ), .ZN(_00656_ ) );
NAND3_X1 _16659_ ( .A1(_00513_ ), .A2(_00514_ ), .A3(_07916_ ), .ZN(_00657_ ) );
OAI211_X1 _16660_ ( .A(_00657_ ), .B(_07696_ ), .C1(_07499_ ), .C2(_07697_ ), .ZN(_00658_ ) );
AND3_X1 _16661_ ( .A1(_00656_ ), .A2(_07799_ ), .A3(_00658_ ), .ZN(_00659_ ) );
NOR4_X1 _16662_ ( .A1(_00653_ ), .A2(_00654_ ), .A3(_00655_ ), .A4(_00659_ ), .ZN(_00660_ ) );
NAND3_X1 _16663_ ( .A1(_00646_ ), .A2(_00650_ ), .A3(_00660_ ), .ZN(_00661_ ) );
AOI21_X1 _16664_ ( .A(_00644_ ), .B1(_00661_ ), .B2(_08125_ ), .ZN(_00662_ ) );
OAI21_X1 _16665_ ( .A(_08089_ ), .B1(_05556_ ), .B2(_04783_ ), .ZN(_00663_ ) );
OAI21_X1 _16666_ ( .A(_00638_ ), .B1(_00662_ ), .B2(_00663_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
NAND3_X1 _16667_ ( .A1(_05577_ ), .A2(_06706_ ), .A3(_05584_ ), .ZN(_00664_ ) );
OAI21_X1 _16668_ ( .A(_04472_ ), .B1(_07121_ ), .B2(_03793_ ), .ZN(_00665_ ) );
AOI21_X1 _16669_ ( .A(_04478_ ), .B1(_00665_ ), .B2(_03839_ ), .ZN(_00666_ ) );
XNOR2_X1 _16670_ ( .A(_00666_ ), .B(_03817_ ), .ZN(_00667_ ) );
NAND2_X1 _16671_ ( .A1(_00667_ ), .A2(_07126_ ), .ZN(_00668_ ) );
AOI22_X1 _16672_ ( .A1(_05575_ ), .A2(_07110_ ), .B1(\ID_EX_imm [23] ), .B2(_07114_ ), .ZN(_00669_ ) );
AOI21_X1 _16673_ ( .A(_07418_ ), .B1(_00668_ ), .B2(_00669_ ), .ZN(_00670_ ) );
OR2_X1 _16674_ ( .A1(_00670_ ), .A2(_07662_ ), .ZN(_00671_ ) );
OAI21_X1 _16675_ ( .A(_07946_ ), .B1(_07386_ ), .B2(_07394_ ), .ZN(_00672_ ) );
AOI21_X1 _16676_ ( .A(_07950_ ), .B1(_00672_ ), .B2(_07949_ ), .ZN(_00673_ ) );
OR3_X1 _16677_ ( .A1(_00673_ ), .A2(_04540_ ), .A3(_07954_ ), .ZN(_00674_ ) );
OAI21_X1 _16678_ ( .A(_04540_ ), .B1(_00673_ ), .B2(_07954_ ), .ZN(_00675_ ) );
NAND3_X1 _16679_ ( .A1(_00674_ ), .A2(_07404_ ), .A3(_00675_ ), .ZN(_00676_ ) );
NAND3_X1 _16680_ ( .A1(_08178_ ), .A2(_07560_ ), .A3(_07408_ ), .ZN(_00677_ ) );
OAI21_X1 _16681_ ( .A(_07329_ ), .B1(_07149_ ), .B2(_02548_ ), .ZN(_00678_ ) );
AND2_X1 _16682_ ( .A1(_00677_ ), .A2(_00678_ ), .ZN(_00679_ ) );
OAI21_X1 _16683_ ( .A(_07914_ ), .B1(_07802_ ), .B2(_07544_ ), .ZN(_00680_ ) );
NOR2_X1 _16684_ ( .A1(_00680_ ), .A2(_07138_ ), .ZN(_00681_ ) );
AND2_X1 _16685_ ( .A1(_08178_ ), .A2(_07464_ ), .ZN(_00682_ ) );
OAI21_X1 _16686_ ( .A(_07130_ ), .B1(_00681_ ), .B2(_00682_ ), .ZN(_00683_ ) );
NOR3_X1 _16687_ ( .A1(_07793_ ), .A2(_07464_ ), .A3(_07920_ ), .ZN(_00684_ ) );
OR3_X1 _16688_ ( .A1(_07579_ ), .A2(_07580_ ), .A3(_07433_ ), .ZN(_00685_ ) );
NAND2_X1 _16689_ ( .A1(_00558_ ), .A2(_07916_ ), .ZN(_00686_ ) );
AOI21_X1 _16690_ ( .A(_07323_ ), .B1(_00685_ ), .B2(_00686_ ), .ZN(_00687_ ) );
AND3_X1 _16691_ ( .A1(_07795_ ), .A2(_07514_ ), .A3(_07796_ ), .ZN(_00688_ ) );
NOR3_X1 _16692_ ( .A1(_00687_ ), .A2(_00688_ ), .A3(_07284_ ), .ZN(_00689_ ) );
OAI21_X1 _16693_ ( .A(_07254_ ), .B1(_00684_ ), .B2(_00689_ ), .ZN(_00690_ ) );
NAND2_X1 _16694_ ( .A1(_04540_ ), .A2(_07327_ ), .ZN(_00691_ ) );
NAND3_X1 _16695_ ( .A1(_07149_ ), .A2(_02548_ ), .A3(_07409_ ), .ZN(_00692_ ) );
AND4_X1 _16696_ ( .A1(_00683_ ), .A2(_00690_ ), .A3(_00691_ ), .A4(_00692_ ), .ZN(_00693_ ) );
NAND3_X1 _16697_ ( .A1(_00676_ ), .A2(_00679_ ), .A3(_00693_ ), .ZN(_00694_ ) );
AOI21_X1 _16698_ ( .A(_00671_ ), .B1(_00694_ ), .B2(_07420_ ), .ZN(_00695_ ) );
OAI21_X1 _16699_ ( .A(_08089_ ), .B1(_05569_ ), .B2(_04783_ ), .ZN(_00696_ ) );
OAI21_X1 _16700_ ( .A(_00664_ ), .B1(_00695_ ), .B2(_00696_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
OAI211_X1 _16701_ ( .A(_06802_ ), .B(_07082_ ), .C1(_07083_ ), .C2(_07087_ ), .ZN(_00697_ ) );
OAI22_X1 _16702_ ( .A1(_05607_ ), .A2(_07111_ ), .B1(_02523_ ), .B2(_07115_ ), .ZN(_00698_ ) );
OR2_X1 _16703_ ( .A1(_00665_ ), .A2(_03839_ ), .ZN(_00699_ ) );
AOI21_X1 _16704_ ( .A(_07600_ ), .B1(_00665_ ), .B2(_03839_ ), .ZN(_00700_ ) );
AOI21_X1 _16705_ ( .A(_00698_ ), .B1(_00699_ ), .B2(_00700_ ), .ZN(_00701_ ) );
AOI21_X1 _16706_ ( .A(_05495_ ), .B1(_00701_ ), .B2(_05672_ ), .ZN(_00702_ ) );
NAND3_X1 _16707_ ( .A1(_07200_ ), .A2(_07212_ ), .A3(_07828_ ), .ZN(_00703_ ) );
AOI211_X1 _16708_ ( .A(_07138_ ), .B(_07188_ ), .C1(_07187_ ), .C2(_00703_ ), .ZN(_00704_ ) );
AND2_X1 _16709_ ( .A1(_08212_ ), .A2(_07251_ ), .ZN(_00705_ ) );
OAI21_X1 _16710_ ( .A(_07130_ ), .B1(_00704_ ), .B2(_00705_ ), .ZN(_00706_ ) );
NAND3_X1 _16711_ ( .A1(_08212_ ), .A2(_07560_ ), .A3(_07407_ ), .ZN(_00707_ ) );
NAND3_X1 _16712_ ( .A1(_07150_ ), .A2(_02522_ ), .A3(_07409_ ), .ZN(_00708_ ) );
AOI21_X1 _16713_ ( .A(_07524_ ), .B1(_04535_ ), .B2(_07953_ ), .ZN(_00709_ ) );
AOI21_X1 _16714_ ( .A(_00709_ ), .B1(_04536_ ), .B2(_07326_ ), .ZN(_00710_ ) );
NAND4_X1 _16715_ ( .A1(_00706_ ), .A2(_00707_ ), .A3(_00708_ ), .A4(_00710_ ), .ZN(_00711_ ) );
AND3_X1 _16716_ ( .A1(_00672_ ), .A2(_07950_ ), .A3(_07949_ ), .ZN(_00712_ ) );
NOR3_X1 _16717_ ( .A1(_00712_ ), .A2(_00673_ ), .A3(_07808_ ), .ZN(_00713_ ) );
NOR2_X1 _16718_ ( .A1(_07845_ ), .A2(_07920_ ), .ZN(_00714_ ) );
OAI21_X1 _16719_ ( .A(_07254_ ), .B1(_00714_ ), .B2(_07464_ ), .ZN(_00715_ ) );
AND2_X1 _16720_ ( .A1(_07847_ ), .A2(_07848_ ), .ZN(_00716_ ) );
MUX2_X1 _16721_ ( .A(_08004_ ), .B(_00716_ ), .S(_07280_ ), .Z(_00717_ ) );
AOI21_X1 _16722_ ( .A(_00715_ ), .B1(_07560_ ), .B2(_00717_ ), .ZN(_00718_ ) );
OR3_X1 _16723_ ( .A1(_00711_ ), .A2(_00713_ ), .A3(_00718_ ), .ZN(_00719_ ) );
AOI21_X1 _16724_ ( .A(_00702_ ), .B1(_00719_ ), .B2(_07420_ ), .ZN(_00720_ ) );
NAND2_X1 _16725_ ( .A1(_05604_ ), .A2(_07663_ ), .ZN(_00721_ ) );
NAND2_X1 _16726_ ( .A1(_00721_ ), .A2(_07665_ ), .ZN(_00722_ ) );
OAI21_X1 _16727_ ( .A(_00697_ ), .B1(_00720_ ), .B2(_00722_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NAND3_X1 _16728_ ( .A1(_07095_ ), .A2(_06706_ ), .A3(_07100_ ), .ZN(_00723_ ) );
NAND2_X1 _16729_ ( .A1(_05646_ ), .A2(_07428_ ), .ZN(_00724_ ) );
NOR2_X1 _16730_ ( .A1(_08011_ ), .A2(_08012_ ), .ZN(_00725_ ) );
OR3_X1 _16731_ ( .A1(_00725_ ), .A2(_03917_ ), .A3(_04503_ ), .ZN(_00726_ ) );
OAI21_X1 _16732_ ( .A(_03917_ ), .B1(_00725_ ), .B2(_04503_ ), .ZN(_00727_ ) );
NAND3_X1 _16733_ ( .A1(_00726_ ), .A2(_07125_ ), .A3(_00727_ ), .ZN(_00728_ ) );
NAND3_X1 _16734_ ( .A1(_07112_ ), .A2(\ID_EX_imm [31] ), .A3(_07109_ ), .ZN(_00729_ ) );
AND3_X1 _16735_ ( .A1(_00724_ ), .A2(_00728_ ), .A3(_00729_ ), .ZN(_00730_ ) );
AOI21_X1 _16736_ ( .A(_05495_ ), .B1(_00730_ ), .B2(_05672_ ), .ZN(_00731_ ) );
NOR2_X1 _16737_ ( .A1(_07154_ ), .A2(_03310_ ), .ZN(_00732_ ) );
OR3_X4 _16738_ ( .A1(_07971_ ), .A2(_04521_ ), .A3(_00732_ ), .ZN(_00733_ ) );
OAI21_X1 _16739_ ( .A(_04521_ ), .B1(_07971_ ), .B2(_00732_ ), .ZN(_00734_ ) );
AND3_X2 _16740_ ( .A1(_00733_ ), .A2(_07403_ ), .A3(_00734_ ), .ZN(_00735_ ) );
OAI211_X1 _16741_ ( .A(_07241_ ), .B(_07304_ ), .C1(_03310_ ), .C2(_07204_ ), .ZN(_00736_ ) );
OAI21_X1 _16742_ ( .A(_07286_ ), .B1(_07218_ ), .B2(_07244_ ), .ZN(_00737_ ) );
AND3_X1 _16743_ ( .A1(_00736_ ), .A2(_07697_ ), .A3(_00737_ ), .ZN(_00738_ ) );
AND3_X1 _16744_ ( .A1(_00560_ ), .A2(_07650_ ), .A3(_00561_ ), .ZN(_00739_ ) );
OAI21_X1 _16745_ ( .A(_07638_ ), .B1(_00738_ ), .B2(_00739_ ), .ZN(_00740_ ) );
NAND3_X1 _16746_ ( .A1(_00685_ ), .A2(_07920_ ), .A3(_00686_ ), .ZN(_00741_ ) );
AOI21_X1 _16747_ ( .A(_07930_ ), .B1(_00740_ ), .B2(_00741_ ), .ZN(_00742_ ) );
AOI22_X1 _16748_ ( .A1(_07186_ ), .A2(_07725_ ), .B1(_03337_ ), .B2(_07136_ ), .ZN(_00743_ ) );
NOR2_X1 _16749_ ( .A1(_00743_ ), .A2(_07804_ ), .ZN(_00744_ ) );
AND3_X1 _16750_ ( .A1(_07794_ ), .A2(_07797_ ), .A3(_07979_ ), .ZN(_00745_ ) );
AND3_X1 _16751_ ( .A1(_04758_ ), .A2(_03337_ ), .A3(_04419_ ), .ZN(_00746_ ) );
OR3_X1 _16752_ ( .A1(_07789_ ), .A2(_04630_ ), .A3(_07852_ ), .ZN(_00747_ ) );
OAI21_X1 _16753_ ( .A(_07329_ ), .B1(_04758_ ), .B2(_03337_ ), .ZN(_00748_ ) );
OAI211_X1 _16754_ ( .A(_00747_ ), .B(_00748_ ), .C1(_04520_ ), .C2(_07753_ ), .ZN(_00749_ ) );
OR4_X1 _16755_ ( .A1(_00744_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_00749_ ), .ZN(_00750_ ) );
OR3_X2 _16756_ ( .A1(_00735_ ), .A2(_00742_ ), .A3(_00750_ ), .ZN(_00751_ ) );
AOI21_X1 _16757_ ( .A(_00731_ ), .B1(_00751_ ), .B2(_07420_ ), .ZN(_00752_ ) );
OAI21_X1 _16758_ ( .A(_08089_ ), .B1(_05659_ ), .B2(_04783_ ), .ZN(_00753_ ) );
OAI21_X1 _16759_ ( .A(_00723_ ), .B1(_00752_ ), .B2(_00753_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
AOI21_X1 _16760_ ( .A(_02389_ ), .B1(_02355_ ), .B2(_02402_ ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _16761_ ( .A1(_05983_ ), .A2(IDU_valid_EXU ), .ZN(_00754_ ) );
OAI21_X1 _16762_ ( .A(_00754_ ), .B1(_05854_ ), .B2(_05870_ ), .ZN(_00755_ ) );
NAND2_X1 _16763_ ( .A1(_05920_ ), .A2(_00754_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
AND2_X1 _16764_ ( .A1(_00755_ ), .A2(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16765_ ( .A1(_05871_ ), .A2(_05920_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16766_ ( .A1(_05871_ ), .A2(_05920_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND4_X1 _16767_ ( .A1(_06257_ ), .A2(_06426_ ), .A3(_05759_ ), .A4(_05917_ ), .ZN(_00756_ ) );
NOR2_X1 _16768_ ( .A1(_05871_ ), .A2(_00756_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16769_ ( .A1(_06252_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_05718_ ), .A4(_05918_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16770_ ( .A(_06426_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16771_ ( .A1(_05919_ ), .A2(_05983_ ), .B1(_02272_ ), .B2(_02405_ ), .ZN(_00757_ ) );
INV_X1 _16772_ ( .A(loaduse_clear ), .ZN(_00758_ ) );
AOI221_X4 _16773_ ( .A(_00757_ ), .B1(\myidu.state [2] ), .B2(_00758_ ), .C1(_05871_ ), .C2(_06426_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16774_ ( .A(_05970_ ), .ZN(_00759_ ) );
OAI21_X1 _16775_ ( .A(_05966_ ), .B1(_00759_ ), .B2(_05709_ ), .ZN(_00760_ ) );
AND3_X1 _16776_ ( .A1(_05919_ ), .A2(IDU_ready_IFU ), .A3(_05703_ ), .ZN(_00761_ ) );
NOR3_X1 _16777_ ( .A1(_05836_ ), .A2(_05824_ ), .A3(_05840_ ), .ZN(_00762_ ) );
NAND4_X1 _16778_ ( .A1(_00762_ ), .A2(_05796_ ), .A3(_05985_ ), .A4(_05987_ ), .ZN(_00763_ ) );
OAI21_X1 _16779_ ( .A(_05980_ ), .B1(_05870_ ), .B2(_00763_ ), .ZN(_00764_ ) );
NAND3_X1 _16780_ ( .A1(_00760_ ), .A2(_00761_ ), .A3(_00764_ ), .ZN(_00765_ ) );
OR3_X1 _16781_ ( .A1(_05704_ ), .A2(_02405_ ), .A3(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_00766_ ) );
NAND3_X1 _16782_ ( .A1(_05759_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_00767_ ) );
NAND3_X1 _16783_ ( .A1(_00765_ ), .A2(_00766_ ), .A3(_00767_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16784_ ( .A(_04868_ ), .B(_05759_ ), .C1(_05919_ ), .C2(_05983_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
NAND2_X1 _16785_ ( .A1(_00760_ ), .A2(_00764_ ), .ZN(_00768_ ) );
NAND2_X1 _16786_ ( .A1(_00768_ ), .A2(_00761_ ), .ZN(_00769_ ) );
NAND3_X1 _16787_ ( .A1(_05759_ ), .A2(\myidu.state [2] ), .A3(_00758_ ), .ZN(_00770_ ) );
NAND2_X1 _16788_ ( .A1(_00769_ ), .A2(_00770_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16789_ ( .A1(_05916_ ), .A2(IDU_ready_IFU ), .ZN(_00771_ ) );
OAI21_X1 _16790_ ( .A(_01886_ ), .B1(_05916_ ), .B2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00772_ ) );
INV_X1 _16791_ ( .A(\myifu.state [0] ), .ZN(_00773_ ) );
AOI211_X1 _16792_ ( .A(_00771_ ), .B(_00772_ ), .C1(_00773_ ), .C2(_05916_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
OR3_X1 _16793_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06547_ ), .ZN(_00774_ ) );
OAI21_X1 _16794_ ( .A(_00774_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06548_ ), .ZN(_00775_ ) );
MUX2_X1 _16795_ ( .A(\io_master_rdata [31] ), .B(_00775_ ), .S(_02317_ ), .Z(_00776_ ) );
AND2_X1 _16796_ ( .A1(_00776_ ), .A2(_06527_ ), .ZN(\myifu.data_in [31] ) );
CLKBUF_X2 _16797_ ( .A(_02319_ ), .Z(_00777_ ) );
CLKBUF_X2 _16798_ ( .A(_06547_ ), .Z(_00778_ ) );
OR3_X1 _16799_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00779_ ) );
OAI211_X1 _16800_ ( .A(_02368_ ), .B(_00779_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00780_ ) );
BUF_X2 _16801_ ( .A(_02367_ ), .Z(_00781_ ) );
BUF_X4 _16802_ ( .A(_00781_ ), .Z(_00782_ ) );
OAI21_X1 _16803_ ( .A(_00780_ ), .B1(\io_master_rdata [30] ), .B2(_00782_ ), .ZN(_00783_ ) );
BUF_X4 _16804_ ( .A(_06516_ ), .Z(_00784_ ) );
NOR2_X1 _16805_ ( .A1(_00783_ ), .A2(_00784_ ), .ZN(\myifu.data_in [30] ) );
OR2_X1 _16806_ ( .A1(_00781_ ), .A2(\io_master_rdata [21] ), .ZN(_00785_ ) );
BUF_X2 _16807_ ( .A(_02367_ ), .Z(_00786_ ) );
OR3_X1 _16808_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00787_ ) );
OAI211_X1 _16809_ ( .A(_00786_ ), .B(_00787_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00788_ ) );
AND3_X1 _16810_ ( .A1(_00785_ ), .A2(_00788_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [21] ) );
OR2_X1 _16811_ ( .A1(_00781_ ), .A2(\io_master_rdata [20] ), .ZN(_00789_ ) );
OR3_X1 _16812_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00790_ ) );
OAI211_X1 _16813_ ( .A(_00786_ ), .B(_00790_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00791_ ) );
AND3_X1 _16814_ ( .A1(_00789_ ), .A2(_00791_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [20] ) );
OR2_X1 _16815_ ( .A1(_00781_ ), .A2(\io_master_rdata [19] ), .ZN(_00792_ ) );
OR3_X1 _16816_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00793_ ) );
OAI211_X1 _16817_ ( .A(_00786_ ), .B(_00793_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00794_ ) );
AND3_X1 _16818_ ( .A1(_00792_ ), .A2(_00794_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [19] ) );
OR2_X1 _16819_ ( .A1(_00781_ ), .A2(\io_master_rdata [18] ), .ZN(_00795_ ) );
OR3_X1 _16820_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00796_ ) );
OAI211_X1 _16821_ ( .A(_00786_ ), .B(_00796_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00797_ ) );
AND3_X1 _16822_ ( .A1(_00795_ ), .A2(_00797_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [18] ) );
OR2_X1 _16823_ ( .A1(_00781_ ), .A2(\io_master_rdata [17] ), .ZN(_00798_ ) );
OR3_X1 _16824_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00799_ ) );
OAI211_X1 _16825_ ( .A(_00786_ ), .B(_00799_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00800_ ) );
AND3_X1 _16826_ ( .A1(_00798_ ), .A2(_00800_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [17] ) );
OR2_X1 _16827_ ( .A1(_00781_ ), .A2(\io_master_rdata [16] ), .ZN(_00801_ ) );
OR3_X1 _16828_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00802_ ) );
OAI211_X1 _16829_ ( .A(_00781_ ), .B(_00802_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00803_ ) );
CLKBUF_X2 _16830_ ( .A(_06527_ ), .Z(_00804_ ) );
AND3_X1 _16831_ ( .A1(_00801_ ), .A2(_00803_ ), .A3(_00804_ ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16832_ ( .A1(_02251_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06547_ ), .ZN(_00805_ ) );
OAI211_X1 _16833_ ( .A(_02367_ ), .B(_00805_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06548_ ), .ZN(_00806_ ) );
OAI21_X2 _16834_ ( .A(_00806_ ), .B1(\io_master_rdata [15] ), .B2(_02367_ ), .ZN(_00807_ ) );
NOR2_X1 _16835_ ( .A1(_00807_ ), .A2(_00784_ ), .ZN(\myifu.data_in [15] ) );
OR2_X1 _16836_ ( .A1(_02368_ ), .A2(\io_master_rdata [14] ), .ZN(_00808_ ) );
CLKBUF_X2 _16837_ ( .A(_00778_ ), .Z(_00809_ ) );
OR3_X1 _16838_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00810_ ) );
OAI211_X1 _16839_ ( .A(_00782_ ), .B(_00810_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00811_ ) );
AND3_X1 _16840_ ( .A1(_00808_ ), .A2(_00811_ ), .A3(_00804_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16841_ ( .A1(_02368_ ), .A2(\io_master_rdata [13] ), .ZN(_00812_ ) );
CLKBUF_X2 _16842_ ( .A(_00778_ ), .Z(_00813_ ) );
OR3_X1 _16843_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00814_ ) );
BUF_X4 _16844_ ( .A(_06548_ ), .Z(_00815_ ) );
OAI211_X1 _16845_ ( .A(_00782_ ), .B(_00814_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00816_ ) );
AND3_X1 _16846_ ( .A1(_00812_ ), .A2(_00816_ ), .A3(_00804_ ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _16847_ ( .A1(_02368_ ), .A2(\io_master_rdata [12] ), .ZN(_00817_ ) );
OR3_X1 _16848_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00818_ ) );
OAI211_X1 _16849_ ( .A(_00782_ ), .B(_00818_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00819_ ) );
AND3_X1 _16850_ ( .A1(_00817_ ), .A2(_00819_ ), .A3(_00804_ ), .ZN(\myifu.data_in [12] ) );
OR2_X1 _16851_ ( .A1(_00786_ ), .A2(\io_master_rdata [29] ), .ZN(_00820_ ) );
OR3_X1 _16852_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00821_ ) );
OAI211_X1 _16853_ ( .A(_02368_ ), .B(_00821_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00822_ ) );
AND3_X1 _16854_ ( .A1(_00820_ ), .A2(_00822_ ), .A3(_00804_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16855_ ( .A1(_02369_ ), .A2(\io_master_rdata [11] ), .ZN(_00823_ ) );
OR3_X1 _16856_ ( .A1(_02321_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00824_ ) );
OAI211_X1 _16857_ ( .A(_02369_ ), .B(_00824_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00825_ ) );
AND3_X1 _16858_ ( .A1(_00823_ ), .A2(_00825_ ), .A3(_00804_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16859_ ( .A1(_02369_ ), .A2(\io_master_rdata [10] ), .ZN(_00826_ ) );
OR3_X1 _16860_ ( .A1(_02321_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00827_ ) );
OAI211_X1 _16861_ ( .A(_02369_ ), .B(_00827_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00828_ ) );
AND3_X1 _16862_ ( .A1(_00826_ ), .A2(_00828_ ), .A3(_00804_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16863_ ( .A1(_02369_ ), .A2(\io_master_rdata [9] ), .ZN(_00829_ ) );
OR3_X1 _16864_ ( .A1(_02321_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00830_ ) );
OAI211_X1 _16865_ ( .A(_02369_ ), .B(_00830_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00831_ ) );
AND3_X1 _16866_ ( .A1(_00829_ ), .A2(_00831_ ), .A3(_00804_ ), .ZN(\myifu.data_in [9] ) );
BUF_X2 _16867_ ( .A(_00781_ ), .Z(_00832_ ) );
OR2_X1 _16868_ ( .A1(_00832_ ), .A2(\io_master_rdata [8] ), .ZN(_00833_ ) );
OR3_X1 _16869_ ( .A1(_02321_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00834_ ) );
OAI211_X1 _16870_ ( .A(_02369_ ), .B(_00834_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00835_ ) );
AND3_X1 _16871_ ( .A1(_00833_ ), .A2(_00835_ ), .A3(_00804_ ), .ZN(\myifu.data_in [8] ) );
OR3_X1 _16872_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06547_ ), .ZN(_00836_ ) );
OAI211_X1 _16873_ ( .A(_02367_ ), .B(_00836_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06548_ ), .ZN(_00837_ ) );
OAI21_X1 _16874_ ( .A(_00837_ ), .B1(\io_master_rdata [7] ), .B2(_02367_ ), .ZN(_00838_ ) );
NOR2_X1 _16875_ ( .A1(_00838_ ), .A2(_00784_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16876_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00839_ ) );
OAI211_X1 _16877_ ( .A(_00782_ ), .B(_00839_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00840_ ) );
OAI21_X1 _16878_ ( .A(_00840_ ), .B1(\io_master_rdata [6] ), .B2(_00832_ ), .ZN(_00841_ ) );
NOR2_X1 _16879_ ( .A1(_00841_ ), .A2(_00784_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16880_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00842_ ) );
OAI211_X1 _16881_ ( .A(_00782_ ), .B(_00842_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00843_ ) );
OAI21_X1 _16882_ ( .A(_00843_ ), .B1(\io_master_rdata [5] ), .B2(_00832_ ), .ZN(_00844_ ) );
NOR2_X1 _16883_ ( .A1(_00844_ ), .A2(_00784_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16884_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00845_ ) );
OAI211_X1 _16885_ ( .A(_00782_ ), .B(_00845_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00846_ ) );
OAI21_X1 _16886_ ( .A(_00846_ ), .B1(\io_master_rdata [4] ), .B2(_00832_ ), .ZN(_00847_ ) );
NOR2_X1 _16887_ ( .A1(_00847_ ), .A2(_00784_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16888_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00848_ ) );
OAI211_X1 _16889_ ( .A(_00782_ ), .B(_00848_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00849_ ) );
OAI21_X1 _16890_ ( .A(_00849_ ), .B1(\io_master_rdata [3] ), .B2(_00832_ ), .ZN(_00850_ ) );
NOR2_X1 _16891_ ( .A1(_00850_ ), .A2(_00784_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16892_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00851_ ) );
OAI211_X1 _16893_ ( .A(_00782_ ), .B(_00851_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00852_ ) );
OAI21_X1 _16894_ ( .A(_00852_ ), .B1(\io_master_rdata [2] ), .B2(_00832_ ), .ZN(_00853_ ) );
NOR2_X1 _16895_ ( .A1(_00853_ ), .A2(_00784_ ), .ZN(\myifu.data_in [2] ) );
OR2_X1 _16896_ ( .A1(_00786_ ), .A2(\io_master_rdata [28] ), .ZN(_00854_ ) );
OR3_X1 _16897_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00855_ ) );
OAI211_X1 _16898_ ( .A(_02368_ ), .B(_00855_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00856_ ) );
AND3_X1 _16899_ ( .A1(_00854_ ), .A2(_00856_ ), .A3(_00804_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16900_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00857_ ) );
OAI211_X1 _16901_ ( .A(_00782_ ), .B(_00857_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00858_ ) );
OAI21_X1 _16902_ ( .A(_00858_ ), .B1(\io_master_rdata [1] ), .B2(_00832_ ), .ZN(_00859_ ) );
NOR2_X1 _16903_ ( .A1(_00859_ ), .A2(_00784_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16904_ ( .A1(_00777_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00813_ ), .ZN(_00860_ ) );
OAI211_X1 _16905_ ( .A(_02368_ ), .B(_00860_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(_00815_ ), .ZN(_00861_ ) );
OAI21_X1 _16906_ ( .A(_00861_ ), .B1(\io_master_rdata [0] ), .B2(_00832_ ), .ZN(_00862_ ) );
NOR2_X1 _16907_ ( .A1(_00862_ ), .A2(_00784_ ), .ZN(\myifu.data_in [0] ) );
OR2_X1 _16908_ ( .A1(_00832_ ), .A2(\io_master_rdata [27] ), .ZN(_00863_ ) );
OR3_X1 _16909_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00864_ ) );
OAI211_X1 _16910_ ( .A(_02369_ ), .B(_00864_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00865_ ) );
AND3_X1 _16911_ ( .A1(_00863_ ), .A2(_00865_ ), .A3(_06527_ ), .ZN(\myifu.data_in [27] ) );
OR2_X1 _16912_ ( .A1(_00786_ ), .A2(\io_master_rdata [26] ), .ZN(_00866_ ) );
OR3_X1 _16913_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00867_ ) );
OAI211_X1 _16914_ ( .A(_02368_ ), .B(_00867_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00815_ ), .ZN(_00868_ ) );
AND3_X1 _16915_ ( .A1(_00866_ ), .A2(_00868_ ), .A3(_06527_ ), .ZN(\myifu.data_in [26] ) );
OR2_X1 _16916_ ( .A1(_00832_ ), .A2(\io_master_rdata [25] ), .ZN(_00869_ ) );
OR3_X1 _16917_ ( .A1(_02320_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00809_ ), .ZN(_00870_ ) );
OAI211_X1 _16918_ ( .A(_02369_ ), .B(_00870_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00871_ ) );
AND3_X1 _16919_ ( .A1(_00869_ ), .A2(_00871_ ), .A3(_06527_ ), .ZN(\myifu.data_in [25] ) );
OR2_X1 _16920_ ( .A1(_00786_ ), .A2(\io_master_rdata [24] ), .ZN(_00872_ ) );
OR3_X1 _16921_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00813_ ), .ZN(_00873_ ) );
OAI211_X1 _16922_ ( .A(_02368_ ), .B(_00873_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00874_ ) );
AND3_X1 _16923_ ( .A1(_00872_ ), .A2(_00874_ ), .A3(_06527_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16924_ ( .A1(_02319_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06547_ ), .ZN(_00875_ ) );
OAI211_X1 _16925_ ( .A(_02367_ ), .B(_00875_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06548_ ), .ZN(_00876_ ) );
OAI21_X1 _16926_ ( .A(_00876_ ), .B1(\io_master_rdata [23] ), .B2(_02367_ ), .ZN(_00877_ ) );
NOR2_X1 _16927_ ( .A1(_00877_ ), .A2(_06516_ ), .ZN(\myifu.data_in [23] ) );
OR2_X1 _16928_ ( .A1(_00781_ ), .A2(\io_master_rdata [22] ), .ZN(_00878_ ) );
OR3_X1 _16929_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00778_ ), .ZN(_00879_ ) );
OAI211_X1 _16930_ ( .A(_00786_ ), .B(_00879_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06549_ ), .ZN(_00880_ ) );
AND3_X1 _16931_ ( .A1(_00878_ ), .A2(_00880_ ), .A3(_06527_ ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16932_ ( .A(_00242_ ), .ZN(_00881_ ) );
NAND2_X1 _16933_ ( .A1(_00881_ ), .A2(_02357_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16934_ ( .A1(_06346_ ), .A2(fanout_net_8 ), .ZN(_00882_ ) );
INV_X1 _16935_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00883_ ) );
OAI21_X1 _16936_ ( .A(_02357_ ), .B1(_00882_ ), .B2(_00883_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16937_ ( .A1(_06355_ ), .A2(fanout_net_12 ), .ZN(_00884_ ) );
OAI21_X1 _16938_ ( .A(_02357_ ), .B1(_00884_ ), .B2(_00883_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16939_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .ZN(_00885_ ) );
OAI21_X1 _16940_ ( .A(_02357_ ), .B1(_00885_ ), .B2(_00883_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
OAI21_X1 _16941_ ( .A(\IF_ID_inst [8] ), .B1(_05996_ ), .B2(_05988_ ), .ZN(_00886_ ) );
NOR2_X1 _16942_ ( .A1(_05996_ ), .A2(_05988_ ), .ZN(_00887_ ) );
AND2_X1 _16943_ ( .A1(_00887_ ), .A2(_06008_ ), .ZN(_00888_ ) );
NOR4_X1 _16944_ ( .A1(_05941_ ), .A2(_05943_ ), .A3(_05783_ ), .A4(_05836_ ), .ZN(_00889_ ) );
NAND3_X1 _16945_ ( .A1(_00888_ ), .A2(_00889_ ), .A3(_05869_ ), .ZN(_00890_ ) );
AND2_X1 _16946_ ( .A1(_00890_ ), .A2(_06144_ ), .ZN(_00891_ ) );
OAI221_X1 _16947_ ( .A(_00886_ ), .B1(_05924_ ), .B2(_05701_ ), .C1(_00891_ ), .C2(_05707_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
AND3_X1 _16948_ ( .A1(_06048_ ), .A2(\IF_ID_inst [31] ), .A3(_05724_ ), .ZN(_00892_ ) );
INV_X1 _16949_ ( .A(_00892_ ), .ZN(_00893_ ) );
BUF_X2 _16950_ ( .A(_05970_ ), .Z(_00894_ ) );
OAI221_X1 _16951_ ( .A(_00893_ ), .B1(_05702_ ), .B2(_00888_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
NOR2_X1 _16952_ ( .A1(_05970_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00895_ ) );
NOR2_X1 _16953_ ( .A1(_00887_ ), .A2(_05702_ ), .ZN(_00896_ ) );
NOR2_X1 _16954_ ( .A1(_00895_ ), .A2(_00896_ ), .ZN(_00897_ ) );
BUF_X4 _16955_ ( .A(_00897_ ), .Z(_00898_ ) );
BUF_X4 _16956_ ( .A(_00893_ ), .Z(_00899_ ) );
BUF_X4 _16957_ ( .A(_06008_ ), .Z(_00900_ ) );
OAI211_X1 _16958_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05706_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16959_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05707_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16960_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05710_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
OAI21_X1 _16961_ ( .A(\IF_ID_inst [31] ), .B1(_05996_ ), .B2(_05988_ ), .ZN(_00901_ ) );
OAI221_X1 _16962_ ( .A(_00901_ ), .B1(_05793_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI221_X1 _16963_ ( .A(_00901_ ), .B1(_05794_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI221_X1 _16964_ ( .A(_00901_ ), .B1(_05795_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16965_ ( .A(_00901_ ), .B1(_05924_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _16966_ ( .A(_00901_ ), .B1(_05760_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16967_ ( .A(_00901_ ), .B1(_05814_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16968_ ( .A(_00901_ ), .B1(_05754_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16969_ ( .A(_00901_ ), .B1(_05749_ ), .B2(_05790_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16970_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05711_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
AOI22_X1 _16971_ ( .A1(\IF_ID_inst [31] ), .A2(_05996_ ), .B1(_05988_ ), .B2(\IF_ID_inst [7] ), .ZN(_00902_ ) );
OAI211_X1 _16972_ ( .A(_06123_ ), .B(_00902_ ), .C1(_00894_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
OAI221_X1 _16973_ ( .A(_06116_ ), .B1(_00887_ ), .B2(_05706_ ), .C1(_05970_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
OAI21_X1 _16974_ ( .A(\IF_ID_inst [29] ), .B1(_05996_ ), .B2(_05988_ ), .ZN(_00903_ ) );
OAI221_X1 _16975_ ( .A(_00903_ ), .B1(_05711_ ), .B2(_06144_ ), .C1(_05970_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16976_ ( .A(_06108_ ), .ZN(_00904_ ) );
OAI221_X1 _16977_ ( .A(_00904_ ), .B1(_00887_ ), .B2(_05712_ ), .C1(_05970_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
INV_X1 _16978_ ( .A(_06101_ ), .ZN(_00905_ ) );
OAI221_X1 _16979_ ( .A(_00905_ ), .B1(_00887_ ), .B2(_05713_ ), .C1(_05970_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
OAI221_X1 _16980_ ( .A(_06063_ ), .B1(_00887_ ), .B2(_05714_ ), .C1(_05970_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
OAI21_X1 _16981_ ( .A(\IF_ID_inst [25] ), .B1(_05996_ ), .B2(_05988_ ), .ZN(_00906_ ) );
OAI221_X1 _16982_ ( .A(_00906_ ), .B1(_05715_ ), .B2(_06144_ ), .C1(_05970_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16983_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05712_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16984_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05713_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16985_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05714_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16986_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05715_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16987_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05716_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16988_ ( .A(_00898_ ), .B(_00899_ ), .C1(_05717_ ), .C2(_00900_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16989_ ( .A(_00897_ ), .B(_00893_ ), .C1(_05719_ ), .C2(_06008_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16990_ ( .A(\IF_ID_inst [11] ), .B1(_05996_ ), .B2(_05988_ ), .ZN(_00907_ ) );
OAI221_X1 _16991_ ( .A(_00907_ ), .B1(_05793_ ), .B2(_05700_ ), .C1(_00891_ ), .C2(_05716_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16992_ ( .A(\IF_ID_inst [10] ), .B1(_05996_ ), .B2(_05988_ ), .ZN(_00908_ ) );
OAI221_X1 _16993_ ( .A(_00908_ ), .B1(_05794_ ), .B2(_05700_ ), .C1(_00891_ ), .C2(_05717_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16994_ ( .A(\IF_ID_inst [9] ), .B1(_05996_ ), .B2(_05988_ ), .ZN(_00909_ ) );
OAI221_X1 _16995_ ( .A(_00909_ ), .B1(_05795_ ), .B2(_05700_ ), .C1(_00891_ ), .C2(_05719_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16996_ ( .A1(_05796_ ), .A2(_05726_ ), .ZN(_00910_ ) );
OAI221_X1 _16997_ ( .A(_00910_ ), .B1(_05760_ ), .B2(_05700_ ), .C1(_00890_ ), .C2(_05710_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AND2_X2 _16998_ ( .A1(_06421_ ), .A2(_06414_ ), .ZN(_00911_ ) );
BUF_X4 _16999_ ( .A(_00911_ ), .Z(_00912_ ) );
BUF_X4 _17000_ ( .A(_00912_ ), .Z(_00913_ ) );
AOI21_X1 _17001_ ( .A(\IF_ID_pc [1] ), .B1(_06423_ ), .B2(\IF_ID_pc [2] ), .ZN(_00914_ ) );
INV_X1 _17002_ ( .A(_00914_ ), .ZN(_00915_ ) );
OAI21_X1 _17003_ ( .A(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .B1(_06423_ ), .B2(\IF_ID_pc [2] ), .ZN(_00916_ ) );
NOR2_X1 _17004_ ( .A1(_00915_ ), .A2(_00916_ ), .ZN(_00917_ ) );
BUF_X4 _17005_ ( .A(_00917_ ), .Z(_00918_ ) );
BUF_X4 _17006_ ( .A(_00918_ ), .Z(_00919_ ) );
NAND2_X1 _17007_ ( .A1(_00833_ ), .A2(_00835_ ), .ZN(_00920_ ) );
BUF_X4 _17008_ ( .A(_06515_ ), .Z(_00921_ ) );
OAI211_X1 _17009_ ( .A(_00913_ ), .B(_00919_ ), .C1(_00920_ ), .C2(_00921_ ), .ZN(_00922_ ) );
AND2_X2 _17010_ ( .A1(_00911_ ), .A2(_00917_ ), .ZN(_00923_ ) );
OAI211_X1 _17011_ ( .A(_00922_ ), .B(\myifu.state [2] ), .C1(_00923_ ), .C2(_06087_ ), .ZN(_00924_ ) );
AND3_X1 _17012_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00925_ ) );
AND3_X1 _17013_ ( .A1(_06345_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00926_ ) );
AOI211_X1 _17014_ ( .A(_00925_ ), .B(_00926_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_06504_ ), .ZN(_00927_ ) );
NAND2_X1 _17015_ ( .A1(_00883_ ), .A2(\IF_ID_pc [2] ), .ZN(_00928_ ) );
BUF_X2 _17016_ ( .A(_00928_ ), .Z(_00929_ ) );
NAND2_X1 _17017_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00930_ ) );
BUF_X4 _17018_ ( .A(_00930_ ), .Z(_00931_ ) );
BUF_X4 _17019_ ( .A(_00931_ ), .Z(_00932_ ) );
NAND3_X1 _17020_ ( .A1(_06355_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00933_ ) );
NAND4_X1 _17021_ ( .A1(_00927_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_00933_ ), .ZN(_00934_ ) );
NOR2_X1 _17022_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00935_ ) );
BUF_X2 _17023_ ( .A(_00935_ ), .Z(_00936_ ) );
BUF_X4 _17024_ ( .A(_00936_ ), .Z(_00937_ ) );
BUF_X4 _17025_ ( .A(_06095_ ), .Z(_00938_ ) );
BUF_X4 _17026_ ( .A(_00938_ ), .Z(_00939_ ) );
NAND3_X1 _17027_ ( .A1(_00939_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00940_ ) );
NAND3_X1 _17028_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00941_ ) );
AND2_X1 _17029_ ( .A1(_00940_ ), .A2(_00941_ ), .ZN(_00942_ ) );
NAND2_X1 _17030_ ( .A1(_00928_ ), .A2(_00930_ ), .ZN(_00943_ ) );
BUF_X2 _17031_ ( .A(_00943_ ), .Z(_00944_ ) );
BUF_X4 _17032_ ( .A(_06353_ ), .Z(_00945_ ) );
BUF_X4 _17033_ ( .A(_00945_ ), .Z(_00946_ ) );
NAND3_X1 _17034_ ( .A1(_00946_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00947_ ) );
BUF_X4 _17035_ ( .A(_06354_ ), .Z(_00948_ ) );
NAND3_X1 _17036_ ( .A1(_06346_ ), .A2(_00948_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00949_ ) );
NAND4_X1 _17037_ ( .A1(_00942_ ), .A2(_00944_ ), .A3(_00947_ ), .A4(_00949_ ), .ZN(_00950_ ) );
NAND3_X1 _17038_ ( .A1(_00934_ ), .A2(_00937_ ), .A3(_00950_ ), .ZN(_00951_ ) );
NAND2_X1 _17039_ ( .A1(_00924_ ), .A2(_00951_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _17040_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00952_ ) );
AND3_X1 _17041_ ( .A1(_00938_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00953_ ) );
BUF_X4 _17042_ ( .A(_06503_ ), .Z(_00954_ ) );
AOI211_X1 _17043_ ( .A(_00952_ ), .B(_00953_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00954_ ), .ZN(_00955_ ) );
BUF_X4 _17044_ ( .A(_00928_ ), .Z(_00956_ ) );
NAND3_X1 _17045_ ( .A1(_00948_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00957_ ) );
NAND4_X1 _17046_ ( .A1(_00955_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_00957_ ), .ZN(_00958_ ) );
BUF_X4 _17047_ ( .A(_06095_ ), .Z(_00959_ ) );
BUF_X4 _17048_ ( .A(_00959_ ), .Z(_00960_ ) );
NAND3_X1 _17049_ ( .A1(_00960_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00961_ ) );
NAND3_X1 _17050_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00962_ ) );
AND2_X1 _17051_ ( .A1(_00961_ ), .A2(_00962_ ), .ZN(_00963_ ) );
BUF_X4 _17052_ ( .A(_00943_ ), .Z(_00964_ ) );
NAND3_X1 _17053_ ( .A1(_00945_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00965_ ) );
NAND3_X1 _17054_ ( .A1(_00939_ ), .A2(_00945_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00966_ ) );
NAND4_X1 _17055_ ( .A1(_00963_ ), .A2(_00964_ ), .A3(_00965_ ), .A4(_00966_ ), .ZN(_00967_ ) );
NAND3_X1 _17056_ ( .A1(_00958_ ), .A2(_00936_ ), .A3(_00967_ ), .ZN(_00968_ ) );
INV_X2 _17057_ ( .A(_00923_ ), .ZN(_00969_ ) );
BUF_X4 _17058_ ( .A(_00969_ ), .Z(_00970_ ) );
NOR2_X1 _17059_ ( .A1(_00970_ ), .A2(\myifu.data_in [31] ), .ZN(_00971_ ) );
OAI21_X1 _17060_ ( .A(\myifu.state [2] ), .B1(_00923_ ), .B2(_06130_ ), .ZN(_00972_ ) );
OAI21_X1 _17061_ ( .A(_00968_ ), .B1(_00971_ ), .B2(_00972_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
INV_X1 _17062_ ( .A(\myifu.state [2] ), .ZN(_00973_ ) );
BUF_X4 _17063_ ( .A(_00973_ ), .Z(_00974_ ) );
AOI21_X1 _17064_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_00975_ ) );
BUF_X4 _17065_ ( .A(_00912_ ), .Z(_00976_ ) );
BUF_X4 _17066_ ( .A(_00918_ ), .Z(_00977_ ) );
BUF_X4 _17067_ ( .A(_06515_ ), .Z(_00978_ ) );
OAI211_X1 _17068_ ( .A(_00976_ ), .B(_00977_ ), .C1(_00783_ ), .C2(_00978_ ), .ZN(_00979_ ) );
NAND2_X1 _17069_ ( .A1(_00975_ ), .A2(_00979_ ), .ZN(_00980_ ) );
AND3_X1 _17070_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00981_ ) );
AND3_X1 _17071_ ( .A1(_06345_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00982_ ) );
AOI211_X1 _17072_ ( .A(_00981_ ), .B(_00982_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_06504_ ), .ZN(_00983_ ) );
NAND3_X1 _17073_ ( .A1(_06355_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00984_ ) );
NAND4_X1 _17074_ ( .A1(_00983_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_00984_ ), .ZN(_00985_ ) );
NAND3_X1 _17075_ ( .A1(_00939_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00986_ ) );
NAND3_X1 _17076_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00987_ ) );
AND2_X1 _17077_ ( .A1(_00986_ ), .A2(_00987_ ), .ZN(_00988_ ) );
NAND3_X1 _17078_ ( .A1(_00946_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00989_ ) );
NAND3_X1 _17079_ ( .A1(_06346_ ), .A2(_00948_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00990_ ) );
NAND4_X1 _17080_ ( .A1(_00988_ ), .A2(_00944_ ), .A3(_00989_ ), .A4(_00990_ ), .ZN(_00991_ ) );
NAND3_X1 _17081_ ( .A1(_00985_ ), .A2(_00937_ ), .A3(_00991_ ), .ZN(_00992_ ) );
NAND2_X1 _17082_ ( .A1(_00980_ ), .A2(_00992_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
NAND2_X1 _17083_ ( .A1(_00785_ ), .A2(_00788_ ), .ZN(_00993_ ) );
OAI211_X1 _17084_ ( .A(_00912_ ), .B(_00918_ ), .C1(_00993_ ), .C2(_06515_ ), .ZN(_00994_ ) );
NAND2_X1 _17085_ ( .A1(_00994_ ), .A2(\myifu.state [2] ), .ZN(_00995_ ) );
BUF_X4 _17086_ ( .A(_00969_ ), .Z(_00996_ ) );
AOI21_X1 _17087_ ( .A(_00995_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00996_ ), .ZN(_00997_ ) );
AND3_X1 _17088_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00998_ ) );
AND3_X1 _17089_ ( .A1(_00959_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00999_ ) );
AOI211_X1 _17090_ ( .A(_00998_ ), .B(_00999_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_00954_ ), .ZN(_01000_ ) );
BUF_X4 _17091_ ( .A(_06353_ ), .Z(_01001_ ) );
NAND3_X1 _17092_ ( .A1(_01001_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_01002_ ) );
NAND4_X1 _17093_ ( .A1(_01000_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_01002_ ), .ZN(_01003_ ) );
NAND3_X1 _17094_ ( .A1(_00938_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_01004_ ) );
NAND3_X1 _17095_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_01005_ ) );
AND2_X1 _17096_ ( .A1(_01004_ ), .A2(_01005_ ), .ZN(_01006_ ) );
NAND3_X1 _17097_ ( .A1(_06354_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_01007_ ) );
BUF_X4 _17098_ ( .A(_06352_ ), .Z(_01008_ ) );
NAND3_X1 _17099_ ( .A1(_00960_ ), .A2(_01008_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_01009_ ) );
NAND4_X1 _17100_ ( .A1(_01006_ ), .A2(_00964_ ), .A3(_01007_ ), .A4(_01009_ ), .ZN(_01010_ ) );
AND3_X1 _17101_ ( .A1(_01003_ ), .A2(_00936_ ), .A3(_01010_ ), .ZN(_01011_ ) );
OR2_X1 _17102_ ( .A1(_00997_ ), .A2(_01011_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
NAND2_X1 _17103_ ( .A1(_00789_ ), .A2(_00791_ ), .ZN(_01012_ ) );
OAI211_X1 _17104_ ( .A(_00912_ ), .B(_00918_ ), .C1(_01012_ ), .C2(_06515_ ), .ZN(_01013_ ) );
NAND2_X1 _17105_ ( .A1(_01013_ ), .A2(\myifu.state [2] ), .ZN(_01014_ ) );
AOI21_X1 _17106_ ( .A(_01014_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00996_ ), .ZN(_01015_ ) );
AND3_X1 _17107_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_01016_ ) );
AND3_X1 _17108_ ( .A1(_00959_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_01017_ ) );
AOI211_X1 _17109_ ( .A(_01016_ ), .B(_01017_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_00954_ ), .ZN(_01018_ ) );
NAND3_X1 _17110_ ( .A1(_01001_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_01019_ ) );
NAND4_X1 _17111_ ( .A1(_01018_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_01019_ ), .ZN(_01020_ ) );
NAND3_X1 _17112_ ( .A1(_00938_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_01021_ ) );
NAND3_X1 _17113_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_01022_ ) );
AND2_X1 _17114_ ( .A1(_01021_ ), .A2(_01022_ ), .ZN(_01023_ ) );
BUF_X4 _17115_ ( .A(_00943_ ), .Z(_01024_ ) );
NAND3_X1 _17116_ ( .A1(_06354_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_01025_ ) );
BUF_X4 _17117_ ( .A(_00959_ ), .Z(_01026_ ) );
NAND3_X1 _17118_ ( .A1(_01026_ ), .A2(_01008_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_01027_ ) );
NAND4_X1 _17119_ ( .A1(_01023_ ), .A2(_01024_ ), .A3(_01025_ ), .A4(_01027_ ), .ZN(_01028_ ) );
AND3_X1 _17120_ ( .A1(_01020_ ), .A2(_00936_ ), .A3(_01028_ ), .ZN(_01029_ ) );
OR2_X1 _17121_ ( .A1(_01015_ ), .A2(_01029_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
NAND2_X1 _17122_ ( .A1(_00792_ ), .A2(_00794_ ), .ZN(_01030_ ) );
OAI211_X1 _17123_ ( .A(_00912_ ), .B(_00918_ ), .C1(_01030_ ), .C2(_06515_ ), .ZN(_01031_ ) );
NAND2_X1 _17124_ ( .A1(_01031_ ), .A2(\myifu.state [2] ), .ZN(_01032_ ) );
AOI21_X1 _17125_ ( .A(_01032_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00996_ ), .ZN(_01033_ ) );
AND3_X1 _17126_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_01034_ ) );
AND3_X1 _17127_ ( .A1(_00959_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_01035_ ) );
AOI211_X1 _17128_ ( .A(_01034_ ), .B(_01035_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_00954_ ), .ZN(_01036_ ) );
NAND3_X1 _17129_ ( .A1(_01001_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_01037_ ) );
NAND4_X1 _17130_ ( .A1(_01036_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_01037_ ), .ZN(_01038_ ) );
NAND3_X1 _17131_ ( .A1(_00938_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_01039_ ) );
NAND3_X1 _17132_ ( .A1(fanout_net_12 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_01040_ ) );
AND2_X1 _17133_ ( .A1(_01039_ ), .A2(_01040_ ), .ZN(_01041_ ) );
NAND3_X1 _17134_ ( .A1(_06354_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_01042_ ) );
NAND3_X1 _17135_ ( .A1(_01026_ ), .A2(_01008_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_01043_ ) );
NAND4_X1 _17136_ ( .A1(_01041_ ), .A2(_01024_ ), .A3(_01042_ ), .A4(_01043_ ), .ZN(_01044_ ) );
AND3_X1 _17137_ ( .A1(_01038_ ), .A2(_00936_ ), .A3(_01044_ ), .ZN(_01045_ ) );
OR2_X1 _17138_ ( .A1(_01033_ ), .A2(_01045_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
AOI21_X1 _17139_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01046_ ) );
NAND2_X1 _17140_ ( .A1(_00795_ ), .A2(_00797_ ), .ZN(_01047_ ) );
OAI211_X1 _17141_ ( .A(_00976_ ), .B(_00977_ ), .C1(_01047_ ), .C2(_00978_ ), .ZN(_01048_ ) );
NAND2_X1 _17142_ ( .A1(_01046_ ), .A2(_01048_ ), .ZN(_01049_ ) );
AND3_X1 _17143_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_01050_ ) );
AND3_X1 _17144_ ( .A1(_06345_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_01051_ ) );
AOI211_X1 _17145_ ( .A(_01050_ ), .B(_01051_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_06504_ ), .ZN(_01052_ ) );
NAND3_X1 _17146_ ( .A1(_06355_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_01053_ ) );
NAND4_X1 _17147_ ( .A1(_01052_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_01053_ ), .ZN(_01054_ ) );
NAND3_X1 _17148_ ( .A1(_00939_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_01055_ ) );
NAND3_X1 _17149_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_01056_ ) );
AND2_X1 _17150_ ( .A1(_01055_ ), .A2(_01056_ ), .ZN(_01057_ ) );
NAND3_X1 _17151_ ( .A1(_00946_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_01058_ ) );
NAND3_X1 _17152_ ( .A1(_06346_ ), .A2(_00948_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_01059_ ) );
NAND4_X1 _17153_ ( .A1(_01057_ ), .A2(_00944_ ), .A3(_01058_ ), .A4(_01059_ ), .ZN(_01060_ ) );
NAND3_X1 _17154_ ( .A1(_01054_ ), .A2(_00937_ ), .A3(_01060_ ), .ZN(_01061_ ) );
NAND2_X1 _17155_ ( .A1(_01049_ ), .A2(_01061_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
NAND2_X1 _17156_ ( .A1(_00798_ ), .A2(_00800_ ), .ZN(_01062_ ) );
OAI211_X1 _17157_ ( .A(_00912_ ), .B(_00918_ ), .C1(_01062_ ), .C2(_06515_ ), .ZN(_01063_ ) );
NAND2_X1 _17158_ ( .A1(_01063_ ), .A2(\myifu.state [2] ), .ZN(_01064_ ) );
AOI21_X1 _17159_ ( .A(_01064_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00996_ ), .ZN(_01065_ ) );
AND3_X1 _17160_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_01066_ ) );
AND3_X1 _17161_ ( .A1(_06344_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_01067_ ) );
AOI211_X1 _17162_ ( .A(_01066_ ), .B(_01067_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_00954_ ), .ZN(_01068_ ) );
NAND3_X1 _17163_ ( .A1(_01001_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_01069_ ) );
NAND4_X1 _17164_ ( .A1(_01068_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_01069_ ), .ZN(_01070_ ) );
NAND3_X1 _17165_ ( .A1(_00938_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_01071_ ) );
NAND3_X1 _17166_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_01072_ ) );
AND2_X1 _17167_ ( .A1(_01071_ ), .A2(_01072_ ), .ZN(_01073_ ) );
NAND3_X1 _17168_ ( .A1(_06354_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_01074_ ) );
NAND3_X1 _17169_ ( .A1(_01026_ ), .A2(_01008_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_01075_ ) );
NAND4_X1 _17170_ ( .A1(_01073_ ), .A2(_01024_ ), .A3(_01074_ ), .A4(_01075_ ), .ZN(_01076_ ) );
AND3_X1 _17171_ ( .A1(_01070_ ), .A2(_00936_ ), .A3(_01076_ ), .ZN(_01077_ ) );
OR2_X1 _17172_ ( .A1(_01065_ ), .A2(_01077_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
AOI21_X1 _17173_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01078_ ) );
NAND2_X1 _17174_ ( .A1(_00801_ ), .A2(_00803_ ), .ZN(_01079_ ) );
OAI211_X1 _17175_ ( .A(_00976_ ), .B(_00977_ ), .C1(_01079_ ), .C2(_00978_ ), .ZN(_01080_ ) );
NAND2_X1 _17176_ ( .A1(_01078_ ), .A2(_01080_ ), .ZN(_01081_ ) );
AND3_X1 _17177_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_01082_ ) );
AND3_X1 _17178_ ( .A1(_06345_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_01083_ ) );
AOI211_X1 _17179_ ( .A(_01082_ ), .B(_01083_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_06504_ ), .ZN(_01084_ ) );
NAND3_X1 _17180_ ( .A1(_06355_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_01085_ ) );
NAND4_X1 _17181_ ( .A1(_01084_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_01085_ ), .ZN(_01086_ ) );
BUF_X4 _17182_ ( .A(_00938_ ), .Z(_01087_ ) );
NAND3_X1 _17183_ ( .A1(_01087_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_01088_ ) );
NAND3_X1 _17184_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_01089_ ) );
AND2_X1 _17185_ ( .A1(_01088_ ), .A2(_01089_ ), .ZN(_01090_ ) );
BUF_X4 _17186_ ( .A(_00964_ ), .Z(_01091_ ) );
NAND3_X1 _17187_ ( .A1(_00946_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_01092_ ) );
NAND3_X1 _17188_ ( .A1(_06346_ ), .A2(_00948_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_01093_ ) );
NAND4_X1 _17189_ ( .A1(_01090_ ), .A2(_01091_ ), .A3(_01092_ ), .A4(_01093_ ), .ZN(_01094_ ) );
NAND3_X1 _17190_ ( .A1(_01086_ ), .A2(_00937_ ), .A3(_01094_ ), .ZN(_01095_ ) );
NAND2_X1 _17191_ ( .A1(_01081_ ), .A2(_01095_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
OAI211_X1 _17192_ ( .A(_00912_ ), .B(_00918_ ), .C1(_00807_ ), .C2(_06515_ ), .ZN(_01096_ ) );
NAND2_X1 _17193_ ( .A1(_01096_ ), .A2(\myifu.state [2] ), .ZN(_01097_ ) );
AOI21_X1 _17194_ ( .A(_01097_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00996_ ), .ZN(_01098_ ) );
AND3_X1 _17195_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_01099_ ) );
AND3_X1 _17196_ ( .A1(_06344_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_01100_ ) );
AOI211_X1 _17197_ ( .A(_01099_ ), .B(_01100_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_06503_ ), .ZN(_01101_ ) );
NAND3_X1 _17198_ ( .A1(_01001_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_01102_ ) );
NAND4_X1 _17199_ ( .A1(_01101_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_01102_ ), .ZN(_01103_ ) );
NAND3_X1 _17200_ ( .A1(_00938_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_01104_ ) );
NAND3_X1 _17201_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_01105_ ) );
AND2_X1 _17202_ ( .A1(_01104_ ), .A2(_01105_ ), .ZN(_01106_ ) );
NAND3_X1 _17203_ ( .A1(_06354_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_01107_ ) );
NAND3_X1 _17204_ ( .A1(_01026_ ), .A2(_06353_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_01108_ ) );
NAND4_X1 _17205_ ( .A1(_01106_ ), .A2(_01024_ ), .A3(_01107_ ), .A4(_01108_ ), .ZN(_01109_ ) );
AND3_X1 _17206_ ( .A1(_01103_ ), .A2(_00936_ ), .A3(_01109_ ), .ZN(_01110_ ) );
OR2_X1 _17207_ ( .A1(_01098_ ), .A2(_01110_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
NAND2_X1 _17208_ ( .A1(_00808_ ), .A2(_00811_ ), .ZN(_01111_ ) );
OAI211_X1 _17209_ ( .A(_00912_ ), .B(_00918_ ), .C1(_01111_ ), .C2(_06515_ ), .ZN(_01112_ ) );
NAND2_X1 _17210_ ( .A1(_01112_ ), .A2(\myifu.state [2] ), .ZN(_01113_ ) );
AOI21_X1 _17211_ ( .A(_01113_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00969_ ), .ZN(_01114_ ) );
AND3_X1 _17212_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_01115_ ) );
AND3_X1 _17213_ ( .A1(_06344_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_01116_ ) );
AOI211_X1 _17214_ ( .A(_01115_ ), .B(_01116_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_06503_ ), .ZN(_01117_ ) );
NAND3_X1 _17215_ ( .A1(_01001_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_01118_ ) );
NAND4_X1 _17216_ ( .A1(_01117_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_01118_ ), .ZN(_01119_ ) );
NAND3_X1 _17217_ ( .A1(_00938_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_01120_ ) );
NAND3_X1 _17218_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_01121_ ) );
AND2_X1 _17219_ ( .A1(_01120_ ), .A2(_01121_ ), .ZN(_01122_ ) );
NAND3_X1 _17220_ ( .A1(_01008_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_01123_ ) );
NAND3_X1 _17221_ ( .A1(_01026_ ), .A2(_06353_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_01124_ ) );
NAND4_X1 _17222_ ( .A1(_01122_ ), .A2(_01024_ ), .A3(_01123_ ), .A4(_01124_ ), .ZN(_01125_ ) );
AND3_X1 _17223_ ( .A1(_01119_ ), .A2(_00936_ ), .A3(_01125_ ), .ZN(_01126_ ) );
OR2_X1 _17224_ ( .A1(_01114_ ), .A2(_01126_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
AOI21_X1 _17225_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01127_ ) );
NAND2_X1 _17226_ ( .A1(_00812_ ), .A2(_00816_ ), .ZN(_01128_ ) );
OAI211_X1 _17227_ ( .A(_00976_ ), .B(_00977_ ), .C1(_01128_ ), .C2(_00978_ ), .ZN(_01129_ ) );
NAND2_X1 _17228_ ( .A1(_01127_ ), .A2(_01129_ ), .ZN(_01130_ ) );
AND3_X1 _17229_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_01131_ ) );
AND3_X1 _17230_ ( .A1(_06345_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_01132_ ) );
AOI211_X1 _17231_ ( .A(_01131_ ), .B(_01132_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_06504_ ), .ZN(_01133_ ) );
NAND3_X1 _17232_ ( .A1(_06355_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_01134_ ) );
NAND4_X1 _17233_ ( .A1(_01133_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_01134_ ), .ZN(_01135_ ) );
NAND3_X1 _17234_ ( .A1(_01087_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_01136_ ) );
NAND3_X1 _17235_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_01137_ ) );
AND2_X1 _17236_ ( .A1(_01136_ ), .A2(_01137_ ), .ZN(_01138_ ) );
NAND3_X1 _17237_ ( .A1(_00946_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_01139_ ) );
BUF_X4 _17238_ ( .A(_00960_ ), .Z(_01140_ ) );
BUF_X4 _17239_ ( .A(_06354_ ), .Z(_01141_ ) );
NAND3_X1 _17240_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_01142_ ) );
NAND4_X1 _17241_ ( .A1(_01138_ ), .A2(_01091_ ), .A3(_01139_ ), .A4(_01142_ ), .ZN(_01143_ ) );
NAND3_X1 _17242_ ( .A1(_01135_ ), .A2(_00937_ ), .A3(_01143_ ), .ZN(_01144_ ) );
NAND2_X1 _17243_ ( .A1(_01130_ ), .A2(_01144_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
NAND2_X1 _17244_ ( .A1(_00817_ ), .A2(_00819_ ), .ZN(_01145_ ) );
OAI211_X1 _17245_ ( .A(_00912_ ), .B(_00918_ ), .C1(_01145_ ), .C2(_06515_ ), .ZN(_01146_ ) );
NAND2_X1 _17246_ ( .A1(_01146_ ), .A2(\myifu.state [2] ), .ZN(_01147_ ) );
AOI21_X1 _17247_ ( .A(_01147_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00969_ ), .ZN(_01148_ ) );
AND3_X1 _17248_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_01149_ ) );
AND3_X1 _17249_ ( .A1(_06344_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_01150_ ) );
AOI211_X1 _17250_ ( .A(_01149_ ), .B(_01150_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_06503_ ), .ZN(_01151_ ) );
NAND3_X1 _17251_ ( .A1(_01001_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_01152_ ) );
NAND4_X1 _17252_ ( .A1(_01151_ ), .A2(_00956_ ), .A3(_00930_ ), .A4(_01152_ ), .ZN(_01153_ ) );
NAND3_X1 _17253_ ( .A1(_00959_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_01154_ ) );
NAND3_X1 _17254_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_01155_ ) );
AND2_X1 _17255_ ( .A1(_01154_ ), .A2(_01155_ ), .ZN(_01156_ ) );
NAND3_X1 _17256_ ( .A1(_01008_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_01157_ ) );
NAND3_X1 _17257_ ( .A1(_01026_ ), .A2(_06353_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_01158_ ) );
NAND4_X1 _17258_ ( .A1(_01156_ ), .A2(_01024_ ), .A3(_01157_ ), .A4(_01158_ ), .ZN(_01159_ ) );
AND3_X1 _17259_ ( .A1(_01153_ ), .A2(_00936_ ), .A3(_01159_ ), .ZN(_01160_ ) );
OR2_X1 _17260_ ( .A1(_01148_ ), .A2(_01160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
NAND2_X1 _17261_ ( .A1(_00820_ ), .A2(_00822_ ), .ZN(_01161_ ) );
OAI211_X1 _17262_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01161_ ), .C2(_00921_ ), .ZN(_01162_ ) );
OAI211_X1 _17263_ ( .A(_01162_ ), .B(\myifu.state [2] ), .C1(_00923_ ), .C2(_06057_ ), .ZN(_01163_ ) );
AND3_X1 _17264_ ( .A1(fanout_net_13 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_01164_ ) );
AND3_X1 _17265_ ( .A1(_06345_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_01165_ ) );
AOI211_X1 _17266_ ( .A(_01164_ ), .B(_01165_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_06504_ ), .ZN(_01166_ ) );
BUF_X4 _17267_ ( .A(_00945_ ), .Z(_01167_ ) );
NAND3_X1 _17268_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_01168_ ) );
NAND4_X1 _17269_ ( .A1(_01166_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_01168_ ), .ZN(_01169_ ) );
NAND3_X1 _17270_ ( .A1(_01087_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_01170_ ) );
NAND3_X1 _17271_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_01171_ ) );
AND2_X1 _17272_ ( .A1(_01170_ ), .A2(_01171_ ), .ZN(_01172_ ) );
BUF_X4 _17273_ ( .A(_01001_ ), .Z(_01173_ ) );
NAND3_X1 _17274_ ( .A1(_01173_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_01174_ ) );
NAND3_X1 _17275_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_01175_ ) );
NAND4_X1 _17276_ ( .A1(_01172_ ), .A2(_01091_ ), .A3(_01174_ ), .A4(_01175_ ), .ZN(_01176_ ) );
NAND3_X1 _17277_ ( .A1(_01169_ ), .A2(_00937_ ), .A3(_01176_ ), .ZN(_01177_ ) );
NAND2_X1 _17278_ ( .A1(_01163_ ), .A2(_01177_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AOI21_X1 _17279_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_01178_ ) );
NAND2_X1 _17280_ ( .A1(_00823_ ), .A2(_00825_ ), .ZN(_01179_ ) );
OAI211_X1 _17281_ ( .A(_00976_ ), .B(_00977_ ), .C1(_01179_ ), .C2(_00978_ ), .ZN(_01180_ ) );
NAND2_X1 _17282_ ( .A1(_01178_ ), .A2(_01180_ ), .ZN(_01181_ ) );
AND3_X1 _17283_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_01182_ ) );
AND3_X1 _17284_ ( .A1(_06345_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_01183_ ) );
BUF_X4 _17285_ ( .A(_00954_ ), .Z(_01184_ ) );
AOI211_X1 _17286_ ( .A(_01182_ ), .B(_01183_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_01184_ ), .ZN(_01185_ ) );
NAND3_X1 _17287_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_01186_ ) );
NAND4_X1 _17288_ ( .A1(_01185_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_01186_ ), .ZN(_01187_ ) );
NAND3_X1 _17289_ ( .A1(_01087_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_01188_ ) );
NAND3_X1 _17290_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_01189_ ) );
AND2_X1 _17291_ ( .A1(_01188_ ), .A2(_01189_ ), .ZN(_01190_ ) );
NAND3_X1 _17292_ ( .A1(_01173_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_01191_ ) );
NAND3_X1 _17293_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_01192_ ) );
NAND4_X1 _17294_ ( .A1(_01190_ ), .A2(_01091_ ), .A3(_01191_ ), .A4(_01192_ ), .ZN(_01193_ ) );
NAND3_X1 _17295_ ( .A1(_01187_ ), .A2(_00937_ ), .A3(_01193_ ), .ZN(_01194_ ) );
NAND2_X1 _17296_ ( .A1(_01181_ ), .A2(_01194_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
NAND2_X1 _17297_ ( .A1(_00826_ ), .A2(_00828_ ), .ZN(_01195_ ) );
OAI211_X1 _17298_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01195_ ), .C2(_00921_ ), .ZN(_01196_ ) );
OAI211_X1 _17299_ ( .A(_01196_ ), .B(\myifu.state [2] ), .C1(_00923_ ), .C2(_06076_ ), .ZN(_01197_ ) );
AND3_X1 _17300_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_01198_ ) );
AND3_X1 _17301_ ( .A1(_06345_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_01199_ ) );
AOI211_X1 _17302_ ( .A(_01198_ ), .B(_01199_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_01184_ ), .ZN(_01200_ ) );
NAND3_X1 _17303_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_01201_ ) );
NAND4_X1 _17304_ ( .A1(_01200_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_01201_ ), .ZN(_01202_ ) );
NAND3_X1 _17305_ ( .A1(_01087_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_01203_ ) );
NAND3_X1 _17306_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_01204_ ) );
AND2_X1 _17307_ ( .A1(_01203_ ), .A2(_01204_ ), .ZN(_01205_ ) );
NAND3_X1 _17308_ ( .A1(_01173_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_01206_ ) );
NAND3_X1 _17309_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_01207_ ) );
NAND4_X1 _17310_ ( .A1(_01205_ ), .A2(_01091_ ), .A3(_01206_ ), .A4(_01207_ ), .ZN(_01208_ ) );
NAND3_X1 _17311_ ( .A1(_01202_ ), .A2(_00937_ ), .A3(_01208_ ), .ZN(_01209_ ) );
NAND2_X1 _17312_ ( .A1(_01197_ ), .A2(_01209_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
AOI21_X1 _17313_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_01210_ ) );
NAND2_X1 _17314_ ( .A1(_00829_ ), .A2(_00831_ ), .ZN(_01211_ ) );
OAI211_X1 _17315_ ( .A(_00976_ ), .B(_00977_ ), .C1(_01211_ ), .C2(_00978_ ), .ZN(_01212_ ) );
NAND2_X1 _17316_ ( .A1(_01210_ ), .A2(_01212_ ), .ZN(_01213_ ) );
AND3_X1 _17317_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_01214_ ) );
AND3_X1 _17318_ ( .A1(_06345_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_01215_ ) );
AOI211_X1 _17319_ ( .A(_01214_ ), .B(_01215_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_01184_ ), .ZN(_01216_ ) );
NAND3_X1 _17320_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_01217_ ) );
NAND4_X1 _17321_ ( .A1(_01216_ ), .A2(_00929_ ), .A3(_00932_ ), .A4(_01217_ ), .ZN(_01218_ ) );
NAND3_X1 _17322_ ( .A1(_01087_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_01219_ ) );
NAND3_X1 _17323_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_01220_ ) );
AND2_X1 _17324_ ( .A1(_01219_ ), .A2(_01220_ ), .ZN(_01221_ ) );
NAND3_X1 _17325_ ( .A1(_01173_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_01222_ ) );
NAND3_X1 _17326_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_01223_ ) );
NAND4_X1 _17327_ ( .A1(_01221_ ), .A2(_01091_ ), .A3(_01222_ ), .A4(_01223_ ), .ZN(_01224_ ) );
NAND3_X1 _17328_ ( .A1(_01218_ ), .A2(_00937_ ), .A3(_01224_ ), .ZN(_01225_ ) );
NAND2_X1 _17329_ ( .A1(_01213_ ), .A2(_01225_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
AOI21_X1 _17330_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_01226_ ) );
OAI211_X1 _17331_ ( .A(_00976_ ), .B(_00977_ ), .C1(_00838_ ), .C2(_00978_ ), .ZN(_01227_ ) );
NAND2_X1 _17332_ ( .A1(_01226_ ), .A2(_01227_ ), .ZN(_01228_ ) );
AND3_X1 _17333_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_01229_ ) );
CLKBUF_X2 _17334_ ( .A(_06344_ ), .Z(_01230_ ) );
AND3_X1 _17335_ ( .A1(_01230_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_01231_ ) );
AOI211_X1 _17336_ ( .A(_01229_ ), .B(_01231_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_01184_ ), .ZN(_01232_ ) );
BUF_X4 _17337_ ( .A(_00956_ ), .Z(_01233_ ) );
BUF_X4 _17338_ ( .A(_00931_ ), .Z(_01234_ ) );
NAND3_X1 _17339_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_01235_ ) );
NAND4_X1 _17340_ ( .A1(_01232_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01235_ ), .ZN(_01236_ ) );
NAND3_X1 _17341_ ( .A1(_01087_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_01237_ ) );
NAND3_X1 _17342_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_01238_ ) );
AND2_X1 _17343_ ( .A1(_01237_ ), .A2(_01238_ ), .ZN(_01239_ ) );
NAND3_X1 _17344_ ( .A1(_01173_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_01240_ ) );
NAND3_X1 _17345_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_01241_ ) );
NAND4_X1 _17346_ ( .A1(_01239_ ), .A2(_01091_ ), .A3(_01240_ ), .A4(_01241_ ), .ZN(_01242_ ) );
NAND3_X1 _17347_ ( .A1(_01236_ ), .A2(_00937_ ), .A3(_01242_ ), .ZN(_01243_ ) );
NAND2_X1 _17348_ ( .A1(_01228_ ), .A2(_01243_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AOI21_X1 _17349_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01244_ ) );
OAI211_X1 _17350_ ( .A(_00976_ ), .B(_00977_ ), .C1(_00841_ ), .C2(_00978_ ), .ZN(_01245_ ) );
NAND2_X1 _17351_ ( .A1(_01244_ ), .A2(_01245_ ), .ZN(_01246_ ) );
AND3_X1 _17352_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_01247_ ) );
AND3_X1 _17353_ ( .A1(_01230_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_01248_ ) );
AOI211_X1 _17354_ ( .A(_01247_ ), .B(_01248_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_01184_ ), .ZN(_01249_ ) );
NAND3_X1 _17355_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_01250_ ) );
NAND4_X1 _17356_ ( .A1(_01249_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01250_ ), .ZN(_01251_ ) );
BUF_X4 _17357_ ( .A(_00936_ ), .Z(_01252_ ) );
NAND3_X1 _17358_ ( .A1(_01087_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_01253_ ) );
NAND3_X1 _17359_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_01254_ ) );
AND2_X1 _17360_ ( .A1(_01253_ ), .A2(_01254_ ), .ZN(_01255_ ) );
NAND3_X1 _17361_ ( .A1(_01173_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_01256_ ) );
NAND3_X1 _17362_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_01257_ ) );
NAND4_X1 _17363_ ( .A1(_01255_ ), .A2(_01091_ ), .A3(_01256_ ), .A4(_01257_ ), .ZN(_01258_ ) );
NAND3_X1 _17364_ ( .A1(_01251_ ), .A2(_01252_ ), .A3(_01258_ ), .ZN(_01259_ ) );
NAND2_X1 _17365_ ( .A1(_01246_ ), .A2(_01259_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
AOI21_X1 _17366_ ( .A(_00974_ ), .B1(_00970_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01260_ ) );
OAI211_X1 _17367_ ( .A(_00976_ ), .B(_00977_ ), .C1(_00844_ ), .C2(_00978_ ), .ZN(_01261_ ) );
NAND2_X1 _17368_ ( .A1(_01260_ ), .A2(_01261_ ), .ZN(_01262_ ) );
AND3_X1 _17369_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_01263_ ) );
AND3_X1 _17370_ ( .A1(_01230_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_01264_ ) );
AOI211_X1 _17371_ ( .A(_01263_ ), .B(_01264_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_01184_ ), .ZN(_01265_ ) );
NAND3_X1 _17372_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_01266_ ) );
NAND4_X1 _17373_ ( .A1(_01265_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01266_ ), .ZN(_01267_ ) );
NAND3_X1 _17374_ ( .A1(_01087_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_01268_ ) );
NAND3_X1 _17375_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_01269_ ) );
AND2_X1 _17376_ ( .A1(_01268_ ), .A2(_01269_ ), .ZN(_01270_ ) );
NAND3_X1 _17377_ ( .A1(_01173_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_01271_ ) );
NAND3_X1 _17378_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_01272_ ) );
NAND4_X1 _17379_ ( .A1(_01270_ ), .A2(_01091_ ), .A3(_01271_ ), .A4(_01272_ ), .ZN(_01273_ ) );
NAND3_X1 _17380_ ( .A1(_01267_ ), .A2(_01252_ ), .A3(_01273_ ), .ZN(_01274_ ) );
NAND2_X1 _17381_ ( .A1(_01262_ ), .A2(_01274_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
AOI21_X1 _17382_ ( .A(_00974_ ), .B1(_00996_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01275_ ) );
OAI211_X1 _17383_ ( .A(_00976_ ), .B(_00977_ ), .C1(_00847_ ), .C2(_00978_ ), .ZN(_01276_ ) );
NAND2_X1 _17384_ ( .A1(_01275_ ), .A2(_01276_ ), .ZN(_01277_ ) );
AND3_X1 _17385_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_01278_ ) );
AND3_X1 _17386_ ( .A1(_01230_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_01279_ ) );
AOI211_X1 _17387_ ( .A(_01278_ ), .B(_01279_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_01184_ ), .ZN(_01280_ ) );
NAND3_X1 _17388_ ( .A1(_01167_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_01281_ ) );
NAND4_X1 _17389_ ( .A1(_01280_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01281_ ), .ZN(_01282_ ) );
NAND3_X1 _17390_ ( .A1(_01087_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_01283_ ) );
NAND3_X1 _17391_ ( .A1(fanout_net_14 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_01284_ ) );
AND2_X1 _17392_ ( .A1(_01283_ ), .A2(_01284_ ), .ZN(_01285_ ) );
NAND3_X1 _17393_ ( .A1(_01173_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_01286_ ) );
NAND3_X1 _17394_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_01287_ ) );
NAND4_X1 _17395_ ( .A1(_01285_ ), .A2(_01091_ ), .A3(_01286_ ), .A4(_01287_ ), .ZN(_01288_ ) );
NAND3_X1 _17396_ ( .A1(_01282_ ), .A2(_01252_ ), .A3(_01288_ ), .ZN(_01289_ ) );
NAND2_X1 _17397_ ( .A1(_01277_ ), .A2(_01289_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _17398_ ( .A(_00973_ ), .B1(_00996_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01290_ ) );
OAI211_X1 _17399_ ( .A(_00913_ ), .B(_00919_ ), .C1(_00850_ ), .C2(_00921_ ), .ZN(_01291_ ) );
NAND2_X1 _17400_ ( .A1(_01290_ ), .A2(_01291_ ), .ZN(_01292_ ) );
AND3_X1 _17401_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_01293_ ) );
AND3_X1 _17402_ ( .A1(_01230_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_01294_ ) );
AOI211_X1 _17403_ ( .A(_01293_ ), .B(_01294_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_01184_ ), .ZN(_01295_ ) );
NAND3_X1 _17404_ ( .A1(_01167_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_01296_ ) );
NAND4_X1 _17405_ ( .A1(_01295_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01296_ ), .ZN(_01297_ ) );
NAND3_X1 _17406_ ( .A1(_00960_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_01298_ ) );
NAND3_X1 _17407_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_01299_ ) );
AND2_X1 _17408_ ( .A1(_01298_ ), .A2(_01299_ ), .ZN(_01300_ ) );
NAND3_X1 _17409_ ( .A1(_01173_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_01301_ ) );
NAND3_X1 _17410_ ( .A1(_01140_ ), .A2(_01141_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_01302_ ) );
NAND4_X1 _17411_ ( .A1(_01300_ ), .A2(_00964_ ), .A3(_01301_ ), .A4(_01302_ ), .ZN(_01303_ ) );
NAND3_X1 _17412_ ( .A1(_01297_ ), .A2(_01252_ ), .A3(_01303_ ), .ZN(_01304_ ) );
NAND2_X1 _17413_ ( .A1(_01292_ ), .A2(_01304_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
OAI211_X1 _17414_ ( .A(_00912_ ), .B(_00918_ ), .C1(_00853_ ), .C2(_02293_ ), .ZN(_01305_ ) );
NAND2_X1 _17415_ ( .A1(_01305_ ), .A2(\myifu.state [2] ), .ZN(_01306_ ) );
AOI21_X1 _17416_ ( .A(_01306_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00969_ ), .ZN(_01307_ ) );
AND3_X1 _17417_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_01308_ ) );
AND3_X1 _17418_ ( .A1(_06344_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_01309_ ) );
AOI211_X1 _17419_ ( .A(_01308_ ), .B(_01309_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_06503_ ), .ZN(_01310_ ) );
NAND3_X1 _17420_ ( .A1(_01001_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_01311_ ) );
NAND4_X1 _17421_ ( .A1(_01310_ ), .A2(_00928_ ), .A3(_00930_ ), .A4(_01311_ ), .ZN(_01312_ ) );
NAND3_X1 _17422_ ( .A1(_00959_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_01313_ ) );
NAND3_X1 _17423_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_01314_ ) );
AND2_X1 _17424_ ( .A1(_01313_ ), .A2(_01314_ ), .ZN(_01315_ ) );
NAND3_X1 _17425_ ( .A1(_01008_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_01316_ ) );
NAND3_X1 _17426_ ( .A1(_01026_ ), .A2(_06353_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_01317_ ) );
NAND4_X1 _17427_ ( .A1(_01315_ ), .A2(_01024_ ), .A3(_01316_ ), .A4(_01317_ ), .ZN(_01318_ ) );
AND3_X1 _17428_ ( .A1(_01312_ ), .A2(_00935_ ), .A3(_01318_ ), .ZN(_01319_ ) );
OR2_X1 _17429_ ( .A1(_01307_ ), .A2(_01319_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
OAI211_X1 _17430_ ( .A(_00911_ ), .B(_00917_ ), .C1(_00859_ ), .C2(_02293_ ), .ZN(_01320_ ) );
NAND2_X1 _17431_ ( .A1(_01320_ ), .A2(\myifu.state [2] ), .ZN(_01321_ ) );
AOI21_X1 _17432_ ( .A(_01321_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00969_ ), .ZN(_01322_ ) );
AND3_X1 _17433_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01323_ ) );
AND3_X1 _17434_ ( .A1(_06344_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01324_ ) );
AOI211_X1 _17435_ ( .A(_01323_ ), .B(_01324_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_06503_ ), .ZN(_01325_ ) );
NAND3_X1 _17436_ ( .A1(_01001_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01326_ ) );
NAND4_X1 _17437_ ( .A1(_01325_ ), .A2(_00928_ ), .A3(_00930_ ), .A4(_01326_ ), .ZN(_01327_ ) );
NAND3_X1 _17438_ ( .A1(_00959_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01328_ ) );
NAND3_X1 _17439_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01329_ ) );
AND2_X1 _17440_ ( .A1(_01328_ ), .A2(_01329_ ), .ZN(_01330_ ) );
NAND3_X1 _17441_ ( .A1(_01008_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01331_ ) );
NAND3_X1 _17442_ ( .A1(_01026_ ), .A2(_06353_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01332_ ) );
NAND4_X1 _17443_ ( .A1(_01330_ ), .A2(_01024_ ), .A3(_01331_ ), .A4(_01332_ ), .ZN(_01333_ ) );
AND3_X1 _17444_ ( .A1(_01327_ ), .A2(_00935_ ), .A3(_01333_ ), .ZN(_01334_ ) );
OR2_X1 _17445_ ( .A1(_01322_ ), .A2(_01334_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
NAND2_X1 _17446_ ( .A1(_00854_ ), .A2(_00856_ ), .ZN(_01335_ ) );
OAI211_X1 _17447_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01335_ ), .C2(_00921_ ), .ZN(_01336_ ) );
OAI211_X1 _17448_ ( .A(_01336_ ), .B(\myifu.state [2] ), .C1(_00923_ ), .C2(_06109_ ), .ZN(_01337_ ) );
AND3_X1 _17449_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01338_ ) );
AND3_X1 _17450_ ( .A1(_01230_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01339_ ) );
AOI211_X1 _17451_ ( .A(_01338_ ), .B(_01339_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_01184_ ), .ZN(_01340_ ) );
NAND3_X1 _17452_ ( .A1(_01167_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01341_ ) );
NAND4_X1 _17453_ ( .A1(_01340_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01341_ ), .ZN(_01342_ ) );
NAND3_X1 _17454_ ( .A1(_00960_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01343_ ) );
NAND3_X1 _17455_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01344_ ) );
AND2_X1 _17456_ ( .A1(_01343_ ), .A2(_01344_ ), .ZN(_01345_ ) );
NAND3_X1 _17457_ ( .A1(_01173_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01346_ ) );
NAND3_X1 _17458_ ( .A1(_00939_ ), .A2(_00945_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01347_ ) );
NAND4_X1 _17459_ ( .A1(_01345_ ), .A2(_00964_ ), .A3(_01346_ ), .A4(_01347_ ), .ZN(_01348_ ) );
NAND3_X1 _17460_ ( .A1(_01342_ ), .A2(_01252_ ), .A3(_01348_ ), .ZN(_01349_ ) );
NAND2_X1 _17461_ ( .A1(_01337_ ), .A2(_01349_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
OAI211_X1 _17462_ ( .A(_00911_ ), .B(_00917_ ), .C1(_00862_ ), .C2(_02293_ ), .ZN(_01350_ ) );
NAND2_X1 _17463_ ( .A1(_01350_ ), .A2(\myifu.state [2] ), .ZN(_01351_ ) );
AOI21_X1 _17464_ ( .A(_01351_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00969_ ), .ZN(_01352_ ) );
AND3_X1 _17465_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01353_ ) );
AND3_X1 _17466_ ( .A1(_06344_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01354_ ) );
AOI211_X1 _17467_ ( .A(_01353_ ), .B(_01354_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_06503_ ), .ZN(_01355_ ) );
NAND3_X1 _17468_ ( .A1(_06354_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01356_ ) );
NAND4_X1 _17469_ ( .A1(_01355_ ), .A2(_00928_ ), .A3(_00930_ ), .A4(_01356_ ), .ZN(_01357_ ) );
NAND3_X1 _17470_ ( .A1(_00959_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01358_ ) );
NAND3_X1 _17471_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01359_ ) );
AND2_X1 _17472_ ( .A1(_01358_ ), .A2(_01359_ ), .ZN(_01360_ ) );
NAND3_X1 _17473_ ( .A1(_01008_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01361_ ) );
NAND3_X1 _17474_ ( .A1(_01026_ ), .A2(_06353_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01362_ ) );
NAND4_X1 _17475_ ( .A1(_01360_ ), .A2(_01024_ ), .A3(_01361_ ), .A4(_01362_ ), .ZN(_01363_ ) );
AND3_X1 _17476_ ( .A1(_01357_ ), .A2(_00935_ ), .A3(_01363_ ), .ZN(_01364_ ) );
OR2_X1 _17477_ ( .A1(_01352_ ), .A2(_01364_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
NAND2_X1 _17478_ ( .A1(_00863_ ), .A2(_00865_ ), .ZN(_01365_ ) );
OAI211_X1 _17479_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01365_ ), .C2(_00921_ ), .ZN(_01366_ ) );
OAI211_X1 _17480_ ( .A(_01366_ ), .B(\myifu.state [2] ), .C1(_00923_ ), .C2(_06102_ ), .ZN(_01367_ ) );
AND3_X1 _17481_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01368_ ) );
AND3_X1 _17482_ ( .A1(_01230_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01369_ ) );
AOI211_X1 _17483_ ( .A(_01368_ ), .B(_01369_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_01184_ ), .ZN(_01370_ ) );
NAND3_X1 _17484_ ( .A1(_00946_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01371_ ) );
NAND4_X1 _17485_ ( .A1(_01370_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01371_ ), .ZN(_01372_ ) );
NAND3_X1 _17486_ ( .A1(_00960_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01373_ ) );
NAND3_X1 _17487_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01374_ ) );
AND2_X1 _17488_ ( .A1(_01373_ ), .A2(_01374_ ), .ZN(_01375_ ) );
NAND3_X1 _17489_ ( .A1(_00948_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01376_ ) );
NAND3_X1 _17490_ ( .A1(_00939_ ), .A2(_00945_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01377_ ) );
NAND4_X1 _17491_ ( .A1(_01375_ ), .A2(_00964_ ), .A3(_01376_ ), .A4(_01377_ ), .ZN(_01378_ ) );
NAND3_X1 _17492_ ( .A1(_01372_ ), .A2(_01252_ ), .A3(_01378_ ), .ZN(_01379_ ) );
NAND2_X1 _17493_ ( .A1(_01367_ ), .A2(_01379_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
AOI21_X1 _17494_ ( .A(_00973_ ), .B1(_00996_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_01380_ ) );
NAND2_X1 _17495_ ( .A1(_00866_ ), .A2(_00868_ ), .ZN(_01381_ ) );
OAI211_X1 _17496_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01381_ ), .C2(_00921_ ), .ZN(_01382_ ) );
NAND2_X1 _17497_ ( .A1(_01380_ ), .A2(_01382_ ), .ZN(_01383_ ) );
AND3_X1 _17498_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01384_ ) );
AND3_X1 _17499_ ( .A1(_01230_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01385_ ) );
AOI211_X1 _17500_ ( .A(_01384_ ), .B(_01385_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_00954_ ), .ZN(_01386_ ) );
NAND3_X1 _17501_ ( .A1(_00946_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01387_ ) );
NAND4_X1 _17502_ ( .A1(_01386_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01387_ ), .ZN(_01388_ ) );
NAND3_X1 _17503_ ( .A1(_00960_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01389_ ) );
NAND3_X1 _17504_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01390_ ) );
AND2_X1 _17505_ ( .A1(_01389_ ), .A2(_01390_ ), .ZN(_01391_ ) );
NAND3_X1 _17506_ ( .A1(_00948_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01392_ ) );
NAND3_X1 _17507_ ( .A1(_00939_ ), .A2(_00945_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01393_ ) );
NAND4_X1 _17508_ ( .A1(_01391_ ), .A2(_00964_ ), .A3(_01392_ ), .A4(_01393_ ), .ZN(_01394_ ) );
NAND3_X1 _17509_ ( .A1(_01388_ ), .A2(_01252_ ), .A3(_01394_ ), .ZN(_01395_ ) );
NAND2_X1 _17510_ ( .A1(_01383_ ), .A2(_01395_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
NAND2_X1 _17511_ ( .A1(_00869_ ), .A2(_00871_ ), .ZN(_01396_ ) );
OAI211_X1 _17512_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01396_ ), .C2(_00921_ ), .ZN(_01397_ ) );
OAI211_X1 _17513_ ( .A(_01397_ ), .B(\myifu.state [2] ), .C1(_00923_ ), .C2(_06068_ ), .ZN(_01398_ ) );
AND3_X1 _17514_ ( .A1(fanout_net_15 ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01399_ ) );
AND3_X1 _17515_ ( .A1(_01230_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01400_ ) );
AOI211_X1 _17516_ ( .A(_01399_ ), .B(_01400_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00954_ ), .ZN(_01401_ ) );
NAND3_X1 _17517_ ( .A1(_00946_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01402_ ) );
NAND4_X1 _17518_ ( .A1(_01401_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01402_ ), .ZN(_01403_ ) );
NAND3_X1 _17519_ ( .A1(_00960_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01404_ ) );
NAND3_X1 _17520_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01405_ ) );
AND2_X1 _17521_ ( .A1(_01404_ ), .A2(_01405_ ), .ZN(_01406_ ) );
NAND3_X1 _17522_ ( .A1(_00948_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01407_ ) );
NAND3_X1 _17523_ ( .A1(_00939_ ), .A2(_00945_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01408_ ) );
NAND4_X1 _17524_ ( .A1(_01406_ ), .A2(_00964_ ), .A3(_01407_ ), .A4(_01408_ ), .ZN(_01409_ ) );
NAND3_X1 _17525_ ( .A1(_01403_ ), .A2(_01252_ ), .A3(_01409_ ), .ZN(_01410_ ) );
NAND2_X1 _17526_ ( .A1(_01398_ ), .A2(_01410_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
AOI21_X1 _17527_ ( .A(_00973_ ), .B1(_00996_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01411_ ) );
NAND2_X1 _17528_ ( .A1(_00872_ ), .A2(_00874_ ), .ZN(_01412_ ) );
OAI211_X1 _17529_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01412_ ), .C2(_00921_ ), .ZN(_01413_ ) );
NAND2_X1 _17530_ ( .A1(_01411_ ), .A2(_01413_ ), .ZN(_01414_ ) );
AND3_X1 _17531_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01415_ ) );
AND3_X1 _17532_ ( .A1(_01230_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01416_ ) );
AOI211_X1 _17533_ ( .A(_01415_ ), .B(_01416_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_00954_ ), .ZN(_01417_ ) );
NAND3_X1 _17534_ ( .A1(_00946_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01418_ ) );
NAND4_X1 _17535_ ( .A1(_01417_ ), .A2(_01233_ ), .A3(_01234_ ), .A4(_01418_ ), .ZN(_01419_ ) );
NAND3_X1 _17536_ ( .A1(_00960_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01420_ ) );
NAND3_X1 _17537_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01421_ ) );
AND2_X1 _17538_ ( .A1(_01420_ ), .A2(_01421_ ), .ZN(_01422_ ) );
NAND3_X1 _17539_ ( .A1(_00948_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01423_ ) );
NAND3_X1 _17540_ ( .A1(_00939_ ), .A2(_00945_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01424_ ) );
NAND4_X1 _17541_ ( .A1(_01422_ ), .A2(_00964_ ), .A3(_01423_ ), .A4(_01424_ ), .ZN(_01425_ ) );
NAND3_X1 _17542_ ( .A1(_01419_ ), .A2(_01252_ ), .A3(_01425_ ), .ZN(_01426_ ) );
NAND2_X1 _17543_ ( .A1(_01414_ ), .A2(_01426_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
OAI211_X1 _17544_ ( .A(_00911_ ), .B(_00917_ ), .C1(_00877_ ), .C2(_02293_ ), .ZN(_01427_ ) );
NAND2_X1 _17545_ ( .A1(_01427_ ), .A2(\myifu.state [2] ), .ZN(_01428_ ) );
AOI21_X1 _17546_ ( .A(_01428_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00969_ ), .ZN(_01429_ ) );
AND3_X1 _17547_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01430_ ) );
AND3_X1 _17548_ ( .A1(_06344_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01431_ ) );
AOI211_X1 _17549_ ( .A(_01430_ ), .B(_01431_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_06503_ ), .ZN(_01432_ ) );
NAND3_X1 _17550_ ( .A1(_06354_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01433_ ) );
NAND4_X1 _17551_ ( .A1(_01432_ ), .A2(_00928_ ), .A3(_00930_ ), .A4(_01433_ ), .ZN(_01434_ ) );
NAND3_X1 _17552_ ( .A1(_00959_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01435_ ) );
NAND3_X1 _17553_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01436_ ) );
AND2_X1 _17554_ ( .A1(_01435_ ), .A2(_01436_ ), .ZN(_01437_ ) );
NAND3_X1 _17555_ ( .A1(_01008_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01438_ ) );
NAND3_X1 _17556_ ( .A1(_01026_ ), .A2(_06353_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01439_ ) );
NAND4_X1 _17557_ ( .A1(_01437_ ), .A2(_01024_ ), .A3(_01438_ ), .A4(_01439_ ), .ZN(_01440_ ) );
AND3_X1 _17558_ ( .A1(_01434_ ), .A2(_00935_ ), .A3(_01440_ ), .ZN(_01441_ ) );
OR2_X1 _17559_ ( .A1(_01429_ ), .A2(_01441_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
AOI21_X1 _17560_ ( .A(_00973_ ), .B1(_00996_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_01442_ ) );
NAND2_X1 _17561_ ( .A1(_00878_ ), .A2(_00880_ ), .ZN(_01443_ ) );
OAI211_X1 _17562_ ( .A(_00913_ ), .B(_00919_ ), .C1(_01443_ ), .C2(_00921_ ), .ZN(_01444_ ) );
NAND2_X1 _17563_ ( .A1(_01442_ ), .A2(_01444_ ), .ZN(_01445_ ) );
AND3_X1 _17564_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01446_ ) );
AND3_X1 _17565_ ( .A1(_00938_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01447_ ) );
AOI211_X1 _17566_ ( .A(_01446_ ), .B(_01447_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_00954_ ), .ZN(_01448_ ) );
NAND3_X1 _17567_ ( .A1(_00946_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01449_ ) );
NAND4_X1 _17568_ ( .A1(_01448_ ), .A2(_00956_ ), .A3(_00931_ ), .A4(_01449_ ), .ZN(_01450_ ) );
NAND3_X1 _17569_ ( .A1(_00960_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01451_ ) );
NAND3_X1 _17570_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01452_ ) );
AND2_X1 _17571_ ( .A1(_01451_ ), .A2(_01452_ ), .ZN(_01453_ ) );
NAND3_X1 _17572_ ( .A1(_00948_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01454_ ) );
NAND3_X1 _17573_ ( .A1(_00939_ ), .A2(_00945_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01455_ ) );
NAND4_X1 _17574_ ( .A1(_01453_ ), .A2(_00964_ ), .A3(_01454_ ), .A4(_01455_ ), .ZN(_01456_ ) );
NAND3_X1 _17575_ ( .A1(_01450_ ), .A2(_01252_ ), .A3(_01456_ ), .ZN(_01457_ ) );
NAND2_X1 _17576_ ( .A1(_01445_ ), .A2(_01457_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI211_X1 _17577_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_05916_ ), .C1(_06257_ ), .C2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _17578_ ( .A1(_06421_ ), .A2(_06414_ ), .A3(\myifu.state [2] ), .A4(_06415_ ), .ZN(_01458_ ) );
NOR2_X1 _17579_ ( .A1(_02246_ ), .A2(_00773_ ), .ZN(_01459_ ) );
INV_X1 _17580_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01460_ ) );
AOI21_X1 _17581_ ( .A(_00771_ ), .B1(_01459_ ), .B2(_01460_ ), .ZN(_01461_ ) );
AOI21_X1 _17582_ ( .A(reset ), .B1(_01458_ ), .B2(_01461_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _17583_ ( .A1(_05675_ ), .A2(_02293_ ), .ZN(_01462_ ) );
AND3_X1 _17584_ ( .A1(_02112_ ), .A2(_02204_ ), .A3(_02245_ ), .ZN(_01463_ ) );
NOR4_X1 _17585_ ( .A1(_01462_ ), .A2(\myidu.stall_quest_fencei ), .A3(_00773_ ), .A4(_01463_ ), .ZN(_01464_ ) );
AND2_X1 _17586_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01465_ ) );
OR4_X1 _17587_ ( .A1(reset ), .A2(_01464_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A4(_01465_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _17588_ ( .A1(_06422_ ), .A2(_03400_ ), .A3(\myifu.state [2] ), .ZN(_01466_ ) );
NAND2_X1 _17589_ ( .A1(_01462_ ), .A2(_02371_ ), .ZN(_01467_ ) );
NAND2_X1 _17590_ ( .A1(_01466_ ), .A2(_01467_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _17591_ ( .A1(_06421_ ), .A2(_06414_ ), .A3(\myifu.state [2] ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17592_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01468_ ) );
NOR3_X1 _17593_ ( .A1(_01468_ ), .A2(_00884_ ), .A3(_00944_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NOR3_X1 _17594_ ( .A1(_01468_ ), .A2(_00885_ ), .A3(_00944_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _17595_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00944_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17596_ ( .A1(\IF_ID_pc [4] ), .A2(_06502_ ), .A3(_06355_ ), .A4(_00944_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
NOR3_X1 _17597_ ( .A1(_01468_ ), .A2(_00882_ ), .A3(_00944_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17598_ ( .A1(_06346_ ), .A2(_06502_ ), .A3(\IF_ID_pc [3] ), .A4(_00944_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
AND3_X1 _17599_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06504_ ), .A3(_00944_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17600_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06504_ ), .A3(_00929_ ), .A4(_00932_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
AND3_X1 _17601_ ( .A1(_02357_ ), .A2(_06504_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
AND3_X1 _17602_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06346_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
AND3_X1 _17603_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_06355_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
AND3_X1 _17604_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
NOR3_X1 _17605_ ( .A1(_05917_ ), .A2(_00771_ ), .A3(_01465_ ), .ZN(_01469_ ) );
NAND3_X1 _17606_ ( .A1(_00773_ ), .A2(_05916_ ), .A3(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01470_ ) );
NAND2_X1 _17607_ ( .A1(_01469_ ), .A2(_01470_ ), .ZN(_01471_ ) );
AOI211_X1 _17608_ ( .A(_01459_ ), .B(_01471_ ), .C1(_06422_ ), .C2(_02248_ ), .ZN(_01472_ ) );
OR2_X1 _17609_ ( .A1(_01462_ ), .A2(_00773_ ), .ZN(_01473_ ) );
AND2_X1 _17610_ ( .A1(_01472_ ), .A2(_01473_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17611_ ( .A1(_06252_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_05918_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
AOI21_X1 _17612_ ( .A(_05920_ ), .B1(_05701_ ), .B2(_05972_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
AOI211_X1 _17613_ ( .A(reset ), .B(_01471_ ), .C1(_02246_ ), .C2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _17614_ ( .A(_06432_ ), .B(_05678_ ), .S(\mylsu.state [0] ), .Z(_01474_ ) );
AOI21_X1 _17615_ ( .A(_01474_ ), .B1(_06573_ ), .B2(\mylsu.state [3] ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17616_ ( .A(_06498_ ), .ZN(_01475_ ) );
AOI211_X1 _17617_ ( .A(_01475_ ), .B(_01474_ ), .C1(_06573_ ), .C2(\mylsu.state [3] ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
NOR2_X1 _17618_ ( .A1(_05680_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01476_ ) );
AND3_X1 _17619_ ( .A1(_05677_ ), .A2(\mylsu.state [0] ), .A3(_01476_ ), .ZN(_01477_ ) );
NAND3_X1 _17620_ ( .A1(_01477_ ), .A2(_02343_ ), .A3(_06488_ ), .ZN(_01478_ ) );
INV_X1 _17621_ ( .A(_06573_ ), .ZN(_01479_ ) );
OAI21_X1 _17622_ ( .A(_01478_ ), .B1(_01479_ ), .B2(_06497_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND2_X1 _17623_ ( .A1(_06477_ ), .A2(\mylsu.state [0] ), .ZN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
OAI211_X1 _17624_ ( .A(_06477_ ), .B(\mylsu.state [0] ), .C1(io_master_awready ), .C2(io_master_wready ), .ZN(_01480_ ) );
NOR4_X1 _17625_ ( .A1(_02325_ ), .A2(_05683_ ), .A3(_02353_ ), .A4(_01480_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
AND2_X1 _17626_ ( .A1(io_master_awready ), .A2(io_master_wready ), .ZN(_01481_ ) );
NOR2_X1 _17627_ ( .A1(_06440_ ), .A2(_01481_ ), .ZN(_01482_ ) );
AND4_X1 _17628_ ( .A1(io_master_awready ), .A2(_01482_ ), .A3(_06552_ ), .A4(_06477_ ), .ZN(_01483_ ) );
NAND4_X1 _17629_ ( .A1(_02379_ ), .A2(\mylsu.state [0] ), .A3(_02384_ ), .A4(_01483_ ), .ZN(_01484_ ) );
OR4_X1 _17630_ ( .A1(_06560_ ), .A2(_02404_ ), .A3(_06429_ ), .A4(io_master_wready ), .ZN(_01485_ ) );
NAND2_X1 _17631_ ( .A1(_01484_ ), .A2(_01485_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
INV_X1 _17632_ ( .A(_06440_ ), .ZN(_01486_ ) );
NAND4_X1 _17633_ ( .A1(_02385_ ), .A2(_01486_ ), .A3(_06555_ ), .A4(_01481_ ), .ZN(_01487_ ) );
AOI221_X4 _17634_ ( .A(_06568_ ), .B1(\mylsu.state [2] ), .B2(io_master_wready ), .C1(\mylsu.state [4] ), .C2(io_master_awready ), .ZN(_01488_ ) );
AOI21_X1 _17635_ ( .A(_01475_ ), .B1(_01487_ ), .B2(_01488_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
NOR3_X1 _17636_ ( .A1(_05677_ ), .A2(_05678_ ), .A3(_05680_ ), .ZN(_01489_ ) );
AND3_X1 _17637_ ( .A1(_01489_ ), .A2(_02343_ ), .A3(_06488_ ), .ZN(_01490_ ) );
NOR4_X1 _17638_ ( .A1(_02324_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A4(_05680_ ), .ZN(_01491_ ) );
NAND2_X1 _17639_ ( .A1(_01491_ ), .A2(_06491_ ), .ZN(_01492_ ) );
AND2_X1 _17640_ ( .A1(_06465_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_01493_ ) );
OR3_X1 _17641_ ( .A1(_05679_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A3(_01493_ ), .ZN(_01494_ ) );
AOI21_X1 _17642_ ( .A(_01475_ ), .B1(_01492_ ), .B2(_01494_ ), .ZN(_01495_ ) );
AND2_X1 _17643_ ( .A1(_01482_ ), .A2(_06477_ ), .ZN(_01496_ ) );
INV_X1 _17644_ ( .A(_01496_ ), .ZN(_01497_ ) );
NOR4_X1 _17645_ ( .A1(_01497_ ), .A2(io_master_awready ), .A3(io_master_wready ), .A4(_05683_ ), .ZN(_01498_ ) );
AND3_X1 _17646_ ( .A1(_02379_ ), .A2(_02384_ ), .A3(_01498_ ), .ZN(_01499_ ) );
AND3_X1 _17647_ ( .A1(_02342_ ), .A2(_06498_ ), .A3(_01476_ ), .ZN(_01500_ ) );
NAND4_X1 _17648_ ( .A1(_02325_ ), .A2(EXU_valid_LSU ), .A3(_06552_ ), .A4(_06488_ ), .ZN(_01501_ ) );
NOR2_X1 _17649_ ( .A1(_01501_ ), .A2(_02353_ ), .ZN(_01502_ ) );
OR4_X1 _17650_ ( .A1(_01495_ ), .A2(_01499_ ), .A3(_01500_ ), .A4(_01502_ ), .ZN(_01503_ ) );
OAI21_X1 _17651_ ( .A(\mylsu.state [0] ), .B1(_01490_ ), .B2(_01503_ ), .ZN(_01504_ ) );
OR2_X1 _17652_ ( .A1(_06573_ ), .A2(_06497_ ), .ZN(_01505_ ) );
NAND4_X1 _17653_ ( .A1(_02381_ ), .A2(_02383_ ), .A3(_06552_ ), .A4(_06498_ ), .ZN(_01506_ ) );
NAND3_X1 _17654_ ( .A1(_01506_ ), .A2(EXU_valid_LSU ), .A3(_01486_ ), .ZN(_01507_ ) );
AOI221_X4 _17655_ ( .A(_01475_ ), .B1(\mylsu.state [1] ), .B2(_06567_ ), .C1(_01507_ ), .C2(\mylsu.state [0] ), .ZN(_01508_ ) );
NAND3_X1 _17656_ ( .A1(_01504_ ), .A2(_01505_ ), .A3(_01508_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND4_X1 _17657_ ( .A1(_02385_ ), .A2(io_master_wready ), .A3(_06555_ ), .A4(_01482_ ), .ZN(_01509_ ) );
AOI211_X1 _17658_ ( .A(io_master_awready ), .B(_01475_ ), .C1(_01509_ ), .C2(_06559_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
BUF_X4 _17659_ ( .A(_06441_ ), .Z(_01510_ ) );
AOI21_X1 _17660_ ( .A(\EX_LS_pc [21] ), .B1(_06436_ ), .B2(_01510_ ), .ZN(_01511_ ) );
BUF_X4 _17661_ ( .A(_05123_ ), .Z(_01512_ ) );
OAI21_X1 _17662_ ( .A(_06441_ ), .B1(_01512_ ), .B2(_06593_ ), .ZN(_01513_ ) );
AOI21_X1 _17663_ ( .A(_01513_ ), .B1(\LS_WB_wdata_csreg [21] ), .B2(_01512_ ), .ZN(_01514_ ) );
AOI21_X1 _17664_ ( .A(_01511_ ), .B1(_06487_ ), .B2(_01514_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
AOI221_X4 _17665_ ( .A(_06443_ ), .B1(\LS_WB_wdata_csreg [20] ), .B2(_05123_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [20] ), .ZN(_01515_ ) );
BUF_X4 _17666_ ( .A(_06436_ ), .Z(_01516_ ) );
BUF_X4 _17667_ ( .A(_06441_ ), .Z(_01517_ ) );
AOI21_X1 _17668_ ( .A(\EX_LS_pc [20] ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01518_ ) );
NOR2_X1 _17669_ ( .A1(_01515_ ), .A2(_01518_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _17670_ ( .A(\LS_WB_wdata_csreg [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_06446_ ), .Z(_01519_ ) );
MUX2_X1 _17671_ ( .A(_01519_ ), .B(\EX_LS_pc [19] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
AOI21_X1 _17672_ ( .A(\EX_LS_pc [18] ), .B1(_06487_ ), .B2(_01517_ ), .ZN(_01520_ ) );
INV_X1 _17673_ ( .A(_06441_ ), .ZN(_01521_ ) );
BUF_X4 _17674_ ( .A(_04998_ ), .Z(_01522_ ) );
MUX2_X1 _17675_ ( .A(\LS_WB_wdata_csreg [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_01522_ ), .Z(_01523_ ) );
AOI211_X1 _17676_ ( .A(_01521_ ), .B(_01523_ ), .C1(_02386_ ), .C2(_06552_ ), .ZN(_01524_ ) );
NOR2_X1 _17677_ ( .A1(_01520_ ), .A2(_01524_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _17678_ ( .A(\LS_WB_wdata_csreg [17] ), .B(\EX_LS_result_csreg_mem [17] ), .S(_06446_ ), .Z(_01525_ ) );
MUX2_X1 _17679_ ( .A(_01525_ ), .B(\EX_LS_pc [17] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _17680_ ( .A(\EX_LS_pc [16] ), .B1(_06436_ ), .B2(_01510_ ), .ZN(_01526_ ) );
OAI21_X1 _17681_ ( .A(_06441_ ), .B1(_01512_ ), .B2(_06605_ ), .ZN(_01527_ ) );
AOI21_X1 _17682_ ( .A(_01527_ ), .B1(\LS_WB_wdata_csreg [16] ), .B2(_01512_ ), .ZN(_01528_ ) );
AOI21_X1 _17683_ ( .A(_01526_ ), .B1(_06487_ ), .B2(_01528_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _17684_ ( .A(\LS_WB_wdata_csreg [15] ), .B(\EX_LS_result_csreg_mem [15] ), .S(_01522_ ), .Z(_01529_ ) );
MUX2_X1 _17685_ ( .A(_01529_ ), .B(\EX_LS_pc [15] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI221_X4 _17686_ ( .A(_06443_ ), .B1(\LS_WB_wdata_csreg [14] ), .B2(_05123_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [14] ), .ZN(_01530_ ) );
AOI21_X1 _17687_ ( .A(\EX_LS_pc [14] ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01531_ ) );
NOR2_X1 _17688_ ( .A1(_01530_ ), .A2(_01531_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _17689_ ( .A(\LS_WB_wdata_csreg [13] ), .B(\EX_LS_result_csreg_mem [13] ), .S(_01522_ ), .Z(_01532_ ) );
MUX2_X1 _17690_ ( .A(_01532_ ), .B(\EX_LS_pc [13] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
AOI221_X4 _17691_ ( .A(_06443_ ), .B1(\LS_WB_wdata_csreg [12] ), .B2(_05123_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [12] ), .ZN(_01533_ ) );
AOI21_X1 _17692_ ( .A(\EX_LS_pc [12] ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01534_ ) );
NOR2_X1 _17693_ ( .A1(_01533_ ), .A2(_01534_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI221_X4 _17694_ ( .A(_06443_ ), .B1(\LS_WB_wdata_csreg [30] ), .B2(_06480_ ), .C1(\EX_LS_result_csreg_mem [30] ), .C2(_06446_ ), .ZN(_01535_ ) );
AOI21_X1 _17695_ ( .A(\EX_LS_pc [30] ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01536_ ) );
NOR2_X1 _17696_ ( .A1(_01535_ ), .A2(_01536_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
AOI21_X1 _17697_ ( .A(\EX_LS_pc [11] ), .B1(_06436_ ), .B2(_01510_ ), .ZN(_01537_ ) );
OAI21_X1 _17698_ ( .A(_06441_ ), .B1(_01512_ ), .B2(_06866_ ), .ZN(_01538_ ) );
AOI21_X1 _17699_ ( .A(_01538_ ), .B1(\LS_WB_wdata_csreg [11] ), .B2(_01512_ ), .ZN(_01539_ ) );
AOI21_X1 _17700_ ( .A(_01537_ ), .B1(_06487_ ), .B2(_01539_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _17701_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_01522_ ), .Z(_01540_ ) );
MUX2_X1 _17702_ ( .A(_01540_ ), .B(\EX_LS_pc [10] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _17703_ ( .A(\LS_WB_wdata_csreg [9] ), .B(\EX_LS_result_csreg_mem [9] ), .S(_01522_ ), .Z(_01541_ ) );
MUX2_X1 _17704_ ( .A(_01541_ ), .B(\EX_LS_pc [9] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
AOI221_X4 _17705_ ( .A(_06443_ ), .B1(\LS_WB_wdata_csreg [8] ), .B2(_06480_ ), .C1(\EX_LS_result_csreg_mem [8] ), .C2(_06446_ ), .ZN(_01542_ ) );
AOI21_X1 _17706_ ( .A(\EX_LS_pc [8] ), .B1(_01516_ ), .B2(_01510_ ), .ZN(_01543_ ) );
NOR2_X1 _17707_ ( .A1(_01542_ ), .A2(_01543_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _17708_ ( .A(\LS_WB_wdata_csreg [7] ), .B(\EX_LS_result_csreg_mem [7] ), .S(_01522_ ), .Z(_01544_ ) );
MUX2_X1 _17709_ ( .A(_01544_ ), .B(\EX_LS_pc [7] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
AOI21_X1 _17710_ ( .A(\EX_LS_pc [6] ), .B1(_06436_ ), .B2(_01510_ ), .ZN(_01545_ ) );
OAI21_X1 _17711_ ( .A(_06441_ ), .B1(_01512_ ), .B2(_06590_ ), .ZN(_01546_ ) );
AOI21_X1 _17712_ ( .A(_01546_ ), .B1(\LS_WB_wdata_csreg [6] ), .B2(_01512_ ), .ZN(_01547_ ) );
AOI21_X1 _17713_ ( .A(_01545_ ), .B1(_06487_ ), .B2(_01547_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _17714_ ( .A(\LS_WB_wdata_csreg [5] ), .B(\EX_LS_result_csreg_mem [5] ), .S(_01522_ ), .Z(_01548_ ) );
MUX2_X1 _17715_ ( .A(_01548_ ), .B(\EX_LS_pc [5] ), .S(_06444_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
OAI22_X1 _17716_ ( .A1(_06446_ ), .A2(_02377_ ), .B1(_06451_ ), .B2(_05366_ ), .ZN(_01549_ ) );
MUX2_X1 _17717_ ( .A(_01549_ ), .B(\EX_LS_pc [4] ), .S(_06443_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
AOI21_X1 _17718_ ( .A(\EX_LS_pc [3] ), .B1(_06436_ ), .B2(_06441_ ), .ZN(_01550_ ) );
OAI21_X1 _17719_ ( .A(_06441_ ), .B1(_01512_ ), .B2(_06579_ ), .ZN(_01551_ ) );
AOI21_X1 _17720_ ( .A(_01551_ ), .B1(\LS_WB_wdata_csreg [3] ), .B2(_01512_ ), .ZN(_01552_ ) );
AOI21_X1 _17721_ ( .A(_01550_ ), .B1(_06487_ ), .B2(_01552_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
AOI221_X4 _17722_ ( .A(_06442_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [2] ), .C1(\LS_WB_wdata_csreg [2] ), .C2(_05123_ ), .ZN(_01553_ ) );
AOI21_X1 _17723_ ( .A(_01553_ ), .B1(_06430_ ), .B2(_06444_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _17724_ ( .A(\LS_WB_wdata_csreg [29] ), .B(\EX_LS_result_csreg_mem [29] ), .S(_01522_ ), .Z(_01554_ ) );
MUX2_X1 _17725_ ( .A(_01554_ ), .B(\EX_LS_pc [29] ), .S(_06443_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
AOI221_X4 _17726_ ( .A(_06443_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [1] ), .C1(\LS_WB_wdata_csreg [1] ), .C2(_05123_ ), .ZN(_01555_ ) );
AOI21_X1 _17727_ ( .A(\EX_LS_pc [1] ), .B1(_01516_ ), .B2(_01510_ ), .ZN(_01556_ ) );
NOR2_X1 _17728_ ( .A1(_01555_ ), .A2(_01556_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI221_X4 _17729_ ( .A(_06443_ ), .B1(_06480_ ), .B2(\LS_WB_wdata_csreg [0] ), .C1(\EX_LS_result_csreg_mem [0] ), .C2(_06446_ ), .ZN(_01557_ ) );
AOI21_X1 _17730_ ( .A(\EX_LS_pc [0] ), .B1(_01516_ ), .B2(_01510_ ), .ZN(_01558_ ) );
NOR2_X1 _17731_ ( .A1(_01557_ ), .A2(_01558_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
AOI21_X1 _17732_ ( .A(\EX_LS_pc [28] ), .B1(_06487_ ), .B2(_01517_ ), .ZN(_01559_ ) );
MUX2_X1 _17733_ ( .A(\LS_WB_wdata_csreg [28] ), .B(\EX_LS_result_csreg_mem [28] ), .S(_01522_ ), .Z(_01560_ ) );
AOI211_X1 _17734_ ( .A(_01521_ ), .B(_01560_ ), .C1(_02386_ ), .C2(_06552_ ), .ZN(_01561_ ) );
NOR2_X1 _17735_ ( .A1(_01559_ ), .A2(_01561_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI221_X4 _17736_ ( .A(_06442_ ), .B1(\LS_WB_wdata_csreg [27] ), .B2(_05123_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [27] ), .ZN(_01562_ ) );
AOI21_X1 _17737_ ( .A(\EX_LS_pc [27] ), .B1(_01516_ ), .B2(_01510_ ), .ZN(_01563_ ) );
NOR2_X1 _17738_ ( .A1(_01562_ ), .A2(_01563_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI21_X1 _17739_ ( .A(\EX_LS_pc [26] ), .B1(_06487_ ), .B2(_01517_ ), .ZN(_01564_ ) );
MUX2_X1 _17740_ ( .A(\LS_WB_wdata_csreg [26] ), .B(\EX_LS_result_csreg_mem [26] ), .S(_01522_ ), .Z(_01565_ ) );
AOI211_X1 _17741_ ( .A(_01521_ ), .B(_01565_ ), .C1(_02386_ ), .C2(_06552_ ), .ZN(_01566_ ) );
NOR2_X1 _17742_ ( .A1(_01564_ ), .A2(_01566_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI221_X4 _17743_ ( .A(_06442_ ), .B1(\LS_WB_wdata_csreg [25] ), .B2(_05123_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [25] ), .ZN(_01567_ ) );
AOI21_X1 _17744_ ( .A(\EX_LS_pc [25] ), .B1(_06436_ ), .B2(_01510_ ), .ZN(_01568_ ) );
NOR2_X1 _17745_ ( .A1(_01567_ ), .A2(_01568_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _17746_ ( .A(\EX_LS_pc [24] ), .B1(_06487_ ), .B2(_01517_ ), .ZN(_01569_ ) );
MUX2_X1 _17747_ ( .A(\LS_WB_wdata_csreg [24] ), .B(\EX_LS_result_csreg_mem [24] ), .S(_05048_ ), .Z(_01570_ ) );
AOI211_X1 _17748_ ( .A(_01521_ ), .B(_01570_ ), .C1(_02386_ ), .C2(_06552_ ), .ZN(_01571_ ) );
NOR2_X1 _17749_ ( .A1(_01569_ ), .A2(_01571_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _17750_ ( .A(\EX_LS_pc [23] ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01572_ ) );
MUX2_X1 _17751_ ( .A(\LS_WB_wdata_csreg [23] ), .B(\EX_LS_result_csreg_mem [23] ), .S(_05048_ ), .Z(_01573_ ) );
AOI211_X1 _17752_ ( .A(_01521_ ), .B(_01573_ ), .C1(_02386_ ), .C2(_06552_ ), .ZN(_01574_ ) );
NOR2_X1 _17753_ ( .A1(_01572_ ), .A2(_01574_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
AOI221_X4 _17754_ ( .A(_06442_ ), .B1(\LS_WB_wdata_csreg [22] ), .B2(_05123_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [22] ), .ZN(_01575_ ) );
AOI21_X1 _17755_ ( .A(\EX_LS_pc [22] ), .B1(_06436_ ), .B2(_01510_ ), .ZN(_01576_ ) );
NOR2_X1 _17756_ ( .A1(_01575_ ), .A2(_01576_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
AOI21_X1 _17757_ ( .A(\EX_LS_pc [31] ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01577_ ) );
MUX2_X1 _17758_ ( .A(\LS_WB_wdata_csreg [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_05048_ ), .Z(_01578_ ) );
AOI211_X1 _17759_ ( .A(_01521_ ), .B(_01578_ ), .C1(_02386_ ), .C2(_06552_ ), .ZN(_01579_ ) );
NOR2_X1 _17760_ ( .A1(_01577_ ), .A2(_01579_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17761_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01580_ ) );
INV_X1 _17762_ ( .A(_01580_ ), .ZN(_01581_ ) );
OR3_X1 _17763_ ( .A1(_00807_ ), .A2(_05676_ ), .A3(_01581_ ), .ZN(_01582_ ) );
NAND3_X1 _17764_ ( .A1(_00776_ ), .A2(_02270_ ), .A3(_01581_ ), .ZN(_01583_ ) );
AND2_X2 _17765_ ( .A1(_01582_ ), .A2(_01583_ ), .ZN(_01584_ ) );
AND2_X1 _17766_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01585_ ) );
INV_X1 _17767_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01586_ ) );
AND2_X2 _17768_ ( .A1(_01585_ ), .A2(_01586_ ), .ZN(_01587_ ) );
AND2_X4 _17769_ ( .A1(_01584_ ), .A2(_01587_ ), .ZN(_01588_ ) );
AND2_X1 _17770_ ( .A1(_01586_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01589_ ) );
INV_X1 _17771_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_01590_ ) );
AND2_X1 _17772_ ( .A1(_01589_ ), .A2(_01590_ ), .ZN(_01591_ ) );
NAND2_X1 _17773_ ( .A1(_01590_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01592_ ) );
NOR2_X1 _17774_ ( .A1(_01592_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01593_ ) );
OR2_X1 _17775_ ( .A1(_01591_ ), .A2(_01593_ ), .ZN(_01594_ ) );
NOR2_X4 _17776_ ( .A1(_01588_ ), .A2(_01594_ ), .ZN(_01595_ ) );
BUF_X8 _17777_ ( .A(_01595_ ), .Z(_01596_ ) );
NAND3_X1 _17778_ ( .A1(_00785_ ), .A2(_00788_ ), .A3(_06550_ ), .ZN(_01597_ ) );
AND2_X2 _17779_ ( .A1(_01585_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01598_ ) );
BUF_X4 _17780_ ( .A(_01598_ ), .Z(_01599_ ) );
NOR2_X1 _17781_ ( .A1(_01597_ ), .A2(_01599_ ), .ZN(_01600_ ) );
OAI21_X1 _17782_ ( .A(_01596_ ), .B1(_01600_ ), .B2(_01587_ ), .ZN(_01601_ ) );
INV_X2 _17783_ ( .A(_01591_ ), .ZN(_01602_ ) );
BUF_X4 _17784_ ( .A(_01602_ ), .Z(_01603_ ) );
NOR2_X2 _17785_ ( .A1(_00807_ ), .A2(_05676_ ), .ZN(_01604_ ) );
AND3_X4 _17786_ ( .A1(_01604_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(_06508_ ), .ZN(_01605_ ) );
NOR2_X1 _17787_ ( .A1(_00838_ ), .A2(_05676_ ), .ZN(_01606_ ) );
AOI21_X4 _17788_ ( .A(_01605_ ), .B1(_01580_ ), .B2(_01606_ ), .ZN(_01607_ ) );
NOR2_X1 _17789_ ( .A1(_00877_ ), .A2(_05676_ ), .ZN(_01608_ ) );
NAND3_X1 _17790_ ( .A1(_01608_ ), .A2(_06512_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01609_ ) );
AND2_X1 _17791_ ( .A1(_00776_ ), .A2(_02270_ ), .ZN(_01610_ ) );
NAND3_X1 _17792_ ( .A1(_01610_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01611_ ) );
AND3_X4 _17793_ ( .A1(_01607_ ), .A2(_01609_ ), .A3(_01611_ ), .ZN(_01612_ ) );
BUF_X8 _17794_ ( .A(_01612_ ), .Z(_01613_ ) );
BUF_X8 _17795_ ( .A(_01613_ ), .Z(_01614_ ) );
OAI21_X1 _17796_ ( .A(_01601_ ), .B1(_01603_ ), .B2(_01614_ ), .ZN(_01615_ ) );
MUX2_X1 _17797_ ( .A(\EX_LS_result_reg [21] ), .B(_01615_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
BUF_X4 _17798_ ( .A(_01587_ ), .Z(_01616_ ) );
NAND3_X1 _17799_ ( .A1(_00789_ ), .A2(_00791_ ), .A3(_06550_ ), .ZN(_01617_ ) );
NOR2_X1 _17800_ ( .A1(_01617_ ), .A2(_01599_ ), .ZN(_01618_ ) );
OAI21_X1 _17801_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01618_ ), .ZN(_01619_ ) );
OAI21_X1 _17802_ ( .A(_01619_ ), .B1(_01603_ ), .B2(_01614_ ), .ZN(_01620_ ) );
MUX2_X1 _17803_ ( .A(\EX_LS_result_reg [20] ), .B(_01620_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NOR2_X4 _17804_ ( .A1(_01613_ ), .A2(_01602_ ), .ZN(_01621_ ) );
NOR2_X2 _17805_ ( .A1(_01621_ ), .A2(_06432_ ), .ZN(_01622_ ) );
NAND3_X1 _17806_ ( .A1(_00792_ ), .A2(_00794_ ), .A3(_06550_ ), .ZN(_01623_ ) );
NOR2_X1 _17807_ ( .A1(_01623_ ), .A2(_01599_ ), .ZN(_01624_ ) );
OAI21_X1 _17808_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01624_ ), .ZN(_01625_ ) );
BUF_X4 _17809_ ( .A(_06432_ ), .Z(_01626_ ) );
AOI22_X1 _17810_ ( .A1(_01622_ ), .A2(_01625_ ), .B1(_01626_ ), .B2(_03652_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _17811_ ( .A1(_00795_ ), .A2(_00797_ ), .A3(_06550_ ), .ZN(_01627_ ) );
NOR2_X1 _17812_ ( .A1(_01627_ ), .A2(_01599_ ), .ZN(_01628_ ) );
OAI21_X1 _17813_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01628_ ), .ZN(_01629_ ) );
OAI21_X1 _17814_ ( .A(_01629_ ), .B1(_01603_ ), .B2(_01614_ ), .ZN(_01630_ ) );
MUX2_X1 _17815_ ( .A(\EX_LS_result_reg [18] ), .B(_01630_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _17816_ ( .A1(_00798_ ), .A2(_00800_ ), .A3(_06550_ ), .ZN(_01631_ ) );
NOR2_X1 _17817_ ( .A1(_01631_ ), .A2(_01599_ ), .ZN(_01632_ ) );
OAI21_X1 _17818_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01632_ ), .ZN(_01633_ ) );
OAI21_X1 _17819_ ( .A(_01633_ ), .B1(_01603_ ), .B2(_01614_ ), .ZN(_01634_ ) );
MUX2_X1 _17820_ ( .A(\EX_LS_result_reg [17] ), .B(_01634_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _17821_ ( .A1(_00801_ ), .A2(_00803_ ), .A3(_02270_ ), .ZN(_01635_ ) );
NOR2_X1 _17822_ ( .A1(_01635_ ), .A2(_01599_ ), .ZN(_01636_ ) );
OAI21_X1 _17823_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01636_ ), .ZN(_01637_ ) );
OAI21_X1 _17824_ ( .A(_01637_ ), .B1(_01603_ ), .B2(_01614_ ), .ZN(_01638_ ) );
MUX2_X1 _17825_ ( .A(\EX_LS_result_reg [16] ), .B(_01638_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
INV_X1 _17826_ ( .A(_01585_ ), .ZN(_01639_ ) );
AOI21_X1 _17827_ ( .A(_01639_ ), .B1(_01582_ ), .B2(_01583_ ), .ZN(_01640_ ) );
OR3_X1 _17828_ ( .A1(_01591_ ), .A2(_01585_ ), .A3(_01593_ ), .ZN(_01641_ ) );
NOR3_X1 _17829_ ( .A1(_00807_ ), .A2(_06506_ ), .A3(_01641_ ), .ZN(_01642_ ) );
NOR2_X1 _17830_ ( .A1(_01640_ ), .A2(_01642_ ), .ZN(_01643_ ) );
AOI22_X1 _17831_ ( .A1(_01622_ ), .A2(_01643_ ), .B1(_01626_ ), .B2(_04151_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
NOR2_X1 _17832_ ( .A1(_01639_ ), .A2(_01580_ ), .ZN(_01644_ ) );
NOR2_X1 _17833_ ( .A1(_05676_ ), .A2(_01644_ ), .ZN(_01645_ ) );
INV_X1 _17834_ ( .A(_01594_ ), .ZN(_01646_ ) );
AND2_X1 _17835_ ( .A1(_01645_ ), .A2(_01646_ ), .ZN(_01647_ ) );
NAND3_X1 _17836_ ( .A1(_00808_ ), .A2(_00811_ ), .A3(_01647_ ), .ZN(_01648_ ) );
NOR2_X1 _17837_ ( .A1(_00783_ ), .A2(_06506_ ), .ZN(_01649_ ) );
NAND2_X1 _17838_ ( .A1(_01649_ ), .A2(_01644_ ), .ZN(_01650_ ) );
OAI211_X1 _17839_ ( .A(_01648_ ), .B(_01650_ ), .C1(_01614_ ), .C2(_01602_ ), .ZN(_01651_ ) );
MUX2_X1 _17840_ ( .A(\EX_LS_result_reg [14] ), .B(_01651_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
AND4_X1 _17841_ ( .A1(_06550_ ), .A2(_00820_ ), .A3(_00822_ ), .A4(_01644_ ), .ZN(_01652_ ) );
AND3_X1 _17842_ ( .A1(_00812_ ), .A2(_00816_ ), .A3(_01645_ ), .ZN(_01653_ ) );
OAI21_X1 _17843_ ( .A(_01646_ ), .B1(_01652_ ), .B2(_01653_ ), .ZN(_01654_ ) );
OAI21_X1 _17844_ ( .A(_01654_ ), .B1(_01614_ ), .B2(_01602_ ), .ZN(_01655_ ) );
MUX2_X1 _17845_ ( .A(\EX_LS_result_reg [13] ), .B(_01655_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
AND4_X1 _17846_ ( .A1(_06550_ ), .A2(_00854_ ), .A3(_00856_ ), .A4(_01644_ ), .ZN(_01656_ ) );
AND3_X1 _17847_ ( .A1(_00817_ ), .A2(_00819_ ), .A3(_01645_ ), .ZN(_01657_ ) );
OAI21_X1 _17848_ ( .A(_01646_ ), .B1(_01656_ ), .B2(_01657_ ), .ZN(_01658_ ) );
OAI21_X1 _17849_ ( .A(_01658_ ), .B1(_01614_ ), .B2(_01602_ ), .ZN(_01659_ ) );
MUX2_X1 _17850_ ( .A(\EX_LS_result_reg [12] ), .B(_01659_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
NOR3_X1 _17851_ ( .A1(_00783_ ), .A2(_06506_ ), .A3(_01599_ ), .ZN(_01660_ ) );
OAI21_X1 _17852_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01660_ ), .ZN(_01661_ ) );
OAI21_X1 _17853_ ( .A(_01661_ ), .B1(_01603_ ), .B2(_01613_ ), .ZN(_01662_ ) );
MUX2_X1 _17854_ ( .A(\EX_LS_result_reg [30] ), .B(_01662_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NAND4_X1 _17855_ ( .A1(_00863_ ), .A2(_00865_ ), .A3(\io_master_arid [1] ), .A4(_01644_ ), .ZN(_01663_ ) );
NAND3_X1 _17856_ ( .A1(_00823_ ), .A2(_00825_ ), .A3(_01647_ ), .ZN(_01664_ ) );
AND2_X1 _17857_ ( .A1(_01663_ ), .A2(_01664_ ), .ZN(_01665_ ) );
AOI22_X1 _17858_ ( .A1(_01622_ ), .A2(_01665_ ), .B1(_01626_ ), .B2(_04245_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
NAND3_X1 _17859_ ( .A1(_00826_ ), .A2(_00828_ ), .A3(_01647_ ), .ZN(_01666_ ) );
NAND4_X1 _17860_ ( .A1(_00866_ ), .A2(_00868_ ), .A3(_06550_ ), .A4(_01644_ ), .ZN(_01667_ ) );
OAI211_X1 _17861_ ( .A(_01666_ ), .B(_01667_ ), .C1(_01614_ ), .C2(_01602_ ), .ZN(_01668_ ) );
MUX2_X1 _17862_ ( .A(\EX_LS_result_reg [10] ), .B(_01668_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
NAND4_X1 _17863_ ( .A1(_00869_ ), .A2(_00871_ ), .A3(\io_master_arid [1] ), .A4(_01644_ ), .ZN(_01669_ ) );
NAND3_X1 _17864_ ( .A1(_00829_ ), .A2(_00831_ ), .A3(_01647_ ), .ZN(_01670_ ) );
AND2_X1 _17865_ ( .A1(_01669_ ), .A2(_01670_ ), .ZN(_01671_ ) );
AOI22_X1 _17866_ ( .A1(_01622_ ), .A2(_01671_ ), .B1(_01626_ ), .B2(_04294_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _17867_ ( .A1(_00833_ ), .A2(_00835_ ), .A3(_01647_ ), .ZN(_01672_ ) );
NAND4_X1 _17868_ ( .A1(_00872_ ), .A2(_00874_ ), .A3(_06550_ ), .A4(_01644_ ), .ZN(_01673_ ) );
OAI211_X1 _17869_ ( .A(_01672_ ), .B(_01673_ ), .C1(_01614_ ), .C2(_01602_ ), .ZN(_01674_ ) );
MUX2_X1 _17870_ ( .A(\EX_LS_result_reg [8] ), .B(_01674_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
OR3_X4 _17871_ ( .A1(_01612_ ), .A2(\mylsu.typ_tmp [2] ), .A3(_01592_ ), .ZN(_01675_ ) );
MUX2_X1 _17872_ ( .A(_01606_ ), .B(_01608_ ), .S(_01644_ ), .Z(_01676_ ) );
OAI21_X1 _17873_ ( .A(_01676_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01592_ ), .ZN(_01677_ ) );
AOI21_X2 _17874_ ( .A(_01591_ ), .B1(_01675_ ), .B2(_01677_ ), .ZN(_01678_ ) );
OR2_X2 _17875_ ( .A1(_01678_ ), .A2(_01621_ ), .ZN(_01679_ ) );
MUX2_X2 _17876_ ( .A(\EX_LS_result_reg [7] ), .B(_01679_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
AND2_X2 _17877_ ( .A1(_01594_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01680_ ) );
NAND2_X1 _17878_ ( .A1(_01641_ ), .A2(_01581_ ), .ZN(_01681_ ) );
NOR2_X1 _17879_ ( .A1(_01680_ ), .A2(_01681_ ), .ZN(_01682_ ) );
AOI221_X4 _17880_ ( .A(_06432_ ), .B1(_01443_ ), .B2(_01682_ ), .C1(_00841_ ), .C2(_01681_ ), .ZN(_01683_ ) );
NOR2_X1 _17881_ ( .A1(_00783_ ), .A2(_06508_ ), .ZN(_01684_ ) );
OAI21_X1 _17882_ ( .A(_01680_ ), .B1(_01111_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01685_ ) );
OAI211_X1 _17883_ ( .A(_01683_ ), .B(\io_master_arid [1] ), .C1(_01684_ ), .C2(_01685_ ), .ZN(_01686_ ) );
NAND2_X1 _17884_ ( .A1(_01626_ ), .A2(\EX_LS_result_reg [6] ), .ZN(_01687_ ) );
NAND2_X1 _17885_ ( .A1(_01686_ ), .A2(_01687_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
AOI221_X4 _17886_ ( .A(_06432_ ), .B1(_00993_ ), .B2(_01682_ ), .C1(_00844_ ), .C2(_01681_ ), .ZN(_01688_ ) );
AND3_X1 _17887_ ( .A1(_00820_ ), .A2(_00822_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01689_ ) );
OAI21_X1 _17888_ ( .A(_01680_ ), .B1(_01128_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01690_ ) );
OAI211_X1 _17889_ ( .A(_01688_ ), .B(\io_master_arid [1] ), .C1(_01689_ ), .C2(_01690_ ), .ZN(_01691_ ) );
NAND2_X1 _17890_ ( .A1(_01626_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01692_ ) );
NAND2_X1 _17891_ ( .A1(_01691_ ), .A2(_01692_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
AOI221_X4 _17892_ ( .A(_06432_ ), .B1(_01012_ ), .B2(_01682_ ), .C1(_00847_ ), .C2(_01681_ ), .ZN(_01693_ ) );
AND3_X1 _17893_ ( .A1(_00854_ ), .A2(_00856_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01694_ ) );
OAI21_X1 _17894_ ( .A(_01680_ ), .B1(_01145_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01695_ ) );
OAI211_X1 _17895_ ( .A(_01693_ ), .B(\io_master_arid [1] ), .C1(_01694_ ), .C2(_01695_ ), .ZN(_01696_ ) );
NAND2_X1 _17896_ ( .A1(_01626_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_01697_ ) );
NAND2_X1 _17897_ ( .A1(_01696_ ), .A2(_01697_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
AOI221_X4 _17898_ ( .A(_06432_ ), .B1(_01030_ ), .B2(_01682_ ), .C1(_00850_ ), .C2(_01681_ ), .ZN(_01698_ ) );
AND3_X1 _17899_ ( .A1(_00863_ ), .A2(_00865_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01699_ ) );
OAI21_X1 _17900_ ( .A(_01680_ ), .B1(_01179_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01700_ ) );
OAI211_X1 _17901_ ( .A(_01698_ ), .B(\io_master_arid [1] ), .C1(_01699_ ), .C2(_01700_ ), .ZN(_01701_ ) );
NAND2_X1 _17902_ ( .A1(_01626_ ), .A2(\EX_LS_result_reg [3] ), .ZN(_01702_ ) );
NAND2_X1 _17903_ ( .A1(_01701_ ), .A2(_01702_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
AOI221_X4 _17904_ ( .A(_06431_ ), .B1(_01047_ ), .B2(_01682_ ), .C1(_00853_ ), .C2(_01681_ ), .ZN(_01703_ ) );
AND3_X1 _17905_ ( .A1(_00866_ ), .A2(_00868_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01704_ ) );
OAI21_X1 _17906_ ( .A(_01680_ ), .B1(_01195_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01705_ ) );
OAI211_X1 _17907_ ( .A(_01703_ ), .B(\io_master_arid [1] ), .C1(_01704_ ), .C2(_01705_ ), .ZN(_01706_ ) );
NAND2_X1 _17908_ ( .A1(_06432_ ), .A2(\EX_LS_result_reg [2] ), .ZN(_01707_ ) );
NAND2_X1 _17909_ ( .A1(_01706_ ), .A2(_01707_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
NOR3_X1 _17910_ ( .A1(_01161_ ), .A2(_06506_ ), .A3(_01599_ ), .ZN(_01708_ ) );
OAI21_X1 _17911_ ( .A(_01595_ ), .B1(_01616_ ), .B2(_01708_ ), .ZN(_01709_ ) );
OAI21_X1 _17912_ ( .A(_01709_ ), .B1(_01603_ ), .B2(_01613_ ), .ZN(_01710_ ) );
MUX2_X1 _17913_ ( .A(\EX_LS_result_reg [29] ), .B(_01710_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
AOI221_X4 _17914_ ( .A(_06431_ ), .B1(_01062_ ), .B2(_01682_ ), .C1(_00859_ ), .C2(_01681_ ), .ZN(_01711_ ) );
AND3_X1 _17915_ ( .A1(_00869_ ), .A2(_00871_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01712_ ) );
OAI21_X1 _17916_ ( .A(_01680_ ), .B1(_01211_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01713_ ) );
OAI211_X1 _17917_ ( .A(_01711_ ), .B(\io_master_arid [1] ), .C1(_01712_ ), .C2(_01713_ ), .ZN(_01714_ ) );
NAND2_X1 _17918_ ( .A1(_06432_ ), .A2(\EX_LS_result_reg [1] ), .ZN(_01715_ ) );
NAND2_X1 _17919_ ( .A1(_01714_ ), .A2(_01715_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
AOI221_X4 _17920_ ( .A(_06431_ ), .B1(_01079_ ), .B2(_01682_ ), .C1(_00862_ ), .C2(_01681_ ), .ZN(_01716_ ) );
AND3_X1 _17921_ ( .A1(_00872_ ), .A2(_00874_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01717_ ) );
OAI21_X1 _17922_ ( .A(_01680_ ), .B1(_00920_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01718_ ) );
OAI211_X1 _17923_ ( .A(_01716_ ), .B(\io_master_arid [1] ), .C1(_01717_ ), .C2(_01718_ ), .ZN(_01719_ ) );
OAI21_X1 _17924_ ( .A(_01719_ ), .B1(\mylsu.state [3] ), .B2(_04079_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
NOR3_X1 _17925_ ( .A1(_01335_ ), .A2(_06506_ ), .A3(_01598_ ), .ZN(_01720_ ) );
OAI21_X1 _17926_ ( .A(_01595_ ), .B1(_01616_ ), .B2(_01720_ ), .ZN(_01721_ ) );
OAI21_X1 _17927_ ( .A(_01721_ ), .B1(_01603_ ), .B2(_01613_ ), .ZN(_01722_ ) );
MUX2_X1 _17928_ ( .A(\EX_LS_result_reg [28] ), .B(_01722_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
NOR3_X1 _17929_ ( .A1(_01365_ ), .A2(_06506_ ), .A3(_01599_ ), .ZN(_01723_ ) );
OAI21_X1 _17930_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01723_ ), .ZN(_01724_ ) );
AOI22_X1 _17931_ ( .A1(_01622_ ), .A2(_01724_ ), .B1(_01626_ ), .B2(_03988_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
NOR3_X1 _17932_ ( .A1(_01381_ ), .A2(_06506_ ), .A3(_01598_ ), .ZN(_01725_ ) );
OAI21_X1 _17933_ ( .A(_01595_ ), .B1(_01587_ ), .B2(_01725_ ), .ZN(_01726_ ) );
OAI21_X1 _17934_ ( .A(_01726_ ), .B1(_01603_ ), .B2(_01613_ ), .ZN(_01727_ ) );
MUX2_X1 _17935_ ( .A(\EX_LS_result_reg [26] ), .B(_01727_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
NOR3_X1 _17936_ ( .A1(_01396_ ), .A2(_06506_ ), .A3(_01599_ ), .ZN(_01728_ ) );
OAI21_X1 _17937_ ( .A(_01596_ ), .B1(_01616_ ), .B2(_01728_ ), .ZN(_01729_ ) );
AOI22_X1 _17938_ ( .A1(_01622_ ), .A2(_01729_ ), .B1(_01626_ ), .B2(_03963_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
NOR3_X1 _17939_ ( .A1(_01412_ ), .A2(_06506_ ), .A3(_01598_ ), .ZN(_01730_ ) );
OAI21_X1 _17940_ ( .A(_01595_ ), .B1(_01587_ ), .B2(_01730_ ), .ZN(_01731_ ) );
OAI21_X1 _17941_ ( .A(_01731_ ), .B1(_01603_ ), .B2(_01613_ ), .ZN(_01732_ ) );
MUX2_X1 _17942_ ( .A(\EX_LS_result_reg [24] ), .B(_01732_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _17943_ ( .A1(_00877_ ), .A2(_05676_ ), .A3(_01598_ ), .ZN(_01733_ ) );
OAI21_X1 _17944_ ( .A(_01595_ ), .B1(_01587_ ), .B2(_01733_ ), .ZN(_01734_ ) );
OAI21_X1 _17945_ ( .A(_01734_ ), .B1(_01602_ ), .B2(_01613_ ), .ZN(_01735_ ) );
MUX2_X1 _17946_ ( .A(\EX_LS_result_reg [23] ), .B(_01735_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _17947_ ( .A1(_01443_ ), .A2(_05676_ ), .A3(_01598_ ), .ZN(_01736_ ) );
OAI21_X1 _17948_ ( .A(_01595_ ), .B1(_01587_ ), .B2(_01736_ ), .ZN(_01737_ ) );
OAI21_X1 _17949_ ( .A(_01737_ ), .B1(_01602_ ), .B2(_01613_ ), .ZN(_01738_ ) );
MUX2_X1 _17950_ ( .A(\EX_LS_result_reg [22] ), .B(_01738_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _17951_ ( .A(_01586_ ), .B(_01610_ ), .S(_01639_ ), .Z(_01739_ ) );
NAND2_X1 _17952_ ( .A1(_01596_ ), .A2(_01739_ ), .ZN(_01740_ ) );
OAI21_X1 _17953_ ( .A(_01740_ ), .B1(_01602_ ), .B2(_01613_ ), .ZN(_01741_ ) );
MUX2_X1 _17954_ ( .A(\EX_LS_result_reg [31] ), .B(_01741_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17955_ ( .A1(\LS_WB_waddr_reg [1] ), .A2(\LS_WB_waddr_reg [0] ), .ZN(_01742_ ) );
INV_X1 _17956_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01743_ ) );
INV_X1 _17957_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01744_ ) );
NAND3_X1 _17958_ ( .A1(_01742_ ), .A2(_01743_ ), .A3(_01744_ ), .ZN(_01745_ ) );
AND2_X1 _17959_ ( .A1(_01773_ ), .A2(LS_WB_wen_reg ), .ZN(_01746_ ) );
NAND2_X1 _17960_ ( .A1(_01745_ ), .A2(_01746_ ), .ZN(_01747_ ) );
BUF_X4 _17961_ ( .A(_01747_ ), .Z(_01748_ ) );
AOI21_X1 _17962_ ( .A(_01748_ ), .B1(_01743_ ), .B2(_01744_ ), .ZN(_01749_ ) );
INV_X1 _17963_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01750_ ) );
INV_X1 _17964_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01751_ ) );
NOR4_X1 _17965_ ( .A1(_01749_ ), .A2(_01750_ ), .A3(_01751_ ), .A4(_01748_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
AOI21_X1 _17966_ ( .A(_01748_ ), .B1(_01750_ ), .B2(_01751_ ), .ZN(_01752_ ) );
NOR2_X1 _17967_ ( .A1(_01747_ ), .A2(_01743_ ), .ZN(_01753_ ) );
NOR4_X1 _17968_ ( .A1(_01752_ ), .A2(_01753_ ), .A3(_01744_ ), .A4(_01748_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
NOR2_X1 _17969_ ( .A1(_01748_ ), .A2(_01744_ ), .ZN(_01754_ ) );
NOR4_X1 _17970_ ( .A1(_01752_ ), .A2(_01754_ ), .A3(_01743_ ), .A4(_01748_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR2_X1 _17971_ ( .A1(_01748_ ), .A2(_01750_ ), .ZN(_01755_ ) );
AND4_X1 _17972_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01755_ ), .A3(_01753_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
NOR2_X1 _17973_ ( .A1(_01747_ ), .A2(_01751_ ), .ZN(_01756_ ) );
AND4_X1 _17974_ ( .A1(_01744_ ), .A2(_01756_ ), .A3(_01753_ ), .A4(_01750_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
CLKBUF_X1 _17975_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17976_ ( .A1(_01749_ ), .A2(_01755_ ), .A3(_01751_ ), .A4(_01748_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17977_ ( .A1(_01743_ ), .A2(_01756_ ), .A3(_01754_ ), .A4(_01750_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17978_ ( .A1(_01743_ ), .A2(_01755_ ), .A3(_01754_ ), .A4(_01751_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
AND4_X1 _17979_ ( .A1(_01743_ ), .A2(_01756_ ), .A3(_01754_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17980_ ( .A1(_01744_ ), .A2(_01756_ ), .A3(_01753_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
NOR4_X1 _17981_ ( .A1(_01752_ ), .A2(_01743_ ), .A3(_01744_ ), .A4(_01748_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17982_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01756_ ), .A3(_01753_ ), .A4(_01750_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17983_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01755_ ), .A3(_01753_ ), .A4(_01751_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17984_ ( .A1(_01744_ ), .A2(_01755_ ), .A3(_01753_ ), .A4(_01751_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17985_ ( .A1(_01749_ ), .A2(_01756_ ), .A3(_01750_ ), .A4(_01748_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17986_ ( .A1(_02249_ ), .A2(_03400_ ), .A3(_02257_ ), .ZN(_01757_ ) );
NAND2_X1 _17987_ ( .A1(_01757_ ), .A2(_03400_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17988_ ( .A(reset ), .B(_02249_ ), .C1(_02250_ ), .C2(_02277_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17989_ ( .A(_01745_ ), .Z(_01758_ ) );
CLKBUF_X2 _17990_ ( .A(_01746_ ), .Z(_01759_ ) );
AND3_X1 _17991_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17992_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17993_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17994_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17995_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17996_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17997_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17998_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17999_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _18000_ ( .A1(_01758_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01759_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _18001_ ( .A(_01745_ ), .Z(_01760_ ) );
CLKBUF_X2 _18002_ ( .A(_01746_ ), .Z(_01761_ ) );
AND3_X1 _18003_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _18004_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _18005_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _18006_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _18007_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _18008_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _18009_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _18010_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _18011_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _18012_ ( .A1(_01760_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01761_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _18013_ ( .A(_01745_ ), .Z(_01762_ ) );
CLKBUF_X2 _18014_ ( .A(_01746_ ), .Z(_01763_ ) );
AND3_X1 _18015_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _18016_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _18017_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _18018_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _18019_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _18020_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _18021_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _18022_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _18023_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _18024_ ( .A1(_01762_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01763_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _18025_ ( .A1(_01745_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01746_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _18026_ ( .A1(_01745_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01746_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_D ) );
AND3_X1 _18027_ ( .A1(_01914_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _18028_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01764_ ) );
AND2_X1 _18029_ ( .A1(_01764_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01765_ ) );
INV_X1 _18030_ ( .A(_01765_ ), .ZN(_01766_ ) );
NOR2_X1 _18031_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01767_ ) );
OAI211_X1 _18032_ ( .A(_01773_ ), .B(\mysc.state [0] ), .C1(_01766_ ), .C2(_01767_ ), .ZN(_01768_ ) );
INV_X1 _18033_ ( .A(_01768_ ), .ZN(_01769_ ) );
OR3_X1 _18034_ ( .A1(_01769_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _18035_ ( .A1(_01766_ ), .A2(reset ), .A3(_01767_ ), .ZN(_01770_ ) );
NAND2_X1 _18036_ ( .A1(_01770_ ), .A2(\mysc.state [0] ), .ZN(_01771_ ) );
OR3_X1 _18037_ ( .A1(_06501_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01772_ ) );
NAND2_X1 _18038_ ( .A1(_01771_ ), .A2(_01772_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _18039_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_08254_ ) );
CLKGATE_X1 _18040_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_08255_ ) );
CLKGATE_X1 _18041_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_08256_ ) );
CLKGATE_X1 _18042_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08257_ ) );
CLKGATE_X1 _18043_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08258_ ) );
CLKGATE_X1 _18044_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08259_ ) );
CLKGATE_X1 _18045_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08260_ ) );
CLKGATE_X1 _18046_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_08261_ ) );
CLKGATE_X1 _18047_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_08262_ ) );
CLKGATE_X1 _18048_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_08263_ ) );
CLKGATE_X1 _18049_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_08264_ ) );
CLKGATE_X1 _18050_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_08265_ ) );
CLKGATE_X1 _18051_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08266_ ) );
CLKGATE_X1 _18052_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08267_ ) );
CLKGATE_X1 _18053_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08268_ ) );
CLKGATE_X1 _18054_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_08269_ ) );
CLKGATE_X1 _18055_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_08270_ ) );
CLKGATE_X1 _18056_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08271_ ) );
CLKGATE_X1 _18057_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_08272_ ) );
CLKGATE_X1 _18058_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ), .GCK(_08273_ ) );
CLKGATE_X1 _18059_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .GCK(_08274_ ) );
CLKGATE_X1 _18060_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08275_ ) );
CLKGATE_X1 _18061_ ( .CK(clock ), .E(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_08276_ ) );
CLKGATE_X1 _18062_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_08277_ ) );
CLKGATE_X1 _18063_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_08278_ ) );
CLKGATE_X1 _18064_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_08279_ ) );
CLKGATE_X1 _18065_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_08280_ ) );
CLKGATE_X1 _18066_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_08281_ ) );
CLKGATE_X1 _18067_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_08282_ ) );
CLKGATE_X1 _18068_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_08283_ ) );
CLKGATE_X1 _18069_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_08284_ ) );
CLKGATE_X1 _18070_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_08285_ ) );
CLKGATE_X1 _18071_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_08286_ ) );
CLKGATE_X1 _18072_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_08287_ ) );
CLKGATE_X1 _18073_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_08288_ ) );
CLKGATE_X1 _18074_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08289_ ) );
CLKGATE_X1 _18075_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08290_ ) );
CLKGATE_X1 _18076_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08291_ ) );
CLKGATE_X1 _18077_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08292_ ) );
CLKGATE_X1 _18078_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08293_ ) );
CLKGATE_X1 _18079_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08294_ ) );
CLKGATE_X1 _18080_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08295_ ) );
CLKGATE_X1 _18081_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08296_ ) );
CLKGATE_X1 _18082_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08297_ ) );
CLKGATE_X1 _18083_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08298_ ) );
CLKGATE_X1 _18084_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_08299_ ) );
CLKGATE_X1 _18085_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08300_ ) );
CLKGATE_X1 _18086_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08301_ ) );
CLKGATE_X1 _18087_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08302_ ) );
CLKGATE_X1 _18088_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08303_ ) );
CLKGATE_X1 _18089_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08304_ ) );
CLKGATE_X1 _18090_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_08305_ ) );
CLKGATE_X1 _18091_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08306_ ) );
CLKGATE_X1 _18092_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08307_ ) );
CLKGATE_X1 _18093_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08308_ ) );
CLKGATE_X1 _18094_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08309_ ) );
CLKGATE_X1 _18095_ ( .CK(clock ), .E(\myexu.pc_out_$_SDFFE_PP0P__Q_E ), .GCK(_08310_ ) );
CLKGATE_X1 _18096_ ( .CK(clock ), .E(\myidu.state_$_ANDNOT__A_Y ), .GCK(_08311_ ) );
CLKGATE_X1 _18097_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08312_ ) );
CLKGATE_X1 _18098_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08313_ ) );
CLKGATE_X1 _18099_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08314_ ) );
CLKGATE_X1 _18100_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ), .GCK(_08315_ ) );
CLKGATE_X1 _18101_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ), .GCK(_08316_ ) );
CLKGATE_X1 _18102_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08317_ ) );
LOGIC1_X1 _18103_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _18104_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08548_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08549_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08550_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08551_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08552_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08553_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08554_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08555_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08556_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08557_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08558_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08559_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08560_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08561_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08562_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08563_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08564_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08565_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08566_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08567_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08568_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08569_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08570_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08571_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08572_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08573_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08574_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08575_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08576_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08577_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08578_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08317_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08579_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08316_ ), .Q(\mtvec [31] ), .QN(_08580_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08316_ ), .Q(\mtvec [30] ), .QN(_08581_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08316_ ), .Q(\mtvec [21] ), .QN(_08582_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08316_ ), .Q(\mtvec [20] ), .QN(_08583_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08316_ ), .Q(\mtvec [19] ), .QN(_08584_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08316_ ), .Q(\mtvec [18] ), .QN(_08585_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08316_ ), .Q(\mtvec [17] ), .QN(_08586_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08316_ ), .Q(\mtvec [16] ), .QN(_08587_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08316_ ), .Q(\mtvec [15] ), .QN(_08588_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08316_ ), .Q(\mtvec [14] ), .QN(_08589_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08316_ ), .Q(\mtvec [13] ), .QN(_08590_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08316_ ), .Q(\mtvec [12] ), .QN(_08591_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08316_ ), .Q(\mtvec [29] ), .QN(_08592_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08316_ ), .Q(\mtvec [11] ), .QN(_08593_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08316_ ), .Q(\mtvec [10] ), .QN(_08594_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08316_ ), .Q(\mtvec [9] ), .QN(_08595_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08316_ ), .Q(\mtvec [8] ), .QN(_08596_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08316_ ), .Q(\mtvec [7] ), .QN(_08597_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08316_ ), .Q(\mtvec [6] ), .QN(_08598_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08316_ ), .Q(\mtvec [5] ), .QN(_08599_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08316_ ), .Q(\mtvec [4] ), .QN(_08600_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08316_ ), .Q(\mtvec [3] ), .QN(_08601_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08316_ ), .Q(\mtvec [2] ), .QN(_08602_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08316_ ), .Q(\mtvec [28] ), .QN(_08603_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08316_ ), .Q(\mtvec [1] ), .QN(_08604_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08316_ ), .Q(\mtvec [0] ), .QN(_08605_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08316_ ), .Q(\mtvec [27] ), .QN(_08606_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08316_ ), .Q(\mtvec [26] ), .QN(_08607_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08316_ ), .Q(\mtvec [25] ), .QN(_08608_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08316_ ), .Q(\mtvec [24] ), .QN(_08609_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08316_ ), .Q(\mtvec [23] ), .QN(_08610_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08316_ ), .Q(\mtvec [22] ), .QN(_08611_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08315_ ), .Q(\mepc [31] ), .QN(_08612_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08315_ ), .Q(\mepc [30] ), .QN(_08613_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08315_ ), .Q(\mepc [21] ), .QN(_08614_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08315_ ), .Q(\mepc [20] ), .QN(_08615_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08315_ ), .Q(\mepc [19] ), .QN(_08616_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08315_ ), .Q(\mepc [18] ), .QN(_08617_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08315_ ), .Q(\mepc [17] ), .QN(_08618_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08315_ ), .Q(\mepc [16] ), .QN(_08619_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08315_ ), .Q(\mepc [15] ), .QN(_08620_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08315_ ), .Q(\mepc [14] ), .QN(_08621_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08315_ ), .Q(\mepc [13] ), .QN(_08622_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08315_ ), .Q(\mepc [12] ), .QN(_08623_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08315_ ), .Q(\mepc [29] ), .QN(_08624_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08315_ ), .Q(\mepc [11] ), .QN(_08625_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08315_ ), .Q(\mepc [10] ), .QN(_08626_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08315_ ), .Q(\mepc [9] ), .QN(_08627_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08315_ ), .Q(\mepc [8] ), .QN(_08628_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08315_ ), .Q(\mepc [7] ), .QN(_08629_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08315_ ), .Q(\mepc [6] ), .QN(_08630_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08315_ ), .Q(\mepc [5] ), .QN(_08631_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08315_ ), .Q(\mepc [4] ), .QN(_08632_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08315_ ), .Q(\mepc [3] ), .QN(_08633_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08315_ ), .Q(\mepc [2] ), .QN(_08634_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08315_ ), .Q(\mepc [28] ), .QN(_08635_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08315_ ), .Q(\mepc [1] ), .QN(_08636_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08315_ ), .Q(\mepc [0] ), .QN(_08637_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08315_ ), .Q(\mepc [27] ), .QN(_08638_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08315_ ), .Q(\mepc [26] ), .QN(_08639_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08315_ ), .Q(\mepc [25] ), .QN(_08640_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08315_ ), .Q(\mepc [24] ), .QN(_08641_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08315_ ), .Q(\mepc [23] ), .QN(_08642_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08315_ ), .Q(\mepc [22] ), .QN(_08643_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08644_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08645_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08646_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08547_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08546_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08545_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08544_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08543_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08542_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08541_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08540_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08539_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08538_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08537_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08536_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08535_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08534_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08533_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08532_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08531_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08530_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08529_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08528_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08527_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08526_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00086_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08525_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00087_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08524_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00088_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08523_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00089_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08522_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00090_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08521_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00091_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08520_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00092_ ), .CK(_08314_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08647_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PN0__Q ( .D(_00093_ ), .CK(clock ), .Q(excp_written ), .QN(_08648_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08519_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08649_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08650_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08651_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08652_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08653_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08654_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08655_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08656_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08657_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08658_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08659_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08660_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08661_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08662_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08663_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08664_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08665_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08666_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08667_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08668_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08669_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08670_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08671_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08672_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08673_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08674_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08675_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08676_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08677_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08678_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08313_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08518_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00094_ ), .CK(_08312_ ), .Q(\myec.state [1] ), .QN(_08517_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00095_ ), .CK(_08312_ ), .Q(\myec.state [0] ), .QN(_08679_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PP0__Q ( .D(_00096_ ), .CK(clock ), .Q(check_quest ), .QN(_08680_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08516_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08681_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08682_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08683_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08684_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08685_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08686_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08687_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08688_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08689_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08690_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08515_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00097_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08514_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00098_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08513_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00099_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08512_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00100_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08511_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00101_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08510_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00102_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08509_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00103_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08508_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00104_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08507_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00105_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08506_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00106_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08505_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00107_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08504_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00108_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08503_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00109_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08502_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00110_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08501_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00111_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08500_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00112_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08499_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00113_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08498_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00114_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08497_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00115_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08496_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00116_ ), .CK(_08311_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08495_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q ( .D(_00117_ ), .CK(_08310_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08494_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_1 ( .D(_00118_ ), .CK(_08310_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08493_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_2 ( .D(_00119_ ), .CK(_08310_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08492_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_3 ( .D(_00120_ ), .CK(_08310_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08491_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_4 ( .D(_00121_ ), .CK(_08310_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08490_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q ( .D(_00123_ ), .CK(clock ), .Q(\myexu.pc_jump [30] ), .QN(_08488_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_1 ( .D(_00124_ ), .CK(clock ), .Q(\myexu.pc_jump [29] ), .QN(_08487_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_10 ( .D(_00125_ ), .CK(clock ), .Q(\myexu.pc_jump [20] ), .QN(_08486_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_11 ( .D(_00126_ ), .CK(clock ), .Q(\myexu.pc_jump [19] ), .QN(_08485_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_12 ( .D(_00127_ ), .CK(clock ), .Q(\myexu.pc_jump [18] ), .QN(_08484_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_13 ( .D(_00128_ ), .CK(clock ), .Q(\myexu.pc_jump [17] ), .QN(_08483_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_14 ( .D(_00129_ ), .CK(clock ), .Q(\myexu.pc_jump [16] ), .QN(_08482_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_15 ( .D(_00130_ ), .CK(clock ), .Q(\myexu.pc_jump [15] ), .QN(_08481_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_16 ( .D(_00131_ ), .CK(clock ), .Q(\myexu.pc_jump [14] ), .QN(_08480_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_17 ( .D(_00132_ ), .CK(clock ), .Q(\myexu.pc_jump [13] ), .QN(_08479_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_18 ( .D(_00133_ ), .CK(clock ), .Q(\myexu.pc_jump [12] ), .QN(_08478_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_19 ( .D(_00134_ ), .CK(clock ), .Q(\myexu.pc_jump [11] ), .QN(_08477_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_2 ( .D(_00135_ ), .CK(clock ), .Q(\myexu.pc_jump [28] ), .QN(_08476_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_20 ( .D(_00136_ ), .CK(clock ), .Q(\myexu.pc_jump [10] ), .QN(_08475_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_21 ( .D(_00137_ ), .CK(clock ), .Q(\myexu.pc_jump [9] ), .QN(_08474_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_22 ( .D(_00138_ ), .CK(clock ), .Q(\myexu.pc_jump [8] ), .QN(_08473_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_23 ( .D(_00139_ ), .CK(clock ), .Q(\myexu.pc_jump [7] ), .QN(_08472_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_24 ( .D(_00140_ ), .CK(clock ), .Q(\myexu.pc_jump [6] ), .QN(_08471_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_25 ( .D(_00141_ ), .CK(clock ), .Q(\myexu.pc_jump [5] ), .QN(_08470_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_26 ( .D(_00142_ ), .CK(clock ), .Q(\myexu.pc_jump [4] ), .QN(_08469_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_27 ( .D(_00143_ ), .CK(clock ), .Q(\myexu.pc_jump [3] ), .QN(_08468_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_28 ( .D(_00144_ ), .CK(clock ), .Q(\myexu.pc_jump [2] ), .QN(_08467_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_29 ( .D(_00145_ ), .CK(clock ), .Q(\myexu.pc_jump [1] ), .QN(_08466_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_3 ( .D(_00146_ ), .CK(clock ), .Q(\myexu.pc_jump [27] ), .QN(_08465_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_30 ( .D(_00147_ ), .CK(clock ), .Q(\myexu.pc_jump [0] ), .QN(_08464_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_4 ( .D(_00148_ ), .CK(clock ), .Q(\myexu.pc_jump [26] ), .QN(_08463_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_5 ( .D(_00149_ ), .CK(clock ), .Q(\myexu.pc_jump [25] ), .QN(_08462_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_6 ( .D(_00150_ ), .CK(clock ), .Q(\myexu.pc_jump [24] ), .QN(_08461_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_7 ( .D(_00151_ ), .CK(clock ), .Q(\myexu.pc_jump [23] ), .QN(_08460_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_8 ( .D(_00152_ ), .CK(clock ), .Q(\myexu.pc_jump [22] ), .QN(_08459_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP0__Q_9 ( .D(_00153_ ), .CK(clock ), .Q(\myexu.pc_jump [21] ), .QN(_08458_ ) );
DFF_X1 \myexu.pc_jump_$_SDFF_PP1__Q ( .D(_00154_ ), .CK(clock ), .Q(\myexu.pc_jump [31] ), .QN(_08457_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q ( .D(_00122_ ), .CK(_08310_ ), .Q(\EX_LS_pc [31] ), .QN(_08489_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_1 ( .D(_00155_ ), .CK(_08310_ ), .Q(\EX_LS_pc [30] ), .QN(_08456_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_10 ( .D(_00156_ ), .CK(_08310_ ), .Q(\EX_LS_pc [21] ), .QN(_08455_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_11 ( .D(_00157_ ), .CK(_08310_ ), .Q(\EX_LS_pc [20] ), .QN(_08454_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_12 ( .D(_00158_ ), .CK(_08310_ ), .Q(\EX_LS_pc [19] ), .QN(_08453_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_13 ( .D(_00159_ ), .CK(_08310_ ), .Q(\EX_LS_pc [18] ), .QN(_08452_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_14 ( .D(_00160_ ), .CK(_08310_ ), .Q(\EX_LS_pc [17] ), .QN(_08451_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_15 ( .D(_00161_ ), .CK(_08310_ ), .Q(\EX_LS_pc [16] ), .QN(_08450_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_16 ( .D(_00162_ ), .CK(_08310_ ), .Q(\EX_LS_pc [15] ), .QN(_08449_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_17 ( .D(_00163_ ), .CK(_08310_ ), .Q(\EX_LS_pc [14] ), .QN(_08448_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_18 ( .D(_00164_ ), .CK(_08310_ ), .Q(\EX_LS_pc [13] ), .QN(_08447_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_19 ( .D(_00165_ ), .CK(_08310_ ), .Q(\EX_LS_pc [12] ), .QN(_08446_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_2 ( .D(_00166_ ), .CK(_08310_ ), .Q(\EX_LS_pc [29] ), .QN(_08445_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_20 ( .D(_00167_ ), .CK(_08310_ ), .Q(\EX_LS_pc [11] ), .QN(_08444_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_21 ( .D(_00168_ ), .CK(_08310_ ), .Q(\EX_LS_pc [10] ), .QN(_08443_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_22 ( .D(_00169_ ), .CK(_08310_ ), .Q(\EX_LS_pc [9] ), .QN(_08442_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_23 ( .D(_00170_ ), .CK(_08310_ ), .Q(\EX_LS_pc [8] ), .QN(_08441_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_24 ( .D(_00171_ ), .CK(_08310_ ), .Q(\EX_LS_pc [7] ), .QN(_08440_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_25 ( .D(_00172_ ), .CK(_08310_ ), .Q(\EX_LS_pc [6] ), .QN(_08439_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_26 ( .D(_00173_ ), .CK(_08310_ ), .Q(\EX_LS_pc [5] ), .QN(_08438_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_27 ( .D(_00174_ ), .CK(_08310_ ), .Q(\EX_LS_pc [4] ), .QN(_08437_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_28 ( .D(_00175_ ), .CK(_08310_ ), .Q(\EX_LS_pc [3] ), .QN(_08436_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_29 ( .D(_00176_ ), .CK(_08310_ ), .Q(\EX_LS_pc [2] ), .QN(_08435_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_3 ( .D(_00177_ ), .CK(_08310_ ), .Q(\EX_LS_pc [28] ), .QN(_08434_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_30 ( .D(_00178_ ), .CK(_08310_ ), .Q(\EX_LS_pc [1] ), .QN(_08433_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_31 ( .D(_00179_ ), .CK(_08310_ ), .Q(\EX_LS_pc [0] ), .QN(_08432_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_4 ( .D(_00180_ ), .CK(_08310_ ), .Q(\EX_LS_pc [27] ), .QN(_08431_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_5 ( .D(_00181_ ), .CK(_08310_ ), .Q(\EX_LS_pc [26] ), .QN(_08430_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_6 ( .D(_00182_ ), .CK(_08310_ ), .Q(\EX_LS_pc [25] ), .QN(_08429_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_7 ( .D(_00183_ ), .CK(_08310_ ), .Q(\EX_LS_pc [24] ), .QN(_08428_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_8 ( .D(_00184_ ), .CK(_08310_ ), .Q(\EX_LS_pc [23] ), .QN(_08427_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_9 ( .D(_00185_ ), .CK(_08310_ ), .Q(\EX_LS_pc [22] ), .QN(_08691_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08692_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08693_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08694_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08695_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08696_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08697_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08698_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08699_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08700_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08701_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08702_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08703_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08704_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08705_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08706_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08707_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08708_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08709_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08710_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08711_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08712_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08713_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08714_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08715_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08716_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08717_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08718_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08719_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08720_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08721_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08722_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08311_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08723_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08311_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PP0__Q ( .D(_00187_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q ( .D(_00186_ ), .CK(_08310_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_1 ( .D(_00188_ ), .CK(_08310_ ), .Q(\EX_LS_flag [1] ), .QN(_08426_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_2 ( .D(_00189_ ), .CK(_08310_ ), .Q(\EX_LS_flag [0] ), .QN(_08425_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_3 ( .D(_00190_ ), .CK(_08310_ ), .Q(\EX_LS_typ [4] ), .QN(_08424_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_4 ( .D(_00191_ ), .CK(_08310_ ), .Q(\EX_LS_typ [3] ), .QN(_08423_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_5 ( .D(_00192_ ), .CK(_08310_ ), .Q(\EX_LS_typ [2] ), .QN(_08422_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_6 ( .D(_00193_ ), .CK(_08310_ ), .Q(\EX_LS_typ [1] ), .QN(_08421_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_7 ( .D(_00194_ ), .CK(_08310_ ), .Q(\EX_LS_typ [0] ), .QN(_08420_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00195_ ), .CK(_08309_ ), .Q(\ID_EX_csr [11] ), .QN(_08419_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00196_ ), .CK(_08309_ ), .Q(\ID_EX_csr [10] ), .QN(_08418_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00197_ ), .CK(_08309_ ), .Q(\ID_EX_csr [1] ), .QN(_08417_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00198_ ), .CK(_08309_ ), .Q(\ID_EX_csr [0] ), .QN(_08416_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00199_ ), .CK(_08309_ ), .Q(\ID_EX_csr [9] ), .QN(_08415_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00200_ ), .CK(_08309_ ), .Q(\ID_EX_csr [8] ), .QN(_08414_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00201_ ), .CK(_08309_ ), .Q(\ID_EX_csr [7] ), .QN(_08413_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00202_ ), .CK(_08309_ ), .Q(\ID_EX_csr [6] ), .QN(_08412_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00203_ ), .CK(_08309_ ), .Q(\ID_EX_csr [5] ), .QN(_08411_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00204_ ), .CK(_08309_ ), .Q(\ID_EX_csr [4] ), .QN(_08410_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00205_ ), .CK(_08309_ ), .Q(\ID_EX_csr [3] ), .QN(_08409_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00206_ ), .CK(_08309_ ), .Q(\ID_EX_csr [2] ), .QN(_08408_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00207_ ), .CK(_08308_ ), .Q(exception_quest_IDU ), .QN(_08407_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00208_ ), .CK(_08307_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08306_ ), .Q(\ID_EX_imm [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08306_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08306_ ), .Q(\ID_EX_imm [21] ), .QN(_08724_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08306_ ), .Q(\ID_EX_imm [20] ), .QN(_08725_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08306_ ), .Q(\ID_EX_imm [19] ), .QN(_08726_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08306_ ), .Q(\ID_EX_imm [18] ), .QN(_08727_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08306_ ), .Q(\ID_EX_imm [17] ), .QN(_08728_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08306_ ), .Q(\ID_EX_imm [16] ), .QN(_08729_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08306_ ), .Q(\ID_EX_imm [15] ), .QN(_08730_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08306_ ), .Q(\ID_EX_imm [14] ), .QN(_08731_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08306_ ), .Q(\ID_EX_imm [13] ), .QN(_08732_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08306_ ), .Q(\ID_EX_imm [12] ), .QN(_08733_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08306_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08306_ ), .Q(\ID_EX_imm [11] ), .QN(_08734_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08306_ ), .Q(\ID_EX_imm [10] ), .QN(_08735_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08306_ ), .Q(\ID_EX_imm [9] ), .QN(_08736_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08306_ ), .Q(\ID_EX_imm [8] ), .QN(_08737_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08306_ ), .Q(\ID_EX_imm [7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08306_ ), .Q(\ID_EX_imm [6] ), .QN(_08738_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08306_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08306_ ), .Q(\ID_EX_imm [4] ), .QN(_08739_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08306_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08306_ ), .Q(\ID_EX_imm [2] ), .QN(_08740_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08306_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08306_ ), .Q(\ID_EX_imm [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08306_ ), .Q(\ID_EX_imm [0] ), .QN(_08741_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08306_ ), .Q(\ID_EX_imm [27] ), .QN(_08742_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08306_ ), .Q(\ID_EX_imm [26] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08306_ ), .Q(\ID_EX_imm [25] ), .QN(_08743_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08306_ ), .Q(\ID_EX_imm [24] ), .QN(_08744_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08306_ ), .Q(\ID_EX_imm [23] ), .QN(_08745_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08306_ ), .Q(\ID_EX_imm [22] ), .QN(_08746_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08305_ ), .Q(\ID_EX_pc [31] ), .QN(_08747_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08305_ ), .Q(\ID_EX_pc [30] ), .QN(_08748_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08305_ ), .Q(\ID_EX_pc [21] ), .QN(_08749_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08305_ ), .Q(\ID_EX_pc [20] ), .QN(_08750_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08305_ ), .Q(\ID_EX_pc [19] ), .QN(_08751_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08305_ ), .Q(\ID_EX_pc [18] ), .QN(_08752_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08305_ ), .Q(\ID_EX_pc [17] ), .QN(_08753_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08305_ ), .Q(\ID_EX_pc [16] ), .QN(_08754_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08305_ ), .Q(\ID_EX_pc [15] ), .QN(_08755_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08305_ ), .Q(\ID_EX_pc [14] ), .QN(_08756_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08305_ ), .Q(\ID_EX_pc [13] ), .QN(_08757_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08305_ ), .Q(\ID_EX_pc [12] ), .QN(_08758_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08305_ ), .Q(\ID_EX_pc [29] ), .QN(_08759_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08305_ ), .Q(\ID_EX_pc [11] ), .QN(_08760_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08305_ ), .Q(\ID_EX_pc [10] ), .QN(_08761_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08305_ ), .Q(\ID_EX_pc [9] ), .QN(_08762_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08305_ ), .Q(\ID_EX_pc [8] ), .QN(_08763_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08305_ ), .Q(\ID_EX_pc [7] ), .QN(_08764_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08305_ ), .Q(\ID_EX_pc [6] ), .QN(_08765_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08305_ ), .Q(\ID_EX_pc [5] ), .QN(_08766_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08305_ ), .Q(\ID_EX_pc [4] ), .QN(_08767_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08305_ ), .Q(\ID_EX_pc [3] ), .QN(_08768_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08305_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08305_ ), .Q(\ID_EX_pc [28] ), .QN(_08769_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08305_ ), .Q(\ID_EX_pc [1] ), .QN(_08770_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08305_ ), .Q(\ID_EX_pc [0] ), .QN(_08771_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08305_ ), .Q(\ID_EX_pc [27] ), .QN(_08772_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08305_ ), .Q(\ID_EX_pc [26] ), .QN(_08773_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08305_ ), .Q(\ID_EX_pc [25] ), .QN(_08774_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08305_ ), .Q(\ID_EX_pc [24] ), .QN(_08775_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08305_ ), .Q(\ID_EX_pc [23] ), .QN(_08776_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08305_ ), .Q(\ID_EX_pc [22] ), .QN(_08406_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00209_ ), .CK(_08304_ ), .Q(\ID_EX_rd [4] ), .QN(_08405_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00210_ ), .CK(_08304_ ), .Q(\ID_EX_rd [3] ), .QN(_08404_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00211_ ), .CK(_08304_ ), .Q(\ID_EX_rd [2] ), .QN(_08403_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00212_ ), .CK(_08304_ ), .Q(\ID_EX_rd [1] ), .QN(_08402_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00213_ ), .CK(_08304_ ), .Q(\ID_EX_rd [0] ), .QN(_08401_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00214_ ), .CK(_08303_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08400_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00215_ ), .CK(_08303_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08399_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00217_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08397_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00216_ ), .CK(_08303_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08398_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00219_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08395_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00218_ ), .CK(_08303_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08396_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00221_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08393_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00220_ ), .CK(_08303_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08394_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00223_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08391_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00222_ ), .CK(_08302_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08392_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00224_ ), .CK(_08302_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08390_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00226_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08388_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00225_ ), .CK(_08302_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08389_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00228_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08386_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00227_ ), .CK(_08302_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08387_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00230_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08384_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00229_ ), .CK(_08302_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08385_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00232_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08382_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_08301_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08383_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00233_ ), .CK(_08300_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08381_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08778_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00234_ ), .CK(_08299_ ), .Q(\ID_EX_typ [7] ), .QN(_08777_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00235_ ), .CK(_08299_ ), .Q(\ID_EX_typ [6] ), .QN(_08380_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00236_ ), .CK(_08299_ ), .Q(\ID_EX_typ [5] ), .QN(_08379_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00237_ ), .CK(_08299_ ), .Q(\ID_EX_typ [4] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00238_ ), .CK(_08299_ ), .Q(\ID_EX_typ [3] ), .QN(_08378_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00239_ ), .CK(_08299_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00240_ ), .CK(_08299_ ), .Q(\ID_EX_typ [1] ), .QN(_08377_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00241_ ), .CK(_08299_ ), .Q(\ID_EX_typ [0] ), .QN(\myexu.pc_jump_$_SDFF_PP0__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08298_ ), .Q(check_assert ), .QN(_08779_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08297_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08297_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08297_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08297_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08297_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08297_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08297_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08297_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08297_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08297_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08297_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08297_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08297_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08297_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08297_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08297_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08297_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08297_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08297_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08297_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08297_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08297_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08297_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08297_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08297_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08297_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08297_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08297_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08297_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08297_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08297_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08297_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08296_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08295_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08855_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08856_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08857_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08858_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08859_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08860_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08861_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08862_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08863_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08864_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08865_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08866_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08867_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08868_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08869_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08870_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08871_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08872_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08873_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08874_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08294_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08875_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08876_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08877_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08878_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08879_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08880_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08881_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08882_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08883_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08884_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08885_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08886_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08887_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08888_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08889_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08890_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08891_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08892_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08893_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08894_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08895_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08896_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08897_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08898_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08899_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08900_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08901_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08902_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08903_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08904_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08905_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08906_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08293_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08907_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08908_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08909_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08910_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08911_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08912_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08913_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08914_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08915_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08916_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08917_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08918_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08919_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08920_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08921_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08922_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08923_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08924_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08925_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08926_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08927_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08928_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08929_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08930_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08931_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08932_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08933_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08934_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08935_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08936_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08937_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08938_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08292_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08939_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08940_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08941_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08942_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08943_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08944_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08945_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08946_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08947_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08948_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08949_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08950_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08951_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08952_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08953_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08954_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08955_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08956_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08957_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08958_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08959_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08960_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08961_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08962_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08963_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08964_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08965_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08966_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08967_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08968_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08969_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08970_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08291_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08971_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08972_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08973_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08974_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08975_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08976_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08977_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08978_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08979_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08980_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08981_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08982_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08983_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08984_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08985_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08986_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08987_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08988_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08989_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08990_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08991_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08992_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08993_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08994_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08995_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08996_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08997_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08998_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08999_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_09000_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_09001_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_09002_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08290_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_09003_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_09004_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_09005_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_09006_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_09007_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_09008_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_09009_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_09010_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_09011_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_09012_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_09013_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_09014_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_09015_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_09016_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_09017_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_09018_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_09019_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_09020_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_09021_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_09022_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_09023_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_09024_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_09025_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_09026_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_09027_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_09028_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_09029_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_09030_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_09031_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_09032_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_09033_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_09034_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08289_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_09035_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_09036_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_09037_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_09038_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_09039_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_09040_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_09041_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_09042_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_09043_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_09044_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_09045_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_09046_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_09047_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_09048_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_09049_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_09050_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_09051_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_09052_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_09053_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_09054_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_09055_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_09056_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_09057_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_09058_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_09059_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_09060_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_09061_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08288_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_09062_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_09063_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_09064_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_09065_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_09066_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_09067_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_09068_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_09069_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_09070_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_09071_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_09072_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_09073_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_09074_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_09075_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_09076_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_09077_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_09078_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_09079_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_09080_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_09081_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_09082_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_09083_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_09084_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_09085_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_09086_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_09087_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_09088_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08287_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_09089_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_09090_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_09091_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_09092_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_09093_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_09094_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_09095_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_09096_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_09097_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_09098_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_09099_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_09100_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_09101_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_09102_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_09103_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_09104_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_09105_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_09106_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_09107_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_09108_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_09109_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_09110_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_09111_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_09112_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_09113_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_09114_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_09115_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08286_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_09116_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_09117_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_09118_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_09119_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_09120_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_09121_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_09122_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_09123_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_09124_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_09125_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_09126_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_09127_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_09128_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_09129_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_09130_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_09131_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_09132_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_09133_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_09134_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_09135_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_09136_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_09137_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_09138_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_09139_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_09140_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_09141_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_09142_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08285_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08376_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00242_ ), .CK(_08284_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08375_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00243_ ), .CK(_08283_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08374_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00244_ ), .CK(_08282_ ), .Q(\myifu.myicache.valid [2] ), .QN(_09143_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_08281_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08373_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_08280_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_08279_ ), .Q(\IF_ID_pc [30] ), .QN(_08372_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00247_ ), .CK(_08279_ ), .Q(\IF_ID_pc [21] ), .QN(_08371_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00248_ ), .CK(_08279_ ), .Q(\IF_ID_pc [20] ), .QN(_08370_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00249_ ), .CK(_08279_ ), .Q(\IF_ID_pc [19] ), .QN(_08369_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00250_ ), .CK(_08279_ ), .Q(\IF_ID_pc [18] ), .QN(_08368_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00251_ ), .CK(_08279_ ), .Q(\IF_ID_pc [17] ), .QN(_08367_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00252_ ), .CK(_08279_ ), .Q(\IF_ID_pc [16] ), .QN(_08366_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00253_ ), .CK(_08279_ ), .Q(\IF_ID_pc [15] ), .QN(_08365_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00254_ ), .CK(_08279_ ), .Q(\IF_ID_pc [14] ), .QN(_08364_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00255_ ), .CK(_08279_ ), .Q(\IF_ID_pc [13] ), .QN(_08363_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00256_ ), .CK(_08279_ ), .Q(\IF_ID_pc [12] ), .QN(_08362_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00257_ ), .CK(_08279_ ), .Q(\IF_ID_pc [29] ), .QN(_08361_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00258_ ), .CK(_08279_ ), .Q(\IF_ID_pc [11] ), .QN(_08360_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00259_ ), .CK(_08279_ ), .Q(\IF_ID_pc [10] ), .QN(_08359_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00260_ ), .CK(_08279_ ), .Q(\IF_ID_pc [9] ), .QN(_08358_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00261_ ), .CK(_08279_ ), .Q(\IF_ID_pc [8] ), .QN(_08357_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00262_ ), .CK(_08279_ ), .Q(\IF_ID_pc [7] ), .QN(_08356_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00263_ ), .CK(_08279_ ), .Q(\IF_ID_pc [6] ), .QN(_08355_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00264_ ), .CK(_08279_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00265_ ), .CK(_08279_ ), .Q(\IF_ID_pc [4] ), .QN(_08354_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00267_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08353_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00266_ ), .CK(_08279_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00269_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08351_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00268_ ), .CK(_08279_ ), .Q(\IF_ID_pc [2] ), .QN(_08352_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00270_ ), .CK(_08279_ ), .Q(\IF_ID_pc [28] ), .QN(_08350_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00271_ ), .CK(_08279_ ), .Q(\IF_ID_pc [1] ), .QN(_08349_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00272_ ), .CK(_08279_ ), .Q(\IF_ID_pc [27] ), .QN(_08348_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00273_ ), .CK(_08279_ ), .Q(\IF_ID_pc [26] ), .QN(_08347_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00274_ ), .CK(_08279_ ), .Q(\IF_ID_pc [25] ), .QN(_08346_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00275_ ), .CK(_08279_ ), .Q(\IF_ID_pc [24] ), .QN(_08345_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00276_ ), .CK(_08279_ ), .Q(\IF_ID_pc [23] ), .QN(_08344_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00277_ ), .CK(_08279_ ), .Q(\IF_ID_pc [22] ), .QN(_08343_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00278_ ), .CK(_08279_ ), .Q(\IF_ID_pc [31] ), .QN(_08342_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_09145_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08341_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00279_ ), .CK(_08278_ ), .Q(\myifu.tmp_offset [2] ), .QN(_09144_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00281_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00280_ ), .CK(_08277_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08340_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_09146_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_09147_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_09148_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_09149_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_09150_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_09151_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_09152_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_09153_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_09154_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_09155_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_09156_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_09157_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_09158_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_09159_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_09160_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_09161_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_09162_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_09163_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_09164_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_09165_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_09166_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_09167_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_09168_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_09169_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_09170_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_09171_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_09172_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_09173_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_09174_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_09175_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_09176_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08276_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_09177_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_09178_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_09179_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_09180_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_09181_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_09182_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_09183_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_09184_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_09185_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_09186_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_09187_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_09188_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_09189_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_09190_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_09191_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_09192_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_09193_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_09194_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_09195_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_09196_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_09197_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_09198_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_09199_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_09200_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_09201_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_09202_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_09203_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_09204_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_09205_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_09206_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_09207_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_09208_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08275_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08339_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PP0P__Q ( .D(_00282_ ), .CK(_08274_ ), .Q(LS_WB_pc ), .QN(_08338_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PP0P__Q ( .D(_00283_ ), .CK(_08273_ ), .Q(\mylsu.previous_load_done ), .QN(_09209_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_09210_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_09211_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_09212_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(_09213_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_08276_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_08276_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_09214_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_08276_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08337_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00284_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08336_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00285_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08335_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00286_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08334_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00287_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08333_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00288_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08332_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00289_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08331_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00290_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08330_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00291_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08329_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00292_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08328_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00293_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08327_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00294_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08326_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00295_ ), .CK(_08276_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_09215_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_08276_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_09216_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_08276_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_09217_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_08276_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_09218_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_08276_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_09219_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_09220_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_09221_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_09222_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_09223_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_09224_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_09225_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_09226_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_09227_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_09228_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_09229_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_09230_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_09231_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_09232_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_09233_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_09234_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_09235_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_09236_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_09237_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_09238_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_09239_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_09240_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_09241_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_09242_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_09243_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_09244_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_09245_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_09246_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_09247_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_09248_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_09249_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_09250_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_08276_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_09251_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_09252_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_09253_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_09254_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_09255_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_09256_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_09257_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_09258_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_09259_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_09260_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_09261_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_09262_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_09263_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_09264_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_09265_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_09266_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_09267_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_09268_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_09269_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_09270_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_09271_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_09272_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_09273_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_09274_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_09275_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_09276_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_09277_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_09278_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_09279_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_09280_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_09281_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_09282_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_08272_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08325_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q ( .D(_00296_ ), .CK(_08271_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_08324_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_1 ( .D(_00297_ ), .CK(_08271_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08323_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_2 ( .D(_00298_ ), .CK(_08271_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08322_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_3 ( .D(_00299_ ), .CK(_08271_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08321_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_4 ( .D(_00300_ ), .CK(_08271_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08320_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_5 ( .D(_00301_ ), .CK(_08271_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08319_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PP0P__Q ( .D(_00302_ ), .CK(_08271_ ), .Q(LS_WB_wen_reg ), .QN(_09283_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_09284_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_09285_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08270_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08269_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08268_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08267_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08266_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08265_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08264_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08263_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08262_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08261_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08260_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08259_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08258_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08257_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08256_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08255_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00303_ ), .CK(_08254_ ), .Q(loaduse_clear ), .QN(_09286_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_09287_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_09288_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08318_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\ID_EX_typ [3] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(excp_written ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_44 ) );

endmodule
